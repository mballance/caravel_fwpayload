VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 28.980 2924.800 30.180 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2374.980 2924.800 2376.180 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2609.580 2924.800 2610.780 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2844.180 2924.800 2845.380 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3078.780 2924.800 3079.980 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3313.380 2924.800 3314.580 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 263.580 2924.800 264.780 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3482.700 2.400 3483.900 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3195.060 2.400 3196.260 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2908.100 2.400 2909.300 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2620.460 2.400 2621.660 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2333.500 2.400 2334.700 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2045.860 2.400 2047.060 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 498.180 2924.800 499.380 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1758.900 2.400 1760.100 ;
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 732.780 2924.800 733.980 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 967.380 2924.800 968.580 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1201.980 2924.800 1203.180 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1436.580 2924.800 1437.780 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1671.180 2924.800 1672.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1905.780 2924.800 1906.980 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2140.380 2924.800 2141.580 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1738.410 84.220 1738.730 84.280 ;
        RECT 1779.810 84.220 1780.130 84.280 ;
        RECT 1738.410 84.080 1780.130 84.220 ;
        RECT 1738.410 84.020 1738.730 84.080 ;
        RECT 1779.810 84.020 1780.130 84.080 ;
        RECT 2572.850 83.880 2573.170 83.940 ;
        RECT 2580.210 83.880 2580.530 83.940 ;
        RECT 2572.850 83.740 2580.530 83.880 ;
        RECT 2572.850 83.680 2573.170 83.740 ;
        RECT 2580.210 83.680 2580.530 83.740 ;
        RECT 1593.510 83.540 1593.830 83.600 ;
        RECT 1598.110 83.540 1598.430 83.600 ;
        RECT 1593.510 83.400 1598.430 83.540 ;
        RECT 1593.510 83.340 1593.830 83.400 ;
        RECT 1598.110 83.340 1598.430 83.400 ;
        RECT 1670.330 83.540 1670.650 83.600 ;
        RECT 1690.570 83.540 1690.890 83.600 ;
        RECT 1670.330 83.400 1690.890 83.540 ;
        RECT 1670.330 83.340 1670.650 83.400 ;
        RECT 1690.570 83.340 1690.890 83.400 ;
        RECT 2621.150 83.540 2621.470 83.600 ;
        RECT 2632.190 83.540 2632.510 83.600 ;
        RECT 2621.150 83.400 2632.510 83.540 ;
        RECT 2621.150 83.340 2621.470 83.400 ;
        RECT 2632.190 83.340 2632.510 83.400 ;
      LAYER via ;
        RECT 1738.440 84.020 1738.700 84.280 ;
        RECT 1779.840 84.020 1780.100 84.280 ;
        RECT 2572.880 83.680 2573.140 83.940 ;
        RECT 2580.240 83.680 2580.500 83.940 ;
        RECT 1593.540 83.340 1593.800 83.600 ;
        RECT 1598.140 83.340 1598.400 83.600 ;
        RECT 1670.360 83.340 1670.620 83.600 ;
        RECT 1690.600 83.340 1690.860 83.600 ;
        RECT 2621.180 83.340 2621.440 83.600 ;
        RECT 2632.220 83.340 2632.480 83.600 ;
      LAYER met2 ;
        RECT 1155.080 3196.410 1155.360 3200.000 ;
        RECT 1156.990 3196.410 1157.270 3196.525 ;
        RECT 1155.080 3196.270 1157.270 3196.410 ;
        RECT 1155.080 3196.000 1155.360 3196.270 ;
        RECT 1156.990 3196.155 1157.270 3196.270 ;
        RECT 1779.830 85.835 1780.110 86.205 ;
        RECT 1255.430 85.155 1255.710 85.525 ;
        RECT 1200.690 83.795 1200.970 84.165 ;
        RECT 1200.760 83.370 1200.900 83.795 ;
        RECT 1255.500 83.485 1255.640 85.155 ;
        RECT 1779.900 84.310 1780.040 85.835 ;
        RECT 2704.430 85.155 2704.710 85.525 ;
        RECT 2028.690 84.475 2028.970 84.845 ;
        RECT 2090.330 84.730 2090.610 84.845 ;
        RECT 2091.250 84.730 2091.530 84.845 ;
        RECT 2090.330 84.590 2091.530 84.730 ;
        RECT 2090.330 84.475 2090.610 84.590 ;
        RECT 2091.250 84.475 2091.530 84.590 ;
        RECT 1738.440 84.165 1738.700 84.310 ;
        RECT 1598.130 83.795 1598.410 84.165 ;
        RECT 1738.430 83.795 1738.710 84.165 ;
        RECT 1779.840 83.990 1780.100 84.310 ;
        RECT 2028.760 84.165 2028.900 84.475 ;
        RECT 2028.690 83.795 2028.970 84.165 ;
        RECT 2283.530 84.050 2283.810 84.165 ;
        RECT 2284.450 84.050 2284.730 84.165 ;
        RECT 2283.530 83.910 2284.730 84.050 ;
        RECT 2283.530 83.795 2283.810 83.910 ;
        RECT 2284.450 83.795 2284.730 83.910 ;
        RECT 2572.870 83.795 2573.150 84.165 ;
        RECT 2580.230 83.795 2580.510 84.165 ;
        RECT 2632.210 83.795 2632.490 84.165 ;
        RECT 1598.200 83.630 1598.340 83.795 ;
        RECT 2572.880 83.650 2573.140 83.795 ;
        RECT 2580.240 83.650 2580.500 83.795 ;
        RECT 2632.280 83.630 2632.420 83.795 ;
        RECT 1593.540 83.485 1593.800 83.630 ;
        RECT 1201.150 83.370 1201.430 83.485 ;
        RECT 1200.760 83.230 1201.430 83.370 ;
        RECT 1201.150 83.115 1201.430 83.230 ;
        RECT 1255.430 83.115 1255.710 83.485 ;
        RECT 1593.530 83.115 1593.810 83.485 ;
        RECT 1598.140 83.310 1598.400 83.630 ;
        RECT 1670.360 83.485 1670.620 83.630 ;
        RECT 1690.600 83.485 1690.860 83.630 ;
        RECT 2621.180 83.485 2621.440 83.630 ;
        RECT 1670.350 83.115 1670.630 83.485 ;
        RECT 1690.590 83.115 1690.870 83.485 ;
        RECT 2621.170 83.115 2621.450 83.485 ;
        RECT 2632.220 83.310 2632.480 83.630 ;
        RECT 2704.500 83.485 2704.640 85.155 ;
        RECT 2801.030 84.475 2801.310 84.845 ;
        RECT 2704.430 83.115 2704.710 83.485 ;
        RECT 2801.100 82.805 2801.240 84.475 ;
        RECT 2863.130 83.795 2863.410 84.165 ;
        RECT 2863.200 83.370 2863.340 83.795 ;
        RECT 2863.590 83.370 2863.870 83.485 ;
        RECT 2863.200 83.230 2863.870 83.370 ;
        RECT 2863.590 83.115 2863.870 83.230 ;
        RECT 2801.030 82.435 2801.310 82.805 ;
      LAYER via2 ;
        RECT 1156.990 3196.200 1157.270 3196.480 ;
        RECT 1779.830 85.880 1780.110 86.160 ;
        RECT 1255.430 85.200 1255.710 85.480 ;
        RECT 1200.690 83.840 1200.970 84.120 ;
        RECT 2704.430 85.200 2704.710 85.480 ;
        RECT 2028.690 84.520 2028.970 84.800 ;
        RECT 2090.330 84.520 2090.610 84.800 ;
        RECT 2091.250 84.520 2091.530 84.800 ;
        RECT 1598.130 83.840 1598.410 84.120 ;
        RECT 1738.430 83.840 1738.710 84.120 ;
        RECT 2028.690 83.840 2028.970 84.120 ;
        RECT 2283.530 83.840 2283.810 84.120 ;
        RECT 2284.450 83.840 2284.730 84.120 ;
        RECT 2572.870 83.840 2573.150 84.120 ;
        RECT 2580.230 83.840 2580.510 84.120 ;
        RECT 2632.210 83.840 2632.490 84.120 ;
        RECT 1201.150 83.160 1201.430 83.440 ;
        RECT 1255.430 83.160 1255.710 83.440 ;
        RECT 1593.530 83.160 1593.810 83.440 ;
        RECT 1670.350 83.160 1670.630 83.440 ;
        RECT 1690.590 83.160 1690.870 83.440 ;
        RECT 2621.170 83.160 2621.450 83.440 ;
        RECT 2801.030 84.520 2801.310 84.800 ;
        RECT 2704.430 83.160 2704.710 83.440 ;
        RECT 2863.130 83.840 2863.410 84.120 ;
        RECT 2863.590 83.160 2863.870 83.440 ;
        RECT 2801.030 82.480 2801.310 82.760 ;
      LAYER met3 ;
        RECT 1156.965 3196.490 1157.295 3196.505 ;
        RECT 1158.550 3196.490 1158.930 3196.500 ;
        RECT 1156.965 3196.190 1158.930 3196.490 ;
        RECT 1156.965 3196.175 1157.295 3196.190 ;
        RECT 1158.550 3196.180 1158.930 3196.190 ;
        RECT 2917.600 88.210 2924.800 88.660 ;
        RECT 2916.710 87.910 2924.800 88.210 ;
        RECT 1297.470 86.850 1297.850 86.860 ;
        RECT 1344.390 86.850 1344.770 86.860 ;
        RECT 1297.470 86.550 1344.770 86.850 ;
        RECT 1297.470 86.540 1297.850 86.550 ;
        RECT 1344.390 86.540 1344.770 86.550 ;
        RECT 1779.805 86.170 1780.135 86.185 ;
        RECT 1786.910 86.170 1787.290 86.180 ;
        RECT 1779.805 85.870 1787.290 86.170 ;
        RECT 1779.805 85.855 1780.135 85.870 ;
        RECT 1786.910 85.860 1787.290 85.870 ;
        RECT 1255.405 85.490 1255.735 85.505 ;
        RECT 1297.470 85.490 1297.850 85.500 ;
        RECT 1255.405 85.190 1297.850 85.490 ;
        RECT 1255.405 85.175 1255.735 85.190 ;
        RECT 1297.470 85.180 1297.850 85.190 ;
        RECT 1835.670 85.490 1836.050 85.500 ;
        RECT 1835.670 85.190 1836.930 85.490 ;
        RECT 1835.670 85.180 1836.050 85.190 ;
        RECT 1532.070 84.810 1532.450 84.820 ;
        RECT 1400.550 84.510 1414.650 84.810 ;
        RECT 1158.550 84.130 1158.930 84.140 ;
        RECT 1200.665 84.130 1200.995 84.145 ;
        RECT 1158.550 83.830 1200.995 84.130 ;
        RECT 1158.550 83.820 1158.930 83.830 ;
        RECT 1200.665 83.815 1200.995 83.830 ;
        RECT 1201.125 83.450 1201.455 83.465 ;
        RECT 1255.405 83.450 1255.735 83.465 ;
        RECT 1400.550 83.450 1400.850 84.510 ;
        RECT 1201.125 83.150 1255.735 83.450 ;
        RECT 1201.125 83.135 1201.455 83.150 ;
        RECT 1255.405 83.135 1255.735 83.150 ;
        RECT 1366.510 83.150 1400.850 83.450 ;
        RECT 1414.350 83.450 1414.650 84.510 ;
        RECT 1519.230 84.510 1532.450 84.810 ;
        RECT 1414.350 83.150 1449.610 83.450 ;
        RECT 1345.310 82.770 1345.690 82.780 ;
        RECT 1366.510 82.770 1366.810 83.150 ;
        RECT 1345.310 82.470 1366.810 82.770 ;
        RECT 1449.310 82.770 1449.610 83.150 ;
        RECT 1519.230 82.770 1519.530 84.510 ;
        RECT 1532.070 84.500 1532.450 84.510 ;
        RECT 1786.910 84.810 1787.290 84.820 ;
        RECT 1836.630 84.810 1836.930 85.190 ;
        RECT 2125.470 85.180 2125.850 85.500 ;
        RECT 2510.030 85.490 2510.410 85.500 ;
        RECT 2476.030 85.190 2510.410 85.490 ;
        RECT 2028.665 84.810 2028.995 84.825 ;
        RECT 2090.305 84.810 2090.635 84.825 ;
        RECT 1786.910 84.510 1788.170 84.810 ;
        RECT 1836.630 84.510 1907.770 84.810 ;
        RECT 1786.910 84.500 1787.290 84.510 ;
        RECT 1598.105 84.130 1598.435 84.145 ;
        RECT 1738.405 84.130 1738.735 84.145 ;
        RECT 1598.105 83.830 1645.570 84.130 ;
        RECT 1598.105 83.815 1598.435 83.830 ;
        RECT 1532.990 83.450 1533.370 83.460 ;
        RECT 1593.505 83.450 1593.835 83.465 ;
        RECT 1532.990 83.150 1593.835 83.450 ;
        RECT 1645.270 83.450 1645.570 83.830 ;
        RECT 1731.750 83.830 1738.735 84.130 ;
        RECT 1787.870 84.130 1788.170 84.510 ;
        RECT 1835.670 84.130 1836.050 84.140 ;
        RECT 1787.870 83.830 1836.050 84.130 ;
        RECT 1907.470 84.130 1907.770 84.510 ;
        RECT 1955.310 84.510 2004.370 84.810 ;
        RECT 1955.310 84.130 1955.610 84.510 ;
        RECT 1907.470 83.830 1955.610 84.130 ;
        RECT 2004.070 84.130 2004.370 84.510 ;
        RECT 2028.665 84.510 2090.635 84.810 ;
        RECT 2028.665 84.495 2028.995 84.510 ;
        RECT 2090.305 84.495 2090.635 84.510 ;
        RECT 2091.225 84.810 2091.555 84.825 ;
        RECT 2125.510 84.810 2125.810 85.180 ;
        RECT 2091.225 84.510 2125.810 84.810 ;
        RECT 2138.390 84.510 2187.450 84.810 ;
        RECT 2091.225 84.495 2091.555 84.510 ;
        RECT 2028.665 84.130 2028.995 84.145 ;
        RECT 2004.070 83.830 2028.995 84.130 ;
        RECT 1670.325 83.450 1670.655 83.465 ;
        RECT 1645.270 83.150 1670.655 83.450 ;
        RECT 1532.990 83.140 1533.370 83.150 ;
        RECT 1593.505 83.135 1593.835 83.150 ;
        RECT 1670.325 83.135 1670.655 83.150 ;
        RECT 1690.565 83.450 1690.895 83.465 ;
        RECT 1731.750 83.450 1732.050 83.830 ;
        RECT 1738.405 83.815 1738.735 83.830 ;
        RECT 1835.670 83.820 1836.050 83.830 ;
        RECT 2028.665 83.815 2028.995 83.830 ;
        RECT 2125.470 84.130 2125.850 84.140 ;
        RECT 2138.390 84.130 2138.690 84.510 ;
        RECT 2125.470 83.830 2138.690 84.130 ;
        RECT 2125.470 83.820 2125.850 83.830 ;
        RECT 1690.565 83.150 1732.050 83.450 ;
        RECT 2187.150 83.450 2187.450 84.510 ;
        RECT 2283.505 84.130 2283.835 84.145 ;
        RECT 2235.910 83.830 2283.835 84.130 ;
        RECT 2235.910 83.450 2236.210 83.830 ;
        RECT 2283.505 83.815 2283.835 83.830 ;
        RECT 2284.425 84.130 2284.755 84.145 ;
        RECT 2476.030 84.130 2476.330 85.190 ;
        RECT 2510.030 85.180 2510.410 85.190 ;
        RECT 2656.310 85.490 2656.690 85.500 ;
        RECT 2704.405 85.490 2704.735 85.505 ;
        RECT 2656.310 85.190 2704.735 85.490 ;
        RECT 2656.310 85.180 2656.690 85.190 ;
        RECT 2704.405 85.175 2704.735 85.190 ;
        RECT 2801.005 84.810 2801.335 84.825 ;
        RECT 2801.005 84.510 2815.810 84.810 ;
        RECT 2801.005 84.495 2801.335 84.510 ;
        RECT 2572.845 84.130 2573.175 84.145 ;
        RECT 2284.425 83.830 2331.890 84.130 ;
        RECT 2284.425 83.815 2284.755 83.830 ;
        RECT 2187.150 83.150 2236.210 83.450 ;
        RECT 2331.590 83.450 2331.890 83.830 ;
        RECT 2332.510 83.830 2414.690 84.130 ;
        RECT 2332.510 83.450 2332.810 83.830 ;
        RECT 2331.590 83.150 2332.810 83.450 ;
        RECT 2414.390 83.450 2414.690 83.830 ;
        RECT 2429.110 83.830 2476.330 84.130 ;
        RECT 2525.710 83.830 2573.175 84.130 ;
        RECT 2429.110 83.450 2429.410 83.830 ;
        RECT 2414.390 83.150 2429.410 83.450 ;
        RECT 2510.950 83.450 2511.330 83.460 ;
        RECT 2525.710 83.450 2526.010 83.830 ;
        RECT 2572.845 83.815 2573.175 83.830 ;
        RECT 2580.205 84.130 2580.535 84.145 ;
        RECT 2632.185 84.130 2632.515 84.145 ;
        RECT 2656.310 84.130 2656.690 84.140 ;
        RECT 2752.910 84.130 2753.290 84.140 ;
        RECT 2580.205 83.830 2607.890 84.130 ;
        RECT 2580.205 83.815 2580.535 83.830 ;
        RECT 2510.950 83.150 2526.010 83.450 ;
        RECT 2607.590 83.450 2607.890 83.830 ;
        RECT 2632.185 83.830 2656.690 84.130 ;
        RECT 2632.185 83.815 2632.515 83.830 ;
        RECT 2656.310 83.820 2656.690 83.830 ;
        RECT 2718.910 83.830 2753.290 84.130 ;
        RECT 2621.145 83.450 2621.475 83.465 ;
        RECT 2607.590 83.150 2621.475 83.450 ;
        RECT 1690.565 83.135 1690.895 83.150 ;
        RECT 2510.950 83.140 2511.330 83.150 ;
        RECT 2621.145 83.135 2621.475 83.150 ;
        RECT 2704.405 83.450 2704.735 83.465 ;
        RECT 2718.910 83.450 2719.210 83.830 ;
        RECT 2752.910 83.820 2753.290 83.830 ;
        RECT 2704.405 83.150 2719.210 83.450 ;
        RECT 2815.510 83.450 2815.810 84.510 ;
        RECT 2863.105 84.130 2863.435 84.145 ;
        RECT 2916.710 84.130 2917.010 87.910 ;
        RECT 2917.600 87.460 2924.800 87.910 ;
        RECT 2849.550 83.830 2863.435 84.130 ;
        RECT 2849.550 83.450 2849.850 83.830 ;
        RECT 2863.105 83.815 2863.435 83.830 ;
        RECT 2884.510 83.830 2917.010 84.130 ;
        RECT 2815.510 83.150 2849.850 83.450 ;
        RECT 2863.565 83.450 2863.895 83.465 ;
        RECT 2884.510 83.450 2884.810 83.830 ;
        RECT 2863.565 83.150 2884.810 83.450 ;
        RECT 2704.405 83.135 2704.735 83.150 ;
        RECT 2863.565 83.135 2863.895 83.150 ;
        RECT 1449.310 82.470 1519.530 82.770 ;
        RECT 2752.910 82.770 2753.290 82.780 ;
        RECT 2801.005 82.770 2801.335 82.785 ;
        RECT 2752.910 82.470 2801.335 82.770 ;
        RECT 1345.310 82.460 1345.690 82.470 ;
        RECT 2752.910 82.460 2753.290 82.470 ;
        RECT 2801.005 82.455 2801.335 82.470 ;
      LAYER via3 ;
        RECT 1158.580 3196.180 1158.900 3196.500 ;
        RECT 1297.500 86.540 1297.820 86.860 ;
        RECT 1344.420 86.540 1344.740 86.860 ;
        RECT 1786.940 85.860 1787.260 86.180 ;
        RECT 1297.500 85.180 1297.820 85.500 ;
        RECT 1835.700 85.180 1836.020 85.500 ;
        RECT 1158.580 83.820 1158.900 84.140 ;
        RECT 1345.340 82.460 1345.660 82.780 ;
        RECT 1532.100 84.500 1532.420 84.820 ;
        RECT 1786.940 84.500 1787.260 84.820 ;
        RECT 2125.500 85.180 2125.820 85.500 ;
        RECT 1533.020 83.140 1533.340 83.460 ;
        RECT 1835.700 83.820 1836.020 84.140 ;
        RECT 2125.500 83.820 2125.820 84.140 ;
        RECT 2510.060 85.180 2510.380 85.500 ;
        RECT 2656.340 85.180 2656.660 85.500 ;
        RECT 2510.980 83.140 2511.300 83.460 ;
        RECT 2656.340 83.820 2656.660 84.140 ;
        RECT 2752.940 83.820 2753.260 84.140 ;
        RECT 2752.940 82.460 2753.260 82.780 ;
      LAYER met4 ;
        RECT 1158.575 3196.175 1158.905 3196.505 ;
        RECT 1158.590 84.145 1158.890 3196.175 ;
        RECT 1297.495 86.535 1297.825 86.865 ;
        RECT 1344.415 86.535 1344.745 86.865 ;
        RECT 1532.110 86.550 1533.330 86.850 ;
        RECT 1297.510 85.505 1297.810 86.535 ;
        RECT 1297.495 85.175 1297.825 85.505 ;
        RECT 1158.575 83.815 1158.905 84.145 ;
        RECT 1344.430 83.450 1344.730 86.535 ;
        RECT 1532.110 84.825 1532.410 86.550 ;
        RECT 1532.095 84.495 1532.425 84.825 ;
        RECT 1533.030 83.465 1533.330 86.550 ;
        RECT 1786.935 85.855 1787.265 86.185 ;
        RECT 1786.950 84.825 1787.250 85.855 ;
        RECT 1835.695 85.175 1836.025 85.505 ;
        RECT 2125.495 85.175 2125.825 85.505 ;
        RECT 2510.055 85.175 2510.385 85.505 ;
        RECT 2656.335 85.175 2656.665 85.505 ;
        RECT 1786.935 84.495 1787.265 84.825 ;
        RECT 1835.710 84.145 1836.010 85.175 ;
        RECT 2125.510 84.145 2125.810 85.175 ;
        RECT 1835.695 83.815 1836.025 84.145 ;
        RECT 2125.495 83.815 2125.825 84.145 ;
        RECT 1344.430 83.150 1345.650 83.450 ;
        RECT 1345.350 82.785 1345.650 83.150 ;
        RECT 1533.015 83.135 1533.345 83.465 ;
        RECT 2510.070 83.450 2510.370 85.175 ;
        RECT 2656.350 84.145 2656.650 85.175 ;
        RECT 2656.335 83.815 2656.665 84.145 ;
        RECT 2752.935 83.815 2753.265 84.145 ;
        RECT 2510.975 83.450 2511.305 83.465 ;
        RECT 2510.070 83.150 2511.305 83.450 ;
        RECT 2510.975 83.135 2511.305 83.150 ;
        RECT 2752.950 82.785 2753.250 83.815 ;
        RECT 1345.335 82.455 1345.665 82.785 ;
        RECT 2752.935 82.455 2753.265 82.785 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1549.810 3213.920 1550.130 3213.980 ;
        RECT 2900.830 3213.920 2901.150 3213.980 ;
        RECT 1549.810 3213.780 2901.150 3213.920 ;
        RECT 1549.810 3213.720 1550.130 3213.780 ;
        RECT 2900.830 3213.720 2901.150 3213.780 ;
      LAYER via ;
        RECT 1549.840 3213.720 1550.100 3213.980 ;
        RECT 2900.860 3213.720 2901.120 3213.980 ;
      LAYER met2 ;
        RECT 1549.840 3213.690 1550.100 3214.010 ;
        RECT 2900.860 3213.690 2901.120 3214.010 ;
        RECT 1549.900 3200.000 1550.040 3213.690 ;
        RECT 1549.760 3196.000 1550.040 3200.000 ;
        RECT 2900.920 2434.245 2901.060 3213.690 ;
        RECT 2900.850 2433.875 2901.130 2434.245 ;
      LAYER via2 ;
        RECT 2900.850 2433.920 2901.130 2434.200 ;
      LAYER met3 ;
        RECT 2900.825 2434.210 2901.155 2434.225 ;
        RECT 2917.600 2434.210 2924.800 2434.660 ;
        RECT 2900.825 2433.910 2924.800 2434.210 ;
        RECT 2900.825 2433.895 2901.155 2433.910 ;
        RECT 2917.600 2433.460 2924.800 2433.910 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1588.930 3213.835 1589.210 3214.205 ;
        RECT 1589.000 3200.000 1589.140 3213.835 ;
        RECT 1588.860 3196.000 1589.140 3200.000 ;
      LAYER via2 ;
        RECT 1588.930 3213.880 1589.210 3214.160 ;
      LAYER met3 ;
        RECT 1588.905 3214.170 1589.235 3214.185 ;
        RECT 2636.990 3214.170 2637.370 3214.180 ;
        RECT 1588.905 3213.870 2637.370 3214.170 ;
        RECT 1588.905 3213.855 1589.235 3213.870 ;
        RECT 2636.990 3213.860 2637.370 3213.870 ;
        RECT 2637.910 3187.340 2638.290 3187.660 ;
        RECT 2637.950 3186.970 2638.250 3187.340 ;
        RECT 2640.670 3186.970 2641.050 3186.980 ;
        RECT 2637.950 3186.670 2641.050 3186.970 ;
        RECT 2640.670 3186.660 2641.050 3186.670 ;
        RECT 2640.670 3140.730 2641.050 3140.740 ;
        RECT 2637.030 3140.430 2641.050 3140.730 ;
        RECT 2637.030 3140.060 2637.330 3140.430 ;
        RECT 2640.670 3140.420 2641.050 3140.430 ;
        RECT 2636.990 3139.740 2637.370 3140.060 ;
        RECT 2636.990 3105.370 2637.370 3105.380 ;
        RECT 2641.590 3105.370 2641.970 3105.380 ;
        RECT 2636.990 3105.070 2641.970 3105.370 ;
        RECT 2636.990 3105.060 2637.370 3105.070 ;
        RECT 2641.590 3105.060 2641.970 3105.070 ;
        RECT 2641.590 3090.780 2641.970 3091.100 ;
        RECT 2641.630 3090.410 2641.930 3090.780 ;
        RECT 2644.350 3090.410 2644.730 3090.420 ;
        RECT 2641.630 3090.110 2644.730 3090.410 ;
        RECT 2644.350 3090.100 2644.730 3090.110 ;
        RECT 2642.510 3043.490 2642.890 3043.500 ;
        RECT 2644.350 3043.490 2644.730 3043.500 ;
        RECT 2642.510 3043.190 2644.730 3043.490 ;
        RECT 2642.510 3043.180 2642.890 3043.190 ;
        RECT 2644.350 3043.180 2644.730 3043.190 ;
        RECT 2637.910 3008.810 2638.290 3008.820 ;
        RECT 2642.510 3008.810 2642.890 3008.820 ;
        RECT 2637.910 3008.510 2642.890 3008.810 ;
        RECT 2637.910 3008.500 2638.290 3008.510 ;
        RECT 2642.510 3008.500 2642.890 3008.510 ;
        RECT 2637.910 2960.900 2638.290 2961.220 ;
        RECT 2637.950 2959.860 2638.250 2960.900 ;
        RECT 2637.910 2959.540 2638.290 2959.860 ;
        RECT 2636.990 2947.610 2637.370 2947.620 ;
        RECT 2637.910 2947.610 2638.290 2947.620 ;
        RECT 2636.990 2947.310 2638.290 2947.610 ;
        RECT 2636.990 2947.300 2637.370 2947.310 ;
        RECT 2637.910 2947.300 2638.290 2947.310 ;
        RECT 2637.910 2851.050 2638.290 2851.060 ;
        RECT 2637.030 2850.750 2638.290 2851.050 ;
        RECT 2637.030 2850.380 2637.330 2850.750 ;
        RECT 2637.910 2850.740 2638.290 2850.750 ;
        RECT 2636.990 2850.060 2637.370 2850.380 ;
        RECT 2636.990 2842.890 2637.370 2842.900 ;
        RECT 2640.670 2842.890 2641.050 2842.900 ;
        RECT 2636.990 2842.590 2641.050 2842.890 ;
        RECT 2636.990 2842.580 2637.370 2842.590 ;
        RECT 2640.670 2842.580 2641.050 2842.590 ;
        RECT 2640.670 2795.970 2641.050 2795.980 ;
        RECT 2637.950 2795.670 2641.050 2795.970 ;
        RECT 2637.950 2795.300 2638.250 2795.670 ;
        RECT 2640.670 2795.660 2641.050 2795.670 ;
        RECT 2637.910 2794.980 2638.290 2795.300 ;
        RECT 2637.910 2769.820 2638.290 2770.140 ;
        RECT 2637.950 2768.770 2638.250 2769.820 ;
        RECT 2639.750 2768.770 2640.130 2768.780 ;
        RECT 2637.950 2768.470 2640.130 2768.770 ;
        RECT 2639.750 2768.460 2640.130 2768.470 ;
        RECT 2639.750 2766.730 2640.130 2766.740 ;
        RECT 2637.950 2766.430 2640.130 2766.730 ;
        RECT 2637.950 2765.380 2638.250 2766.430 ;
        RECT 2639.750 2766.420 2640.130 2766.430 ;
        RECT 2637.910 2765.060 2638.290 2765.380 ;
        RECT 2917.600 2669.490 2924.800 2669.940 ;
        RECT 2916.710 2669.190 2924.800 2669.490 ;
        RECT 2637.910 2668.500 2638.290 2668.820 ;
        RECT 2637.950 2664.050 2638.250 2668.500 ;
        RECT 2691.310 2665.110 2739.450 2665.410 ;
        RECT 2691.310 2664.050 2691.610 2665.110 ;
        RECT 2739.150 2664.730 2739.450 2665.110 ;
        RECT 2787.910 2665.110 2836.050 2665.410 ;
        RECT 2739.150 2664.430 2787.290 2664.730 ;
        RECT 2637.950 2663.750 2691.610 2664.050 ;
        RECT 2786.990 2664.050 2787.290 2664.430 ;
        RECT 2787.910 2664.050 2788.210 2665.110 ;
        RECT 2835.750 2664.730 2836.050 2665.110 ;
        RECT 2835.750 2664.430 2883.890 2664.730 ;
        RECT 2786.990 2663.750 2788.210 2664.050 ;
        RECT 2883.590 2664.050 2883.890 2664.430 ;
        RECT 2916.710 2664.050 2917.010 2669.190 ;
        RECT 2917.600 2668.740 2924.800 2669.190 ;
        RECT 2883.590 2663.750 2917.010 2664.050 ;
      LAYER via3 ;
        RECT 2637.020 3213.860 2637.340 3214.180 ;
        RECT 2637.940 3187.340 2638.260 3187.660 ;
        RECT 2640.700 3186.660 2641.020 3186.980 ;
        RECT 2640.700 3140.420 2641.020 3140.740 ;
        RECT 2637.020 3139.740 2637.340 3140.060 ;
        RECT 2637.020 3105.060 2637.340 3105.380 ;
        RECT 2641.620 3105.060 2641.940 3105.380 ;
        RECT 2641.620 3090.780 2641.940 3091.100 ;
        RECT 2644.380 3090.100 2644.700 3090.420 ;
        RECT 2642.540 3043.180 2642.860 3043.500 ;
        RECT 2644.380 3043.180 2644.700 3043.500 ;
        RECT 2637.940 3008.500 2638.260 3008.820 ;
        RECT 2642.540 3008.500 2642.860 3008.820 ;
        RECT 2637.940 2960.900 2638.260 2961.220 ;
        RECT 2637.940 2959.540 2638.260 2959.860 ;
        RECT 2637.020 2947.300 2637.340 2947.620 ;
        RECT 2637.940 2947.300 2638.260 2947.620 ;
        RECT 2637.940 2850.740 2638.260 2851.060 ;
        RECT 2637.020 2850.060 2637.340 2850.380 ;
        RECT 2637.020 2842.580 2637.340 2842.900 ;
        RECT 2640.700 2842.580 2641.020 2842.900 ;
        RECT 2640.700 2795.660 2641.020 2795.980 ;
        RECT 2637.940 2794.980 2638.260 2795.300 ;
        RECT 2637.940 2769.820 2638.260 2770.140 ;
        RECT 2639.780 2768.460 2640.100 2768.780 ;
        RECT 2639.780 2766.420 2640.100 2766.740 ;
        RECT 2637.940 2765.060 2638.260 2765.380 ;
        RECT 2637.940 2668.500 2638.260 2668.820 ;
      LAYER met4 ;
        RECT 2637.015 3213.855 2637.345 3214.185 ;
        RECT 2637.030 3189.010 2637.330 3213.855 ;
        RECT 2637.030 3188.710 2638.250 3189.010 ;
        RECT 2637.950 3187.665 2638.250 3188.710 ;
        RECT 2637.935 3187.335 2638.265 3187.665 ;
        RECT 2640.695 3186.655 2641.025 3186.985 ;
        RECT 2640.710 3140.745 2641.010 3186.655 ;
        RECT 2640.695 3140.415 2641.025 3140.745 ;
        RECT 2637.015 3139.735 2637.345 3140.065 ;
        RECT 2637.030 3105.385 2637.330 3139.735 ;
        RECT 2637.015 3105.055 2637.345 3105.385 ;
        RECT 2641.615 3105.055 2641.945 3105.385 ;
        RECT 2641.630 3091.105 2641.930 3105.055 ;
        RECT 2641.615 3090.775 2641.945 3091.105 ;
        RECT 2644.375 3090.095 2644.705 3090.425 ;
        RECT 2644.390 3043.505 2644.690 3090.095 ;
        RECT 2642.535 3043.175 2642.865 3043.505 ;
        RECT 2644.375 3043.175 2644.705 3043.505 ;
        RECT 2642.550 3008.825 2642.850 3043.175 ;
        RECT 2637.935 3008.495 2638.265 3008.825 ;
        RECT 2642.535 3008.495 2642.865 3008.825 ;
        RECT 2637.950 2961.225 2638.250 3008.495 ;
        RECT 2637.935 2960.895 2638.265 2961.225 ;
        RECT 2637.935 2959.535 2638.265 2959.865 ;
        RECT 2637.950 2947.625 2638.250 2959.535 ;
        RECT 2637.015 2947.295 2637.345 2947.625 ;
        RECT 2637.935 2947.295 2638.265 2947.625 ;
        RECT 2637.030 2946.250 2637.330 2947.295 ;
        RECT 2637.030 2945.950 2639.170 2946.250 ;
        RECT 2638.870 2942.850 2639.170 2945.950 ;
        RECT 2637.950 2942.550 2639.170 2942.850 ;
        RECT 2637.950 2898.650 2638.250 2942.550 ;
        RECT 2637.950 2898.350 2639.170 2898.650 ;
        RECT 2638.870 2864.650 2639.170 2898.350 ;
        RECT 2637.950 2864.350 2639.170 2864.650 ;
        RECT 2637.950 2851.065 2638.250 2864.350 ;
        RECT 2637.935 2850.735 2638.265 2851.065 ;
        RECT 2637.015 2850.055 2637.345 2850.385 ;
        RECT 2637.030 2842.905 2637.330 2850.055 ;
        RECT 2637.015 2842.575 2637.345 2842.905 ;
        RECT 2640.695 2842.575 2641.025 2842.905 ;
        RECT 2640.710 2795.985 2641.010 2842.575 ;
        RECT 2640.695 2795.655 2641.025 2795.985 ;
        RECT 2637.935 2794.975 2638.265 2795.305 ;
        RECT 2637.950 2770.145 2638.250 2794.975 ;
        RECT 2637.935 2769.815 2638.265 2770.145 ;
        RECT 2639.775 2768.455 2640.105 2768.785 ;
        RECT 2639.790 2766.745 2640.090 2768.455 ;
        RECT 2639.775 2766.415 2640.105 2766.745 ;
        RECT 2637.935 2765.055 2638.265 2765.385 ;
        RECT 2637.950 2668.825 2638.250 2765.055 ;
        RECT 2637.935 2668.495 2638.265 2668.825 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1629.850 3198.960 1630.170 3199.020 ;
        RECT 2648.290 3198.960 2648.610 3199.020 ;
        RECT 1629.850 3198.820 2648.610 3198.960 ;
        RECT 1629.850 3198.760 1630.170 3198.820 ;
        RECT 2648.290 3198.760 2648.610 3198.820 ;
        RECT 2648.290 2904.860 2648.610 2904.920 ;
        RECT 2900.370 2904.860 2900.690 2904.920 ;
        RECT 2648.290 2904.720 2900.690 2904.860 ;
        RECT 2648.290 2904.660 2648.610 2904.720 ;
        RECT 2900.370 2904.660 2900.690 2904.720 ;
      LAYER via ;
        RECT 1629.880 3198.760 1630.140 3199.020 ;
        RECT 2648.320 3198.760 2648.580 3199.020 ;
        RECT 2648.320 2904.660 2648.580 2904.920 ;
        RECT 2900.400 2904.660 2900.660 2904.920 ;
      LAYER met2 ;
        RECT 1628.420 3199.130 1628.700 3200.000 ;
        RECT 1628.420 3199.050 1630.080 3199.130 ;
        RECT 1628.420 3198.990 1630.140 3199.050 ;
        RECT 1628.420 3196.000 1628.700 3198.990 ;
        RECT 1629.880 3198.730 1630.140 3198.990 ;
        RECT 2648.320 3198.730 2648.580 3199.050 ;
        RECT 2648.380 2904.950 2648.520 3198.730 ;
        RECT 2648.320 2904.630 2648.580 2904.950 ;
        RECT 2900.400 2904.630 2900.660 2904.950 ;
        RECT 2900.460 2904.125 2900.600 2904.630 ;
        RECT 2900.390 2903.755 2900.670 2904.125 ;
      LAYER via2 ;
        RECT 2900.390 2903.800 2900.670 2904.080 ;
      LAYER met3 ;
        RECT 2900.365 2904.090 2900.695 2904.105 ;
        RECT 2917.600 2904.090 2924.800 2904.540 ;
        RECT 2900.365 2903.790 2924.800 2904.090 ;
        RECT 2900.365 2903.775 2900.695 2903.790 ;
        RECT 2917.600 2903.340 2924.800 2903.790 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1669.410 3199.300 1669.730 3199.360 ;
        RECT 2648.750 3199.300 2649.070 3199.360 ;
        RECT 1669.410 3199.160 2649.070 3199.300 ;
        RECT 1669.410 3199.100 1669.730 3199.160 ;
        RECT 2648.750 3199.100 2649.070 3199.160 ;
        RECT 2648.750 3139.460 2649.070 3139.520 ;
        RECT 2900.370 3139.460 2900.690 3139.520 ;
        RECT 2648.750 3139.320 2900.690 3139.460 ;
        RECT 2648.750 3139.260 2649.070 3139.320 ;
        RECT 2900.370 3139.260 2900.690 3139.320 ;
      LAYER via ;
        RECT 1669.440 3199.100 1669.700 3199.360 ;
        RECT 2648.780 3199.100 2649.040 3199.360 ;
        RECT 2648.780 3139.260 2649.040 3139.520 ;
        RECT 2900.400 3139.260 2900.660 3139.520 ;
      LAYER met2 ;
        RECT 1667.980 3199.130 1668.260 3200.000 ;
        RECT 1669.440 3199.130 1669.700 3199.390 ;
        RECT 1667.980 3199.070 1669.700 3199.130 ;
        RECT 2648.780 3199.070 2649.040 3199.390 ;
        RECT 1667.980 3198.990 1669.640 3199.070 ;
        RECT 1667.980 3196.000 1668.260 3198.990 ;
        RECT 2648.840 3139.550 2648.980 3199.070 ;
        RECT 2648.780 3139.230 2649.040 3139.550 ;
        RECT 2900.400 3139.230 2900.660 3139.550 ;
        RECT 2900.460 3138.725 2900.600 3139.230 ;
        RECT 2900.390 3138.355 2900.670 3138.725 ;
      LAYER via2 ;
        RECT 2900.390 3138.400 2900.670 3138.680 ;
      LAYER met3 ;
        RECT 2900.365 3138.690 2900.695 3138.705 ;
        RECT 2917.600 3138.690 2924.800 3139.140 ;
        RECT 2900.365 3138.390 2924.800 3138.690 ;
        RECT 2900.365 3138.375 2900.695 3138.390 ;
        RECT 2917.600 3137.940 2924.800 3138.390 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1710.810 3367.600 1711.130 3367.660 ;
        RECT 2900.830 3367.600 2901.150 3367.660 ;
        RECT 1710.810 3367.460 2901.150 3367.600 ;
        RECT 1710.810 3367.400 1711.130 3367.460 ;
        RECT 2900.830 3367.400 2901.150 3367.460 ;
      LAYER via ;
        RECT 1710.840 3367.400 1711.100 3367.660 ;
        RECT 2900.860 3367.400 2901.120 3367.660 ;
      LAYER met2 ;
        RECT 2900.850 3372.955 2901.130 3373.325 ;
        RECT 2900.920 3367.690 2901.060 3372.955 ;
        RECT 1710.840 3367.370 1711.100 3367.690 ;
        RECT 2900.860 3367.370 2901.120 3367.690 ;
        RECT 1710.900 3200.490 1711.040 3367.370 ;
        RECT 1709.060 3200.350 1711.040 3200.490 ;
        RECT 1707.540 3199.810 1707.820 3200.000 ;
        RECT 1709.060 3199.810 1709.200 3200.350 ;
        RECT 1707.540 3199.670 1709.200 3199.810 ;
        RECT 1707.540 3196.000 1707.820 3199.670 ;
      LAYER via2 ;
        RECT 2900.850 3373.000 2901.130 3373.280 ;
      LAYER met3 ;
        RECT 2900.825 3373.290 2901.155 3373.305 ;
        RECT 2917.600 3373.290 2924.800 3373.740 ;
        RECT 2900.825 3372.990 2924.800 3373.290 ;
        RECT 2900.825 3372.975 2901.155 3372.990 ;
        RECT 2917.600 3372.540 2924.800 3372.990 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2796.485 3332.765 2796.655 3422.355 ;
        RECT 2796.025 3236.205 2796.195 3284.315 ;
      LAYER mcon ;
        RECT 2796.485 3422.185 2796.655 3422.355 ;
        RECT 2796.025 3284.145 2796.195 3284.315 ;
      LAYER met1 ;
        RECT 2795.490 3443.080 2795.810 3443.140 ;
        RECT 2798.250 3443.080 2798.570 3443.140 ;
        RECT 2795.490 3442.940 2798.570 3443.080 ;
        RECT 2795.490 3442.880 2795.810 3442.940 ;
        RECT 2798.250 3442.880 2798.570 3442.940 ;
        RECT 2795.030 3422.340 2795.350 3422.400 ;
        RECT 2796.425 3422.340 2796.715 3422.385 ;
        RECT 2795.030 3422.200 2796.715 3422.340 ;
        RECT 2795.030 3422.140 2795.350 3422.200 ;
        RECT 2796.425 3422.155 2796.715 3422.200 ;
        RECT 2796.425 3332.920 2796.715 3332.965 ;
        RECT 2796.870 3332.920 2797.190 3332.980 ;
        RECT 2796.425 3332.780 2797.190 3332.920 ;
        RECT 2796.425 3332.735 2796.715 3332.780 ;
        RECT 2796.870 3332.720 2797.190 3332.780 ;
        RECT 2795.950 3284.300 2796.270 3284.360 ;
        RECT 2795.755 3284.160 2796.270 3284.300 ;
        RECT 2795.950 3284.100 2796.270 3284.160 ;
        RECT 2795.965 3236.360 2796.255 3236.405 ;
        RECT 2796.410 3236.360 2796.730 3236.420 ;
        RECT 2795.965 3236.220 2796.730 3236.360 ;
        RECT 2795.965 3236.175 2796.255 3236.220 ;
        RECT 2796.410 3236.160 2796.730 3236.220 ;
        RECT 1747.150 3218.680 1747.470 3218.740 ;
        RECT 2796.410 3218.680 2796.730 3218.740 ;
        RECT 1747.150 3218.540 2796.730 3218.680 ;
        RECT 1747.150 3218.480 1747.470 3218.540 ;
        RECT 2796.410 3218.480 2796.730 3218.540 ;
      LAYER via ;
        RECT 2795.520 3442.880 2795.780 3443.140 ;
        RECT 2798.280 3442.880 2798.540 3443.140 ;
        RECT 2795.060 3422.140 2795.320 3422.400 ;
        RECT 2796.900 3332.720 2797.160 3332.980 ;
        RECT 2795.980 3284.100 2796.240 3284.360 ;
        RECT 2796.440 3236.160 2796.700 3236.420 ;
        RECT 1747.180 3218.480 1747.440 3218.740 ;
        RECT 2796.440 3218.480 2796.700 3218.740 ;
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
        RECT 2798.340 3443.170 2798.480 3517.600 ;
        RECT 2795.520 3442.850 2795.780 3443.170 ;
        RECT 2798.280 3442.850 2798.540 3443.170 ;
        RECT 2795.580 3429.650 2795.720 3442.850 ;
        RECT 2795.120 3429.510 2795.720 3429.650 ;
        RECT 2795.120 3422.430 2795.260 3429.510 ;
        RECT 2795.060 3422.110 2795.320 3422.430 ;
        RECT 2796.900 3332.690 2797.160 3333.010 ;
        RECT 2796.960 3298.410 2797.100 3332.690 ;
        RECT 2796.040 3298.270 2797.100 3298.410 ;
        RECT 2796.040 3284.390 2796.180 3298.270 ;
        RECT 2795.980 3284.070 2796.240 3284.390 ;
        RECT 2796.440 3236.130 2796.700 3236.450 ;
        RECT 2796.500 3218.770 2796.640 3236.130 ;
        RECT 1747.180 3218.450 1747.440 3218.770 ;
        RECT 2796.440 3218.450 2796.700 3218.770 ;
        RECT 1747.240 3200.000 1747.380 3218.450 ;
        RECT 1747.100 3196.000 1747.380 3200.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2470.345 3332.765 2470.515 3380.875 ;
      LAYER mcon ;
        RECT 2470.345 3380.705 2470.515 3380.875 ;
      LAYER met1 ;
        RECT 2470.270 3380.860 2470.590 3380.920 ;
        RECT 2470.075 3380.720 2470.590 3380.860 ;
        RECT 2470.270 3380.660 2470.590 3380.720 ;
        RECT 2470.285 3332.920 2470.575 3332.965 ;
        RECT 2470.730 3332.920 2471.050 3332.980 ;
        RECT 2470.285 3332.780 2471.050 3332.920 ;
        RECT 2470.285 3332.735 2470.575 3332.780 ;
        RECT 2470.730 3332.720 2471.050 3332.780 ;
        RECT 2470.270 3270.700 2470.590 3270.760 ;
        RECT 2471.190 3270.700 2471.510 3270.760 ;
        RECT 2470.270 3270.560 2471.510 3270.700 ;
        RECT 2470.270 3270.500 2470.590 3270.560 ;
        RECT 2471.190 3270.500 2471.510 3270.560 ;
        RECT 1786.710 3219.360 1787.030 3219.420 ;
        RECT 2471.190 3219.360 2471.510 3219.420 ;
        RECT 1786.710 3219.220 2471.510 3219.360 ;
        RECT 1786.710 3219.160 1787.030 3219.220 ;
        RECT 2471.190 3219.160 2471.510 3219.220 ;
      LAYER via ;
        RECT 2470.300 3380.660 2470.560 3380.920 ;
        RECT 2470.760 3332.720 2471.020 3332.980 ;
        RECT 2470.300 3270.500 2470.560 3270.760 ;
        RECT 2471.220 3270.500 2471.480 3270.760 ;
        RECT 1786.740 3219.160 1787.000 3219.420 ;
        RECT 2471.220 3219.160 2471.480 3219.420 ;
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
        RECT 2474.040 3517.370 2474.180 3517.600 ;
        RECT 2474.040 3517.230 2474.640 3517.370 ;
        RECT 2474.500 3430.445 2474.640 3517.230 ;
        RECT 2474.430 3430.075 2474.710 3430.445 ;
        RECT 2471.210 3429.395 2471.490 3429.765 ;
        RECT 2471.280 3394.970 2471.420 3429.395 ;
        RECT 2470.360 3394.830 2471.420 3394.970 ;
        RECT 2470.360 3380.950 2470.500 3394.830 ;
        RECT 2470.300 3380.630 2470.560 3380.950 ;
        RECT 2470.760 3332.690 2471.020 3333.010 ;
        RECT 2470.820 3298.410 2470.960 3332.690 ;
        RECT 2470.820 3298.270 2471.420 3298.410 ;
        RECT 2471.280 3270.790 2471.420 3298.270 ;
        RECT 2470.300 3270.530 2470.560 3270.790 ;
        RECT 2471.220 3270.530 2471.480 3270.790 ;
        RECT 2470.300 3270.470 2471.480 3270.530 ;
        RECT 2470.360 3270.390 2471.420 3270.470 ;
        RECT 2471.280 3219.450 2471.420 3270.390 ;
        RECT 1786.740 3219.130 1787.000 3219.450 ;
        RECT 2471.220 3219.130 2471.480 3219.450 ;
        RECT 1786.800 3200.000 1786.940 3219.130 ;
        RECT 1786.660 3196.000 1786.940 3200.000 ;
      LAYER via2 ;
        RECT 2474.430 3430.120 2474.710 3430.400 ;
        RECT 2471.210 3429.440 2471.490 3429.720 ;
      LAYER met3 ;
        RECT 2474.405 3430.410 2474.735 3430.425 ;
        RECT 2470.510 3430.110 2474.735 3430.410 ;
        RECT 2470.510 3429.730 2470.810 3430.110 ;
        RECT 2474.405 3430.095 2474.735 3430.110 ;
        RECT 2471.185 3429.730 2471.515 3429.745 ;
        RECT 2470.510 3429.430 2471.515 3429.730 ;
        RECT 2471.185 3429.415 2471.515 3429.430 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2147.885 3332.765 2148.055 3422.355 ;
        RECT 2147.425 3236.205 2147.595 3284.315 ;
      LAYER mcon ;
        RECT 2147.885 3422.185 2148.055 3422.355 ;
        RECT 2147.425 3284.145 2147.595 3284.315 ;
      LAYER met1 ;
        RECT 2146.890 3443.080 2147.210 3443.140 ;
        RECT 2149.190 3443.080 2149.510 3443.140 ;
        RECT 2146.890 3442.940 2149.510 3443.080 ;
        RECT 2146.890 3442.880 2147.210 3442.940 ;
        RECT 2149.190 3442.880 2149.510 3442.940 ;
        RECT 2146.430 3422.340 2146.750 3422.400 ;
        RECT 2147.825 3422.340 2148.115 3422.385 ;
        RECT 2146.430 3422.200 2148.115 3422.340 ;
        RECT 2146.430 3422.140 2146.750 3422.200 ;
        RECT 2147.825 3422.155 2148.115 3422.200 ;
        RECT 2147.825 3332.920 2148.115 3332.965 ;
        RECT 2148.270 3332.920 2148.590 3332.980 ;
        RECT 2147.825 3332.780 2148.590 3332.920 ;
        RECT 2147.825 3332.735 2148.115 3332.780 ;
        RECT 2148.270 3332.720 2148.590 3332.780 ;
        RECT 2147.350 3284.300 2147.670 3284.360 ;
        RECT 2147.155 3284.160 2147.670 3284.300 ;
        RECT 2147.350 3284.100 2147.670 3284.160 ;
        RECT 2147.365 3236.360 2147.655 3236.405 ;
        RECT 2147.810 3236.360 2148.130 3236.420 ;
        RECT 2147.365 3236.220 2148.130 3236.360 ;
        RECT 2147.365 3236.175 2147.655 3236.220 ;
        RECT 2147.810 3236.160 2148.130 3236.220 ;
        RECT 1825.810 3220.040 1826.130 3220.100 ;
        RECT 2147.810 3220.040 2148.130 3220.100 ;
        RECT 1825.810 3219.900 2148.130 3220.040 ;
        RECT 1825.810 3219.840 1826.130 3219.900 ;
        RECT 2147.810 3219.840 2148.130 3219.900 ;
      LAYER via ;
        RECT 2146.920 3442.880 2147.180 3443.140 ;
        RECT 2149.220 3442.880 2149.480 3443.140 ;
        RECT 2146.460 3422.140 2146.720 3422.400 ;
        RECT 2148.300 3332.720 2148.560 3332.980 ;
        RECT 2147.380 3284.100 2147.640 3284.360 ;
        RECT 2147.840 3236.160 2148.100 3236.420 ;
        RECT 1825.840 3219.840 1826.100 3220.100 ;
        RECT 2147.840 3219.840 2148.100 3220.100 ;
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
        RECT 2149.280 3443.170 2149.420 3517.600 ;
        RECT 2146.920 3442.850 2147.180 3443.170 ;
        RECT 2149.220 3442.850 2149.480 3443.170 ;
        RECT 2146.980 3429.650 2147.120 3442.850 ;
        RECT 2146.520 3429.510 2147.120 3429.650 ;
        RECT 2146.520 3422.430 2146.660 3429.510 ;
        RECT 2146.460 3422.110 2146.720 3422.430 ;
        RECT 2148.300 3332.690 2148.560 3333.010 ;
        RECT 2148.360 3298.410 2148.500 3332.690 ;
        RECT 2147.440 3298.270 2148.500 3298.410 ;
        RECT 2147.440 3284.390 2147.580 3298.270 ;
        RECT 2147.380 3284.070 2147.640 3284.390 ;
        RECT 2147.840 3236.130 2148.100 3236.450 ;
        RECT 2147.900 3220.130 2148.040 3236.130 ;
        RECT 1825.840 3219.810 1826.100 3220.130 ;
        RECT 2147.840 3219.810 2148.100 3220.130 ;
        RECT 1825.900 3200.000 1826.040 3219.810 ;
        RECT 1825.760 3196.000 1826.040 3200.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1824.890 3498.500 1825.210 3498.560 ;
        RECT 1828.110 3498.500 1828.430 3498.560 ;
        RECT 1824.890 3498.360 1828.430 3498.500 ;
        RECT 1824.890 3498.300 1825.210 3498.360 ;
        RECT 1828.110 3498.300 1828.430 3498.360 ;
        RECT 1828.110 3215.620 1828.430 3215.680 ;
        RECT 1865.370 3215.620 1865.690 3215.680 ;
        RECT 1828.110 3215.480 1865.690 3215.620 ;
        RECT 1828.110 3215.420 1828.430 3215.480 ;
        RECT 1865.370 3215.420 1865.690 3215.480 ;
      LAYER via ;
        RECT 1824.920 3498.300 1825.180 3498.560 ;
        RECT 1828.140 3498.300 1828.400 3498.560 ;
        RECT 1828.140 3215.420 1828.400 3215.680 ;
        RECT 1865.400 3215.420 1865.660 3215.680 ;
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
        RECT 1824.980 3498.590 1825.120 3517.600 ;
        RECT 1824.920 3498.270 1825.180 3498.590 ;
        RECT 1828.140 3498.270 1828.400 3498.590 ;
        RECT 1828.200 3215.710 1828.340 3498.270 ;
        RECT 1828.140 3215.390 1828.400 3215.710 ;
        RECT 1865.400 3215.390 1865.660 3215.710 ;
        RECT 1865.460 3200.000 1865.600 3215.390 ;
        RECT 1865.320 3196.000 1865.600 3200.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1500.590 3498.500 1500.910 3498.560 ;
        RECT 1503.810 3498.500 1504.130 3498.560 ;
        RECT 1500.590 3498.360 1504.130 3498.500 ;
        RECT 1500.590 3498.300 1500.910 3498.360 ;
        RECT 1503.810 3498.300 1504.130 3498.360 ;
        RECT 1503.810 3219.700 1504.130 3219.760 ;
        RECT 1904.930 3219.700 1905.250 3219.760 ;
        RECT 1503.810 3219.560 1905.250 3219.700 ;
        RECT 1503.810 3219.500 1504.130 3219.560 ;
        RECT 1904.930 3219.500 1905.250 3219.560 ;
      LAYER via ;
        RECT 1500.620 3498.300 1500.880 3498.560 ;
        RECT 1503.840 3498.300 1504.100 3498.560 ;
        RECT 1503.840 3219.500 1504.100 3219.760 ;
        RECT 1904.960 3219.500 1905.220 3219.760 ;
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
        RECT 1500.680 3498.590 1500.820 3517.600 ;
        RECT 1500.620 3498.270 1500.880 3498.590 ;
        RECT 1503.840 3498.270 1504.100 3498.590 ;
        RECT 1503.900 3219.790 1504.040 3498.270 ;
        RECT 1503.840 3219.470 1504.100 3219.790 ;
        RECT 1904.960 3219.470 1905.220 3219.790 ;
        RECT 1905.020 3200.000 1905.160 3219.470 ;
        RECT 1904.880 3196.000 1905.160 3200.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1200.210 322.560 1200.530 322.620 ;
        RECT 1241.610 322.560 1241.930 322.620 ;
        RECT 1200.210 322.420 1241.930 322.560 ;
        RECT 1200.210 322.360 1200.530 322.420 ;
        RECT 1241.610 322.360 1241.930 322.420 ;
        RECT 1338.210 319.500 1338.530 319.560 ;
        RECT 1379.610 319.500 1379.930 319.560 ;
        RECT 1338.210 319.360 1379.930 319.500 ;
        RECT 1338.210 319.300 1338.530 319.360 ;
        RECT 1379.610 319.300 1379.930 319.360 ;
        RECT 1777.510 319.160 1777.830 319.220 ;
        RECT 1801.890 319.160 1802.210 319.220 ;
        RECT 1777.510 319.020 1802.210 319.160 ;
        RECT 1777.510 318.960 1777.830 319.020 ;
        RECT 1801.890 318.960 1802.210 319.020 ;
        RECT 1966.570 319.160 1966.890 319.220 ;
        RECT 2028.210 319.160 2028.530 319.220 ;
        RECT 1966.570 319.020 2028.530 319.160 ;
        RECT 1966.570 318.960 1966.890 319.020 ;
        RECT 2028.210 318.960 2028.530 319.020 ;
        RECT 1731.050 318.140 1731.370 318.200 ;
        RECT 1732.430 318.140 1732.750 318.200 ;
        RECT 1731.050 318.000 1732.750 318.140 ;
        RECT 1731.050 317.940 1731.370 318.000 ;
        RECT 1732.430 317.940 1732.750 318.000 ;
        RECT 2608.270 318.140 2608.590 318.200 ;
        RECT 2632.190 318.140 2632.510 318.200 ;
        RECT 2608.270 318.000 2632.510 318.140 ;
        RECT 2608.270 317.940 2608.590 318.000 ;
        RECT 2632.190 317.940 2632.510 318.000 ;
        RECT 1687.350 317.800 1687.670 317.860 ;
        RECT 1724.610 317.800 1724.930 317.860 ;
        RECT 1687.350 317.660 1724.930 317.800 ;
        RECT 1687.350 317.600 1687.670 317.660 ;
        RECT 1724.610 317.600 1724.930 317.660 ;
      LAYER via ;
        RECT 1200.240 322.360 1200.500 322.620 ;
        RECT 1241.640 322.360 1241.900 322.620 ;
        RECT 1338.240 319.300 1338.500 319.560 ;
        RECT 1379.640 319.300 1379.900 319.560 ;
        RECT 1777.540 318.960 1777.800 319.220 ;
        RECT 1801.920 318.960 1802.180 319.220 ;
        RECT 1966.600 318.960 1966.860 319.220 ;
        RECT 2028.240 318.960 2028.500 319.220 ;
        RECT 1731.080 317.940 1731.340 318.200 ;
        RECT 1732.460 317.940 1732.720 318.200 ;
        RECT 2608.300 317.940 2608.560 318.200 ;
        RECT 2632.220 317.940 2632.480 318.200 ;
        RECT 1687.380 317.600 1687.640 317.860 ;
        RECT 1724.640 317.600 1724.900 317.860 ;
      LAYER met2 ;
        RECT 1194.180 3196.410 1194.460 3200.000 ;
        RECT 1195.630 3196.410 1195.910 3196.525 ;
        RECT 1194.180 3196.270 1195.910 3196.410 ;
        RECT 1194.180 3196.000 1194.460 3196.270 ;
        RECT 1195.630 3196.155 1195.910 3196.270 ;
        RECT 1200.230 324.515 1200.510 324.885 ;
        RECT 1200.300 322.650 1200.440 324.515 ;
        RECT 1200.240 322.330 1200.500 322.650 ;
        RECT 1241.640 322.330 1241.900 322.650 ;
        RECT 1241.700 318.085 1241.840 322.330 ;
        RECT 1265.550 321.115 1265.830 321.485 ;
        RECT 1241.630 317.715 1241.910 318.085 ;
        RECT 1265.620 316.725 1265.760 321.115 ;
        RECT 1521.310 320.435 1521.590 320.805 ;
        RECT 1338.240 319.445 1338.500 319.590 ;
        RECT 1379.640 319.445 1379.900 319.590 ;
        RECT 1338.230 319.075 1338.510 319.445 ;
        RECT 1379.630 319.075 1379.910 319.445 ;
        RECT 1386.530 319.075 1386.810 319.445 ;
        RECT 1386.600 318.085 1386.740 319.075 ;
        RECT 1521.380 318.085 1521.520 320.435 ;
        RECT 2704.430 319.755 2704.710 320.125 ;
        RECT 1732.450 319.075 1732.730 319.445 ;
        RECT 1777.530 319.075 1777.810 319.445 ;
        RECT 1732.520 318.230 1732.660 319.075 ;
        RECT 1777.540 318.930 1777.800 319.075 ;
        RECT 1801.920 318.930 1802.180 319.250 ;
        RECT 1966.600 318.930 1966.860 319.250 ;
        RECT 2028.230 319.075 2028.510 319.445 ;
        RECT 2090.330 319.075 2090.610 319.445 ;
        RECT 2028.240 318.930 2028.500 319.075 ;
        RECT 1731.080 318.085 1731.340 318.230 ;
        RECT 1386.530 317.715 1386.810 318.085 ;
        RECT 1521.310 317.715 1521.590 318.085 ;
        RECT 1687.370 317.715 1687.650 318.085 ;
        RECT 1724.630 317.715 1724.910 318.085 ;
        RECT 1731.070 317.715 1731.350 318.085 ;
        RECT 1732.460 317.910 1732.720 318.230 ;
        RECT 1801.980 318.085 1802.120 318.930 ;
        RECT 1966.660 318.765 1966.800 318.930 ;
        RECT 1917.830 318.395 1918.110 318.765 ;
        RECT 1966.590 318.395 1966.870 318.765 ;
        RECT 2090.400 318.650 2090.540 319.075 ;
        RECT 2090.790 318.650 2091.070 318.765 ;
        RECT 2090.400 318.510 2091.070 318.650 ;
        RECT 2090.790 318.395 2091.070 318.510 ;
        RECT 2283.530 318.650 2283.810 318.765 ;
        RECT 2284.450 318.650 2284.730 318.765 ;
        RECT 2283.530 318.510 2284.730 318.650 ;
        RECT 2283.530 318.395 2283.810 318.510 ;
        RECT 2284.450 318.395 2284.730 318.510 ;
        RECT 2572.870 318.395 2573.150 318.765 ;
        RECT 2632.210 318.395 2632.490 318.765 ;
        RECT 1801.910 317.715 1802.190 318.085 ;
        RECT 1687.380 317.570 1687.640 317.715 ;
        RECT 1724.640 317.570 1724.900 317.715 ;
        RECT 1917.900 317.405 1918.040 318.395 ;
        RECT 1917.830 317.035 1918.110 317.405 ;
        RECT 2572.940 316.725 2573.080 318.395 ;
        RECT 2632.280 318.230 2632.420 318.395 ;
        RECT 2608.300 318.085 2608.560 318.230 ;
        RECT 2608.290 317.715 2608.570 318.085 ;
        RECT 2632.220 317.910 2632.480 318.230 ;
        RECT 2704.500 318.085 2704.640 319.755 ;
        RECT 2801.030 319.075 2801.310 319.445 ;
        RECT 2704.430 317.715 2704.710 318.085 ;
        RECT 2801.100 317.405 2801.240 319.075 ;
        RECT 2863.130 318.395 2863.410 318.765 ;
        RECT 2863.200 317.970 2863.340 318.395 ;
        RECT 2863.590 317.970 2863.870 318.085 ;
        RECT 2863.200 317.830 2863.870 317.970 ;
        RECT 2863.590 317.715 2863.870 317.830 ;
        RECT 2801.030 317.035 2801.310 317.405 ;
        RECT 1265.550 316.355 1265.830 316.725 ;
        RECT 2572.870 316.355 2573.150 316.725 ;
      LAYER via2 ;
        RECT 1195.630 3196.200 1195.910 3196.480 ;
        RECT 1200.230 324.560 1200.510 324.840 ;
        RECT 1265.550 321.160 1265.830 321.440 ;
        RECT 1241.630 317.760 1241.910 318.040 ;
        RECT 1521.310 320.480 1521.590 320.760 ;
        RECT 1338.230 319.120 1338.510 319.400 ;
        RECT 1379.630 319.120 1379.910 319.400 ;
        RECT 1386.530 319.120 1386.810 319.400 ;
        RECT 2704.430 319.800 2704.710 320.080 ;
        RECT 1732.450 319.120 1732.730 319.400 ;
        RECT 1777.530 319.120 1777.810 319.400 ;
        RECT 2028.230 319.120 2028.510 319.400 ;
        RECT 2090.330 319.120 2090.610 319.400 ;
        RECT 1386.530 317.760 1386.810 318.040 ;
        RECT 1521.310 317.760 1521.590 318.040 ;
        RECT 1687.370 317.760 1687.650 318.040 ;
        RECT 1724.630 317.760 1724.910 318.040 ;
        RECT 1731.070 317.760 1731.350 318.040 ;
        RECT 1917.830 318.440 1918.110 318.720 ;
        RECT 1966.590 318.440 1966.870 318.720 ;
        RECT 2090.790 318.440 2091.070 318.720 ;
        RECT 2283.530 318.440 2283.810 318.720 ;
        RECT 2284.450 318.440 2284.730 318.720 ;
        RECT 2572.870 318.440 2573.150 318.720 ;
        RECT 2632.210 318.440 2632.490 318.720 ;
        RECT 1801.910 317.760 1802.190 318.040 ;
        RECT 1917.830 317.080 1918.110 317.360 ;
        RECT 2608.290 317.760 2608.570 318.040 ;
        RECT 2801.030 319.120 2801.310 319.400 ;
        RECT 2704.430 317.760 2704.710 318.040 ;
        RECT 2863.130 318.440 2863.410 318.720 ;
        RECT 2863.590 317.760 2863.870 318.040 ;
        RECT 2801.030 317.080 2801.310 317.360 ;
        RECT 1265.550 316.400 1265.830 316.680 ;
        RECT 2572.870 316.400 2573.150 316.680 ;
      LAYER met3 ;
        RECT 1195.605 3196.490 1195.935 3196.505 ;
        RECT 1199.950 3196.490 1200.330 3196.500 ;
        RECT 1195.605 3196.190 1200.330 3196.490 ;
        RECT 1195.605 3196.175 1195.935 3196.190 ;
        RECT 1199.950 3196.180 1200.330 3196.190 ;
        RECT 1200.205 324.860 1200.535 324.865 ;
        RECT 1199.950 324.850 1200.535 324.860 ;
        RECT 1199.750 324.550 1200.535 324.850 ;
        RECT 1199.950 324.540 1200.535 324.550 ;
        RECT 1200.205 324.535 1200.535 324.540 ;
        RECT 2917.600 322.810 2924.800 323.260 ;
        RECT 2916.710 322.510 2924.800 322.810 ;
        RECT 1265.525 321.450 1265.855 321.465 ;
        RECT 1265.525 321.150 1290.450 321.450 ;
        RECT 1265.525 321.135 1265.855 321.150 ;
        RECT 1290.150 320.770 1290.450 321.150 ;
        RECT 1521.285 320.770 1521.615 320.785 ;
        RECT 1290.150 320.470 1318.050 320.770 ;
        RECT 1317.750 319.410 1318.050 320.470 ;
        RECT 1497.150 320.470 1521.615 320.770 ;
        RECT 1338.205 319.410 1338.535 319.425 ;
        RECT 1317.750 319.110 1338.535 319.410 ;
        RECT 1338.205 319.095 1338.535 319.110 ;
        RECT 1379.605 319.410 1379.935 319.425 ;
        RECT 1386.505 319.410 1386.835 319.425 ;
        RECT 1497.150 319.410 1497.450 320.470 ;
        RECT 1521.285 320.455 1521.615 320.470 ;
        RECT 2510.030 320.090 2510.410 320.100 ;
        RECT 2476.030 319.790 2510.410 320.090 ;
        RECT 1379.605 319.110 1386.835 319.410 ;
        RECT 1379.605 319.095 1379.935 319.110 ;
        RECT 1386.505 319.095 1386.835 319.110 ;
        RECT 1434.590 319.110 1497.450 319.410 ;
        RECT 1732.425 319.410 1732.755 319.425 ;
        RECT 1777.505 319.410 1777.835 319.425 ;
        RECT 1732.425 319.110 1777.835 319.410 ;
        RECT 1434.590 318.730 1434.890 319.110 ;
        RECT 1732.425 319.095 1732.755 319.110 ;
        RECT 1777.505 319.095 1777.835 319.110 ;
        RECT 2028.205 319.410 2028.535 319.425 ;
        RECT 2090.305 319.410 2090.635 319.425 ;
        RECT 2028.205 319.110 2042.090 319.410 ;
        RECT 2028.205 319.095 2028.535 319.110 ;
        RECT 1869.710 318.730 1870.090 318.740 ;
        RECT 1386.750 318.430 1434.890 318.730 ;
        RECT 1821.910 318.430 1870.090 318.730 ;
        RECT 1386.750 318.065 1387.050 318.430 ;
        RECT 1241.605 318.050 1241.935 318.065 ;
        RECT 1241.605 317.750 1242.610 318.050 ;
        RECT 1241.605 317.735 1241.935 317.750 ;
        RECT 1242.310 316.690 1242.610 317.750 ;
        RECT 1386.505 317.750 1387.050 318.065 ;
        RECT 1521.285 318.050 1521.615 318.065 ;
        RECT 1545.870 318.050 1546.250 318.060 ;
        RECT 1687.345 318.050 1687.675 318.065 ;
        RECT 1521.285 317.750 1546.250 318.050 ;
        RECT 1386.505 317.735 1386.835 317.750 ;
        RECT 1521.285 317.735 1521.615 317.750 ;
        RECT 1545.870 317.740 1546.250 317.750 ;
        RECT 1651.710 317.750 1687.675 318.050 ;
        RECT 1265.525 316.690 1265.855 316.705 ;
        RECT 1242.310 316.390 1265.855 316.690 ;
        RECT 1265.525 316.375 1265.855 316.390 ;
        RECT 1545.870 316.690 1546.250 316.700 ;
        RECT 1651.710 316.690 1652.010 317.750 ;
        RECT 1687.345 317.735 1687.675 317.750 ;
        RECT 1724.605 318.050 1724.935 318.065 ;
        RECT 1731.045 318.050 1731.375 318.065 ;
        RECT 1724.605 317.750 1731.375 318.050 ;
        RECT 1724.605 317.735 1724.935 317.750 ;
        RECT 1731.045 317.735 1731.375 317.750 ;
        RECT 1801.885 318.050 1802.215 318.065 ;
        RECT 1821.910 318.050 1822.210 318.430 ;
        RECT 1869.710 318.420 1870.090 318.430 ;
        RECT 1917.805 318.730 1918.135 318.745 ;
        RECT 1966.565 318.730 1966.895 318.745 ;
        RECT 1917.805 318.430 1966.895 318.730 ;
        RECT 1917.805 318.415 1918.135 318.430 ;
        RECT 1966.565 318.415 1966.895 318.430 ;
        RECT 1801.885 317.750 1822.210 318.050 ;
        RECT 2041.790 318.050 2042.090 319.110 ;
        RECT 2076.750 319.110 2090.635 319.410 ;
        RECT 2076.750 318.730 2077.050 319.110 ;
        RECT 2090.305 319.095 2090.635 319.110 ;
        RECT 2124.590 319.110 2138.690 319.410 ;
        RECT 2042.710 318.430 2077.050 318.730 ;
        RECT 2090.765 318.730 2091.095 318.745 ;
        RECT 2124.590 318.730 2124.890 319.110 ;
        RECT 2090.765 318.430 2124.890 318.730 ;
        RECT 2042.710 318.050 2043.010 318.430 ;
        RECT 2090.765 318.415 2091.095 318.430 ;
        RECT 2041.790 317.750 2043.010 318.050 ;
        RECT 2138.390 318.050 2138.690 319.110 ;
        RECT 2139.310 319.110 2187.450 319.410 ;
        RECT 2139.310 318.050 2139.610 319.110 ;
        RECT 2138.390 317.750 2139.610 318.050 ;
        RECT 2187.150 318.050 2187.450 319.110 ;
        RECT 2283.505 318.730 2283.835 318.745 ;
        RECT 2235.910 318.430 2283.835 318.730 ;
        RECT 2235.910 318.050 2236.210 318.430 ;
        RECT 2283.505 318.415 2283.835 318.430 ;
        RECT 2284.425 318.730 2284.755 318.745 ;
        RECT 2476.030 318.730 2476.330 319.790 ;
        RECT 2510.030 319.780 2510.410 319.790 ;
        RECT 2656.310 320.090 2656.690 320.100 ;
        RECT 2704.405 320.090 2704.735 320.105 ;
        RECT 2656.310 319.790 2704.735 320.090 ;
        RECT 2656.310 319.780 2656.690 319.790 ;
        RECT 2704.405 319.775 2704.735 319.790 ;
        RECT 2801.005 319.410 2801.335 319.425 ;
        RECT 2801.005 319.110 2815.810 319.410 ;
        RECT 2801.005 319.095 2801.335 319.110 ;
        RECT 2572.845 318.730 2573.175 318.745 ;
        RECT 2284.425 318.430 2331.890 318.730 ;
        RECT 2284.425 318.415 2284.755 318.430 ;
        RECT 2187.150 317.750 2236.210 318.050 ;
        RECT 2331.590 318.050 2331.890 318.430 ;
        RECT 2332.510 318.430 2414.690 318.730 ;
        RECT 2332.510 318.050 2332.810 318.430 ;
        RECT 2331.590 317.750 2332.810 318.050 ;
        RECT 2414.390 318.050 2414.690 318.430 ;
        RECT 2429.110 318.430 2476.330 318.730 ;
        RECT 2525.710 318.430 2573.175 318.730 ;
        RECT 2429.110 318.050 2429.410 318.430 ;
        RECT 2414.390 317.750 2429.410 318.050 ;
        RECT 2510.950 318.050 2511.330 318.060 ;
        RECT 2525.710 318.050 2526.010 318.430 ;
        RECT 2572.845 318.415 2573.175 318.430 ;
        RECT 2632.185 318.730 2632.515 318.745 ;
        RECT 2656.310 318.730 2656.690 318.740 ;
        RECT 2752.910 318.730 2753.290 318.740 ;
        RECT 2632.185 318.430 2656.690 318.730 ;
        RECT 2632.185 318.415 2632.515 318.430 ;
        RECT 2656.310 318.420 2656.690 318.430 ;
        RECT 2718.910 318.430 2753.290 318.730 ;
        RECT 2608.265 318.050 2608.595 318.065 ;
        RECT 2510.950 317.750 2526.010 318.050 ;
        RECT 2607.590 317.750 2608.595 318.050 ;
        RECT 1801.885 317.735 1802.215 317.750 ;
        RECT 2510.950 317.740 2511.330 317.750 ;
        RECT 1869.710 317.370 1870.090 317.380 ;
        RECT 1917.805 317.370 1918.135 317.385 ;
        RECT 1869.710 317.070 1918.135 317.370 ;
        RECT 1869.710 317.060 1870.090 317.070 ;
        RECT 1917.805 317.055 1918.135 317.070 ;
        RECT 1545.870 316.390 1652.010 316.690 ;
        RECT 2572.845 316.690 2573.175 316.705 ;
        RECT 2607.590 316.690 2607.890 317.750 ;
        RECT 2608.265 317.735 2608.595 317.750 ;
        RECT 2704.405 318.050 2704.735 318.065 ;
        RECT 2718.910 318.050 2719.210 318.430 ;
        RECT 2752.910 318.420 2753.290 318.430 ;
        RECT 2704.405 317.750 2719.210 318.050 ;
        RECT 2815.510 318.050 2815.810 319.110 ;
        RECT 2863.105 318.730 2863.435 318.745 ;
        RECT 2916.710 318.730 2917.010 322.510 ;
        RECT 2917.600 322.060 2924.800 322.510 ;
        RECT 2849.550 318.430 2863.435 318.730 ;
        RECT 2849.550 318.050 2849.850 318.430 ;
        RECT 2863.105 318.415 2863.435 318.430 ;
        RECT 2884.510 318.430 2917.010 318.730 ;
        RECT 2815.510 317.750 2849.850 318.050 ;
        RECT 2863.565 318.050 2863.895 318.065 ;
        RECT 2884.510 318.050 2884.810 318.430 ;
        RECT 2863.565 317.750 2884.810 318.050 ;
        RECT 2704.405 317.735 2704.735 317.750 ;
        RECT 2863.565 317.735 2863.895 317.750 ;
        RECT 2752.910 317.370 2753.290 317.380 ;
        RECT 2801.005 317.370 2801.335 317.385 ;
        RECT 2752.910 317.070 2801.335 317.370 ;
        RECT 2752.910 317.060 2753.290 317.070 ;
        RECT 2801.005 317.055 2801.335 317.070 ;
        RECT 2572.845 316.390 2607.890 316.690 ;
        RECT 1545.870 316.380 1546.250 316.390 ;
        RECT 2572.845 316.375 2573.175 316.390 ;
      LAYER via3 ;
        RECT 1199.980 3196.180 1200.300 3196.500 ;
        RECT 1199.980 324.540 1200.300 324.860 ;
        RECT 1545.900 317.740 1546.220 318.060 ;
        RECT 1545.900 316.380 1546.220 316.700 ;
        RECT 1869.740 318.420 1870.060 318.740 ;
        RECT 2510.060 319.780 2510.380 320.100 ;
        RECT 2656.340 319.780 2656.660 320.100 ;
        RECT 2510.980 317.740 2511.300 318.060 ;
        RECT 2656.340 318.420 2656.660 318.740 ;
        RECT 1869.740 317.060 1870.060 317.380 ;
        RECT 2752.940 318.420 2753.260 318.740 ;
        RECT 2752.940 317.060 2753.260 317.380 ;
      LAYER met4 ;
        RECT 1199.975 3196.175 1200.305 3196.505 ;
        RECT 1199.990 324.865 1200.290 3196.175 ;
        RECT 1199.975 324.535 1200.305 324.865 ;
        RECT 2510.055 319.775 2510.385 320.105 ;
        RECT 2656.335 319.775 2656.665 320.105 ;
        RECT 1869.735 318.415 1870.065 318.745 ;
        RECT 1545.895 317.735 1546.225 318.065 ;
        RECT 1545.910 316.705 1546.210 317.735 ;
        RECT 1869.750 317.385 1870.050 318.415 ;
        RECT 2510.070 318.050 2510.370 319.775 ;
        RECT 2656.350 318.745 2656.650 319.775 ;
        RECT 2656.335 318.415 2656.665 318.745 ;
        RECT 2752.935 318.415 2753.265 318.745 ;
        RECT 2510.975 318.050 2511.305 318.065 ;
        RECT 2510.070 317.750 2511.305 318.050 ;
        RECT 2510.975 317.735 2511.305 317.750 ;
        RECT 2752.950 317.385 2753.250 318.415 ;
        RECT 1869.735 317.055 1870.065 317.385 ;
        RECT 2752.935 317.055 2753.265 317.385 ;
        RECT 1545.895 316.375 1546.225 316.705 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1175.830 3498.500 1176.150 3498.560 ;
        RECT 1179.510 3498.500 1179.830 3498.560 ;
        RECT 1175.830 3498.360 1179.830 3498.500 ;
        RECT 1175.830 3498.300 1176.150 3498.360 ;
        RECT 1179.510 3498.300 1179.830 3498.360 ;
        RECT 1179.510 3219.020 1179.830 3219.080 ;
        RECT 1944.490 3219.020 1944.810 3219.080 ;
        RECT 1179.510 3218.880 1944.810 3219.020 ;
        RECT 1179.510 3218.820 1179.830 3218.880 ;
        RECT 1944.490 3218.820 1944.810 3218.880 ;
      LAYER via ;
        RECT 1175.860 3498.300 1176.120 3498.560 ;
        RECT 1179.540 3498.300 1179.800 3498.560 ;
        RECT 1179.540 3218.820 1179.800 3219.080 ;
        RECT 1944.520 3218.820 1944.780 3219.080 ;
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
        RECT 1175.920 3498.590 1176.060 3517.600 ;
        RECT 1175.860 3498.270 1176.120 3498.590 ;
        RECT 1179.540 3498.270 1179.800 3498.590 ;
        RECT 1179.600 3219.110 1179.740 3498.270 ;
        RECT 1179.540 3218.790 1179.800 3219.110 ;
        RECT 1944.520 3218.790 1944.780 3219.110 ;
        RECT 1944.580 3200.000 1944.720 3218.790 ;
        RECT 1944.440 3196.000 1944.720 3200.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 851.530 3503.940 851.850 3504.000 ;
        RECT 1980.370 3503.940 1980.690 3504.000 ;
        RECT 851.530 3503.800 1980.690 3503.940 ;
        RECT 851.530 3503.740 851.850 3503.800 ;
        RECT 1980.370 3503.740 1980.690 3503.800 ;
      LAYER via ;
        RECT 851.560 3503.740 851.820 3504.000 ;
        RECT 1980.400 3503.740 1980.660 3504.000 ;
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
        RECT 851.620 3504.030 851.760 3517.600 ;
        RECT 851.560 3503.710 851.820 3504.030 ;
        RECT 1980.400 3503.710 1980.660 3504.030 ;
        RECT 1980.460 3199.810 1980.600 3503.710 ;
        RECT 1984.000 3199.810 1984.280 3200.000 ;
        RECT 1980.460 3199.670 1984.280 3199.810 ;
        RECT 1984.000 3196.000 1984.280 3199.670 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 527.230 3502.920 527.550 3502.980 ;
        RECT 2021.770 3502.920 2022.090 3502.980 ;
        RECT 527.230 3502.780 2022.090 3502.920 ;
        RECT 527.230 3502.720 527.550 3502.780 ;
        RECT 2021.770 3502.720 2022.090 3502.780 ;
      LAYER via ;
        RECT 527.260 3502.720 527.520 3502.980 ;
        RECT 2021.800 3502.720 2022.060 3502.980 ;
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
        RECT 527.320 3503.010 527.460 3517.600 ;
        RECT 527.260 3502.690 527.520 3503.010 ;
        RECT 2021.800 3502.690 2022.060 3503.010 ;
        RECT 2021.860 3199.810 2022.000 3502.690 ;
        RECT 2023.100 3199.810 2023.380 3200.000 ;
        RECT 2021.860 3199.670 2023.380 3199.810 ;
        RECT 2023.100 3196.000 2023.380 3199.670 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 202.470 3501.900 202.790 3501.960 ;
        RECT 2056.270 3501.900 2056.590 3501.960 ;
        RECT 202.470 3501.760 2056.590 3501.900 ;
        RECT 202.470 3501.700 202.790 3501.760 ;
        RECT 2056.270 3501.700 2056.590 3501.760 ;
      LAYER via ;
        RECT 202.500 3501.700 202.760 3501.960 ;
        RECT 2056.300 3501.700 2056.560 3501.960 ;
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
        RECT 202.560 3501.990 202.700 3517.600 ;
        RECT 202.500 3501.670 202.760 3501.990 ;
        RECT 2056.300 3501.670 2056.560 3501.990 ;
        RECT 2056.360 3199.130 2056.500 3501.670 ;
        RECT 2062.660 3199.130 2062.940 3200.000 ;
        RECT 2056.360 3198.990 2062.940 3199.130 ;
        RECT 2062.660 3196.000 2062.940 3198.990 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.550 3408.740 17.870 3408.800 ;
        RECT 2097.670 3408.740 2097.990 3408.800 ;
        RECT 17.550 3408.600 2097.990 3408.740 ;
        RECT 17.550 3408.540 17.870 3408.600 ;
        RECT 2097.670 3408.540 2097.990 3408.600 ;
      LAYER via ;
        RECT 17.580 3408.540 17.840 3408.800 ;
        RECT 2097.700 3408.540 2097.960 3408.800 ;
      LAYER met2 ;
        RECT 17.570 3411.035 17.850 3411.405 ;
        RECT 17.640 3408.830 17.780 3411.035 ;
        RECT 17.580 3408.510 17.840 3408.830 ;
        RECT 2097.700 3408.510 2097.960 3408.830 ;
        RECT 2097.760 3199.130 2097.900 3408.510 ;
        RECT 2102.220 3199.130 2102.500 3200.000 ;
        RECT 2097.760 3198.990 2102.500 3199.130 ;
        RECT 2102.220 3196.000 2102.500 3198.990 ;
      LAYER via2 ;
        RECT 17.570 3411.080 17.850 3411.360 ;
      LAYER met3 ;
        RECT -4.800 3411.370 2.400 3411.820 ;
        RECT 17.545 3411.370 17.875 3411.385 ;
        RECT -4.800 3411.070 17.875 3411.370 ;
        RECT -4.800 3410.620 2.400 3411.070 ;
        RECT 17.545 3411.055 17.875 3411.070 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2140.525 3196.085 2140.695 3199.655 ;
      LAYER mcon ;
        RECT 2140.525 3199.485 2140.695 3199.655 ;
      LAYER met1 ;
        RECT 2140.450 3199.640 2140.770 3199.700 ;
        RECT 2140.255 3199.500 2140.770 3199.640 ;
        RECT 2140.450 3199.440 2140.770 3199.500 ;
        RECT 33.650 3196.240 33.970 3196.300 ;
        RECT 2140.465 3196.240 2140.755 3196.285 ;
        RECT 33.650 3196.100 2140.755 3196.240 ;
        RECT 33.650 3196.040 33.970 3196.100 ;
        RECT 2140.465 3196.055 2140.755 3196.100 ;
        RECT 15.710 3124.840 16.030 3124.900 ;
        RECT 33.650 3124.840 33.970 3124.900 ;
        RECT 15.710 3124.700 33.970 3124.840 ;
        RECT 15.710 3124.640 16.030 3124.700 ;
        RECT 33.650 3124.640 33.970 3124.700 ;
      LAYER via ;
        RECT 2140.480 3199.440 2140.740 3199.700 ;
        RECT 33.680 3196.040 33.940 3196.300 ;
        RECT 15.740 3124.640 16.000 3124.900 ;
        RECT 33.680 3124.640 33.940 3124.900 ;
      LAYER met2 ;
        RECT 2141.780 3199.810 2142.060 3200.000 ;
        RECT 2140.540 3199.730 2142.060 3199.810 ;
        RECT 2140.480 3199.670 2142.060 3199.730 ;
        RECT 2140.480 3199.410 2140.740 3199.670 ;
        RECT 33.680 3196.010 33.940 3196.330 ;
        RECT 33.740 3124.930 33.880 3196.010 ;
        RECT 2141.780 3196.000 2142.060 3199.670 ;
        RECT 15.740 3124.610 16.000 3124.930 ;
        RECT 33.680 3124.610 33.940 3124.930 ;
        RECT 15.800 3124.445 15.940 3124.610 ;
        RECT 15.730 3124.075 16.010 3124.445 ;
      LAYER via2 ;
        RECT 15.730 3124.120 16.010 3124.400 ;
      LAYER met3 ;
        RECT -4.800 3124.410 2.400 3124.860 ;
        RECT 15.705 3124.410 16.035 3124.425 ;
        RECT -4.800 3124.110 16.035 3124.410 ;
        RECT -4.800 3123.660 2.400 3124.110 ;
        RECT 15.705 3124.095 16.035 3124.110 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2180.545 3195.745 2180.715 3199.655 ;
      LAYER mcon ;
        RECT 2180.545 3199.485 2180.715 3199.655 ;
      LAYER met1 ;
        RECT 2180.470 3199.640 2180.790 3199.700 ;
        RECT 2180.275 3199.500 2180.790 3199.640 ;
        RECT 2180.470 3199.440 2180.790 3199.500 ;
        RECT 33.190 3195.900 33.510 3195.960 ;
        RECT 2180.485 3195.900 2180.775 3195.945 ;
        RECT 33.190 3195.760 2180.775 3195.900 ;
        RECT 33.190 3195.700 33.510 3195.760 ;
        RECT 2180.485 3195.715 2180.775 3195.760 ;
        RECT 15.710 2837.880 16.030 2837.940 ;
        RECT 33.190 2837.880 33.510 2837.940 ;
        RECT 15.710 2837.740 33.510 2837.880 ;
        RECT 15.710 2837.680 16.030 2837.740 ;
        RECT 33.190 2837.680 33.510 2837.740 ;
      LAYER via ;
        RECT 2180.500 3199.440 2180.760 3199.700 ;
        RECT 33.220 3195.700 33.480 3195.960 ;
        RECT 15.740 2837.680 16.000 2837.940 ;
        RECT 33.220 2837.680 33.480 2837.940 ;
      LAYER met2 ;
        RECT 2181.340 3199.810 2181.620 3200.000 ;
        RECT 2180.560 3199.730 2181.620 3199.810 ;
        RECT 2180.500 3199.670 2181.620 3199.730 ;
        RECT 2180.500 3199.410 2180.760 3199.670 ;
        RECT 2181.340 3196.000 2181.620 3199.670 ;
        RECT 33.220 3195.670 33.480 3195.990 ;
        RECT 33.280 2837.970 33.420 3195.670 ;
        RECT 15.740 2837.650 16.000 2837.970 ;
        RECT 33.220 2837.650 33.480 2837.970 ;
        RECT 15.800 2836.805 15.940 2837.650 ;
        RECT 15.730 2836.435 16.010 2836.805 ;
      LAYER via2 ;
        RECT 15.730 2836.480 16.010 2836.760 ;
      LAYER met3 ;
        RECT -4.800 2836.770 2.400 2837.220 ;
        RECT 15.705 2836.770 16.035 2836.785 ;
        RECT -4.800 2836.470 16.035 2836.770 ;
        RECT -4.800 2836.020 2.400 2836.470 ;
        RECT 15.705 2836.455 16.035 2836.470 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2219.185 3195.405 2219.355 3199.655 ;
      LAYER mcon ;
        RECT 2219.185 3199.485 2219.355 3199.655 ;
      LAYER met1 ;
        RECT 2219.110 3199.640 2219.430 3199.700 ;
        RECT 2218.915 3199.500 2219.430 3199.640 ;
        RECT 2219.110 3199.440 2219.430 3199.500 ;
        RECT 32.730 3195.560 33.050 3195.620 ;
        RECT 2219.125 3195.560 2219.415 3195.605 ;
        RECT 32.730 3195.420 2219.415 3195.560 ;
        RECT 32.730 3195.360 33.050 3195.420 ;
        RECT 2219.125 3195.375 2219.415 3195.420 ;
        RECT 16.170 2551.940 16.490 2552.000 ;
        RECT 32.730 2551.940 33.050 2552.000 ;
        RECT 16.170 2551.800 33.050 2551.940 ;
        RECT 16.170 2551.740 16.490 2551.800 ;
        RECT 32.730 2551.740 33.050 2551.800 ;
      LAYER via ;
        RECT 2219.140 3199.440 2219.400 3199.700 ;
        RECT 32.760 3195.360 33.020 3195.620 ;
        RECT 16.200 2551.740 16.460 2552.000 ;
        RECT 32.760 2551.740 33.020 2552.000 ;
      LAYER met2 ;
        RECT 2220.900 3199.810 2221.180 3200.000 ;
        RECT 2219.200 3199.730 2221.180 3199.810 ;
        RECT 2219.140 3199.670 2221.180 3199.730 ;
        RECT 2219.140 3199.410 2219.400 3199.670 ;
        RECT 2220.900 3196.000 2221.180 3199.670 ;
        RECT 32.760 3195.330 33.020 3195.650 ;
        RECT 32.820 2552.030 32.960 3195.330 ;
        RECT 16.200 2551.710 16.460 2552.030 ;
        RECT 32.760 2551.710 33.020 2552.030 ;
        RECT 16.260 2549.845 16.400 2551.710 ;
        RECT 16.190 2549.475 16.470 2549.845 ;
      LAYER via2 ;
        RECT 16.190 2549.520 16.470 2549.800 ;
      LAYER met3 ;
        RECT -4.800 2549.810 2.400 2550.260 ;
        RECT 16.165 2549.810 16.495 2549.825 ;
        RECT -4.800 2549.510 16.495 2549.810 ;
        RECT -4.800 2549.060 2.400 2549.510 ;
        RECT 16.165 2549.495 16.495 2549.510 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2258.745 3195.065 2258.915 3199.655 ;
      LAYER mcon ;
        RECT 2258.745 3199.485 2258.915 3199.655 ;
      LAYER met1 ;
        RECT 2258.670 3199.640 2258.990 3199.700 ;
        RECT 2258.475 3199.500 2258.990 3199.640 ;
        RECT 2258.670 3199.440 2258.990 3199.500 ;
        RECT 32.270 3195.220 32.590 3195.280 ;
        RECT 2258.685 3195.220 2258.975 3195.265 ;
        RECT 32.270 3195.080 2258.975 3195.220 ;
        RECT 32.270 3195.020 32.590 3195.080 ;
        RECT 2258.685 3195.035 2258.975 3195.080 ;
        RECT 15.710 2262.260 16.030 2262.320 ;
        RECT 32.270 2262.260 32.590 2262.320 ;
        RECT 15.710 2262.120 32.590 2262.260 ;
        RECT 15.710 2262.060 16.030 2262.120 ;
        RECT 32.270 2262.060 32.590 2262.120 ;
      LAYER via ;
        RECT 2258.700 3199.440 2258.960 3199.700 ;
        RECT 32.300 3195.020 32.560 3195.280 ;
        RECT 15.740 2262.060 16.000 2262.320 ;
        RECT 32.300 2262.060 32.560 2262.320 ;
      LAYER met2 ;
        RECT 2260.000 3199.810 2260.280 3200.000 ;
        RECT 2258.760 3199.730 2260.280 3199.810 ;
        RECT 2258.700 3199.670 2260.280 3199.730 ;
        RECT 2258.700 3199.410 2258.960 3199.670 ;
        RECT 2260.000 3196.000 2260.280 3199.670 ;
        RECT 32.300 3194.990 32.560 3195.310 ;
        RECT 32.360 2262.350 32.500 3194.990 ;
        RECT 15.740 2262.205 16.000 2262.350 ;
        RECT 15.730 2261.835 16.010 2262.205 ;
        RECT 32.300 2262.030 32.560 2262.350 ;
      LAYER via2 ;
        RECT 15.730 2261.880 16.010 2262.160 ;
      LAYER met3 ;
        RECT -4.800 2262.170 2.400 2262.620 ;
        RECT 15.705 2262.170 16.035 2262.185 ;
        RECT -4.800 2261.870 16.035 2262.170 ;
        RECT -4.800 2261.420 2.400 2261.870 ;
        RECT 15.705 2261.855 16.035 2261.870 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 16.630 3211.200 16.950 3211.260 ;
        RECT 2299.610 3211.200 2299.930 3211.260 ;
        RECT 16.630 3211.060 2299.930 3211.200 ;
        RECT 16.630 3211.000 16.950 3211.060 ;
        RECT 2299.610 3211.000 2299.930 3211.060 ;
      LAYER via ;
        RECT 16.660 3211.000 16.920 3211.260 ;
        RECT 2299.640 3211.000 2299.900 3211.260 ;
      LAYER met2 ;
        RECT 16.660 3210.970 16.920 3211.290 ;
        RECT 2299.640 3210.970 2299.900 3211.290 ;
        RECT 16.720 1975.245 16.860 3210.970 ;
        RECT 2299.700 3200.000 2299.840 3210.970 ;
        RECT 2299.560 3196.000 2299.840 3200.000 ;
        RECT 16.650 1974.875 16.930 1975.245 ;
      LAYER via2 ;
        RECT 16.650 1974.920 16.930 1975.200 ;
      LAYER met3 ;
        RECT -4.800 1975.210 2.400 1975.660 ;
        RECT 16.625 1975.210 16.955 1975.225 ;
        RECT -4.800 1974.910 16.955 1975.210 ;
        RECT -4.800 1974.460 2.400 1974.910 ;
        RECT 16.625 1974.895 16.955 1974.910 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1683.670 553.760 1683.990 553.820 ;
        RECT 1731.050 553.760 1731.370 553.820 ;
        RECT 1683.670 553.620 1731.370 553.760 ;
        RECT 1683.670 553.560 1683.990 553.620 ;
        RECT 1731.050 553.560 1731.370 553.620 ;
        RECT 2125.270 552.740 2125.590 552.800 ;
        RECT 2172.650 552.740 2172.970 552.800 ;
        RECT 2125.270 552.600 2172.970 552.740 ;
        RECT 2125.270 552.540 2125.590 552.600 ;
        RECT 2172.650 552.540 2172.970 552.600 ;
        RECT 2608.270 552.740 2608.590 552.800 ;
        RECT 2632.190 552.740 2632.510 552.800 ;
        RECT 2608.270 552.600 2632.510 552.740 ;
        RECT 2608.270 552.540 2608.590 552.600 ;
        RECT 2632.190 552.540 2632.510 552.600 ;
      LAYER via ;
        RECT 1683.700 553.560 1683.960 553.820 ;
        RECT 1731.080 553.560 1731.340 553.820 ;
        RECT 2125.300 552.540 2125.560 552.800 ;
        RECT 2172.680 552.540 2172.940 552.800 ;
        RECT 2608.300 552.540 2608.560 552.800 ;
        RECT 2632.220 552.540 2632.480 552.800 ;
      LAYER met2 ;
        RECT 1233.740 3196.410 1234.020 3200.000 ;
        RECT 1234.730 3196.410 1235.010 3196.525 ;
        RECT 1233.740 3196.270 1235.010 3196.410 ;
        RECT 1233.740 3196.000 1234.020 3196.270 ;
        RECT 1234.730 3196.155 1235.010 3196.270 ;
        RECT 1393.890 554.355 1394.170 554.725 ;
        RECT 2704.430 554.355 2704.710 554.725 ;
        RECT 1393.960 552.685 1394.100 554.355 ;
        RECT 1490.030 553.675 1490.310 554.045 ;
        RECT 1683.690 553.675 1683.970 554.045 ;
        RECT 1490.100 552.685 1490.240 553.675 ;
        RECT 1683.700 553.530 1683.960 553.675 ;
        RECT 1731.080 553.530 1731.340 553.850 ;
        RECT 2172.670 553.675 2172.950 554.045 ;
        RECT 1731.140 552.685 1731.280 553.530 ;
        RECT 2090.330 552.995 2090.610 553.365 ;
        RECT 1393.890 552.315 1394.170 552.685 ;
        RECT 1490.030 552.315 1490.310 552.685 ;
        RECT 1731.070 552.315 1731.350 552.685 ;
        RECT 2090.400 551.325 2090.540 552.995 ;
        RECT 2172.740 552.830 2172.880 553.675 ;
        RECT 2572.870 552.995 2573.150 553.365 ;
        RECT 2632.210 552.995 2632.490 553.365 ;
        RECT 2125.300 552.685 2125.560 552.830 ;
        RECT 2125.290 552.315 2125.570 552.685 ;
        RECT 2172.680 552.510 2172.940 552.830 ;
        RECT 2572.940 551.325 2573.080 552.995 ;
        RECT 2632.280 552.830 2632.420 552.995 ;
        RECT 2608.300 552.685 2608.560 552.830 ;
        RECT 2608.290 552.315 2608.570 552.685 ;
        RECT 2632.220 552.510 2632.480 552.830 ;
        RECT 2704.500 552.685 2704.640 554.355 ;
        RECT 2801.030 553.675 2801.310 554.045 ;
        RECT 2704.430 552.315 2704.710 552.685 ;
        RECT 2801.100 552.005 2801.240 553.675 ;
        RECT 2863.130 552.995 2863.410 553.365 ;
        RECT 2863.200 552.570 2863.340 552.995 ;
        RECT 2863.590 552.570 2863.870 552.685 ;
        RECT 2863.200 552.430 2863.870 552.570 ;
        RECT 2863.590 552.315 2863.870 552.430 ;
        RECT 2801.030 551.635 2801.310 552.005 ;
        RECT 2090.330 550.955 2090.610 551.325 ;
        RECT 2572.870 550.955 2573.150 551.325 ;
      LAYER via2 ;
        RECT 1234.730 3196.200 1235.010 3196.480 ;
        RECT 1393.890 554.400 1394.170 554.680 ;
        RECT 2704.430 554.400 2704.710 554.680 ;
        RECT 1490.030 553.720 1490.310 554.000 ;
        RECT 1683.690 553.720 1683.970 554.000 ;
        RECT 2172.670 553.720 2172.950 554.000 ;
        RECT 2090.330 553.040 2090.610 553.320 ;
        RECT 1393.890 552.360 1394.170 552.640 ;
        RECT 1490.030 552.360 1490.310 552.640 ;
        RECT 1731.070 552.360 1731.350 552.640 ;
        RECT 2572.870 553.040 2573.150 553.320 ;
        RECT 2632.210 553.040 2632.490 553.320 ;
        RECT 2125.290 552.360 2125.570 552.640 ;
        RECT 2608.290 552.360 2608.570 552.640 ;
        RECT 2801.030 553.720 2801.310 554.000 ;
        RECT 2704.430 552.360 2704.710 552.640 ;
        RECT 2863.130 553.040 2863.410 553.320 ;
        RECT 2863.590 552.360 2863.870 552.640 ;
        RECT 2801.030 551.680 2801.310 551.960 ;
        RECT 2090.330 551.000 2090.610 551.280 ;
        RECT 2572.870 551.000 2573.150 551.280 ;
      LAYER met3 ;
        RECT 1234.705 3196.490 1235.035 3196.505 ;
        RECT 1237.670 3196.490 1238.050 3196.500 ;
        RECT 1234.705 3196.190 1238.050 3196.490 ;
        RECT 1234.705 3196.175 1235.035 3196.190 ;
        RECT 1237.670 3196.180 1238.050 3196.190 ;
        RECT 2917.600 557.410 2924.800 557.860 ;
        RECT 2916.710 557.110 2924.800 557.410 ;
        RECT 1635.110 555.370 1635.490 555.380 ;
        RECT 1635.110 555.070 1683.290 555.370 ;
        RECT 1635.110 555.060 1635.490 555.070 ;
        RECT 1393.865 554.690 1394.195 554.705 ;
        RECT 1345.350 554.390 1394.195 554.690 ;
        RECT 1237.670 553.330 1238.050 553.340 ;
        RECT 1345.350 553.330 1345.650 554.390 ;
        RECT 1393.865 554.375 1394.195 554.390 ;
        RECT 1490.005 554.010 1490.335 554.025 ;
        RECT 1635.110 554.010 1635.490 554.020 ;
        RECT 1490.005 553.710 1491.010 554.010 ;
        RECT 1490.005 553.695 1490.335 553.710 ;
        RECT 1490.710 553.340 1491.010 553.710 ;
        RECT 1558.790 553.710 1635.490 554.010 ;
        RECT 1682.990 554.010 1683.290 555.070 ;
        RECT 2316.830 554.690 2317.210 554.700 ;
        RECT 2510.030 554.690 2510.410 554.700 ;
        RECT 2282.830 554.390 2317.210 554.690 ;
        RECT 1683.665 554.010 1683.995 554.025 ;
        RECT 1786.910 554.010 1787.290 554.020 ;
        RECT 2172.645 554.010 2172.975 554.025 ;
        RECT 1682.990 553.710 1683.995 554.010 ;
        RECT 1237.670 553.030 1345.650 553.330 ;
        RECT 1237.670 553.020 1238.050 553.030 ;
        RECT 1490.670 553.020 1491.050 553.340 ;
        RECT 1393.865 552.650 1394.195 552.665 ;
        RECT 1490.005 552.650 1490.335 552.665 ;
        RECT 1393.865 552.350 1490.335 552.650 ;
        RECT 1393.865 552.335 1394.195 552.350 ;
        RECT 1490.005 552.335 1490.335 552.350 ;
        RECT 1490.670 552.650 1491.050 552.660 ;
        RECT 1558.790 552.650 1559.090 553.710 ;
        RECT 1635.110 553.700 1635.490 553.710 ;
        RECT 1683.665 553.695 1683.995 553.710 ;
        RECT 1755.670 553.710 1787.290 554.010 ;
        RECT 1490.670 552.350 1559.090 552.650 ;
        RECT 1731.045 552.650 1731.375 552.665 ;
        RECT 1755.670 552.650 1755.970 553.710 ;
        RECT 1786.910 553.700 1787.290 553.710 ;
        RECT 1970.030 553.710 1994.250 554.010 ;
        RECT 1970.030 553.330 1970.330 553.710 ;
        RECT 1836.630 553.030 1970.330 553.330 ;
        RECT 1731.045 552.350 1755.970 552.650 ;
        RECT 1787.830 552.650 1788.210 552.660 ;
        RECT 1836.630 552.650 1836.930 553.030 ;
        RECT 1787.830 552.350 1836.930 552.650 ;
        RECT 1993.950 552.650 1994.250 553.710 ;
        RECT 2172.645 553.710 2187.450 554.010 ;
        RECT 2172.645 553.695 2172.975 553.710 ;
        RECT 2090.305 553.330 2090.635 553.345 ;
        RECT 2042.710 553.030 2090.635 553.330 ;
        RECT 2042.710 552.650 2043.010 553.030 ;
        RECT 2090.305 553.015 2090.635 553.030 ;
        RECT 2125.265 552.650 2125.595 552.665 ;
        RECT 1993.950 552.350 2043.010 552.650 ;
        RECT 2124.590 552.350 2125.595 552.650 ;
        RECT 2187.150 552.650 2187.450 553.710 ;
        RECT 2282.830 553.330 2283.130 554.390 ;
        RECT 2316.830 554.380 2317.210 554.390 ;
        RECT 2476.030 554.390 2510.410 554.690 ;
        RECT 2476.030 553.330 2476.330 554.390 ;
        RECT 2510.030 554.380 2510.410 554.390 ;
        RECT 2656.310 554.690 2656.690 554.700 ;
        RECT 2704.405 554.690 2704.735 554.705 ;
        RECT 2656.310 554.390 2704.735 554.690 ;
        RECT 2656.310 554.380 2656.690 554.390 ;
        RECT 2704.405 554.375 2704.735 554.390 ;
        RECT 2801.005 554.010 2801.335 554.025 ;
        RECT 2801.005 553.710 2815.810 554.010 ;
        RECT 2801.005 553.695 2801.335 553.710 ;
        RECT 2572.845 553.330 2573.175 553.345 ;
        RECT 2235.910 553.030 2283.130 553.330 ;
        RECT 2332.510 553.030 2379.730 553.330 ;
        RECT 2235.910 552.650 2236.210 553.030 ;
        RECT 2187.150 552.350 2236.210 552.650 ;
        RECT 2317.750 552.650 2318.130 552.660 ;
        RECT 2332.510 552.650 2332.810 553.030 ;
        RECT 2317.750 552.350 2332.810 552.650 ;
        RECT 2379.430 552.650 2379.730 553.030 ;
        RECT 2429.110 553.030 2476.330 553.330 ;
        RECT 2525.710 553.030 2573.175 553.330 ;
        RECT 2429.110 552.650 2429.410 553.030 ;
        RECT 2379.430 552.350 2429.410 552.650 ;
        RECT 2510.950 552.650 2511.330 552.660 ;
        RECT 2525.710 552.650 2526.010 553.030 ;
        RECT 2572.845 553.015 2573.175 553.030 ;
        RECT 2632.185 553.330 2632.515 553.345 ;
        RECT 2656.310 553.330 2656.690 553.340 ;
        RECT 2752.910 553.330 2753.290 553.340 ;
        RECT 2632.185 553.030 2656.690 553.330 ;
        RECT 2632.185 553.015 2632.515 553.030 ;
        RECT 2656.310 553.020 2656.690 553.030 ;
        RECT 2718.910 553.030 2753.290 553.330 ;
        RECT 2608.265 552.650 2608.595 552.665 ;
        RECT 2510.950 552.350 2526.010 552.650 ;
        RECT 2607.590 552.350 2608.595 552.650 ;
        RECT 1490.670 552.340 1491.050 552.350 ;
        RECT 1731.045 552.335 1731.375 552.350 ;
        RECT 1787.830 552.340 1788.210 552.350 ;
        RECT 2090.305 551.290 2090.635 551.305 ;
        RECT 2124.590 551.290 2124.890 552.350 ;
        RECT 2125.265 552.335 2125.595 552.350 ;
        RECT 2317.750 552.340 2318.130 552.350 ;
        RECT 2510.950 552.340 2511.330 552.350 ;
        RECT 2090.305 550.990 2124.890 551.290 ;
        RECT 2572.845 551.290 2573.175 551.305 ;
        RECT 2607.590 551.290 2607.890 552.350 ;
        RECT 2608.265 552.335 2608.595 552.350 ;
        RECT 2704.405 552.650 2704.735 552.665 ;
        RECT 2718.910 552.650 2719.210 553.030 ;
        RECT 2752.910 553.020 2753.290 553.030 ;
        RECT 2704.405 552.350 2719.210 552.650 ;
        RECT 2815.510 552.650 2815.810 553.710 ;
        RECT 2863.105 553.330 2863.435 553.345 ;
        RECT 2916.710 553.330 2917.010 557.110 ;
        RECT 2917.600 556.660 2924.800 557.110 ;
        RECT 2849.550 553.030 2863.435 553.330 ;
        RECT 2849.550 552.650 2849.850 553.030 ;
        RECT 2863.105 553.015 2863.435 553.030 ;
        RECT 2884.510 553.030 2917.010 553.330 ;
        RECT 2815.510 552.350 2849.850 552.650 ;
        RECT 2863.565 552.650 2863.895 552.665 ;
        RECT 2884.510 552.650 2884.810 553.030 ;
        RECT 2863.565 552.350 2884.810 552.650 ;
        RECT 2704.405 552.335 2704.735 552.350 ;
        RECT 2863.565 552.335 2863.895 552.350 ;
        RECT 2752.910 551.970 2753.290 551.980 ;
        RECT 2801.005 551.970 2801.335 551.985 ;
        RECT 2752.910 551.670 2801.335 551.970 ;
        RECT 2752.910 551.660 2753.290 551.670 ;
        RECT 2801.005 551.655 2801.335 551.670 ;
        RECT 2572.845 550.990 2607.890 551.290 ;
        RECT 2090.305 550.975 2090.635 550.990 ;
        RECT 2572.845 550.975 2573.175 550.990 ;
      LAYER via3 ;
        RECT 1237.700 3196.180 1238.020 3196.500 ;
        RECT 1635.140 555.060 1635.460 555.380 ;
        RECT 1237.700 553.020 1238.020 553.340 ;
        RECT 1490.700 553.020 1491.020 553.340 ;
        RECT 1490.700 552.340 1491.020 552.660 ;
        RECT 1635.140 553.700 1635.460 554.020 ;
        RECT 1786.940 553.700 1787.260 554.020 ;
        RECT 1787.860 552.340 1788.180 552.660 ;
        RECT 2316.860 554.380 2317.180 554.700 ;
        RECT 2510.060 554.380 2510.380 554.700 ;
        RECT 2656.340 554.380 2656.660 554.700 ;
        RECT 2317.780 552.340 2318.100 552.660 ;
        RECT 2510.980 552.340 2511.300 552.660 ;
        RECT 2656.340 553.020 2656.660 553.340 ;
        RECT 2752.940 553.020 2753.260 553.340 ;
        RECT 2752.940 551.660 2753.260 551.980 ;
      LAYER met4 ;
        RECT 1237.695 3196.175 1238.025 3196.505 ;
        RECT 1237.710 553.345 1238.010 3196.175 ;
        RECT 1635.135 555.055 1635.465 555.385 ;
        RECT 1635.150 554.025 1635.450 555.055 ;
        RECT 2316.855 554.375 2317.185 554.705 ;
        RECT 2510.055 554.375 2510.385 554.705 ;
        RECT 2656.335 554.375 2656.665 554.705 ;
        RECT 1635.135 553.695 1635.465 554.025 ;
        RECT 1786.935 553.695 1787.265 554.025 ;
        RECT 1237.695 553.015 1238.025 553.345 ;
        RECT 1490.695 553.015 1491.025 553.345 ;
        RECT 1490.710 552.665 1491.010 553.015 ;
        RECT 1490.695 552.335 1491.025 552.665 ;
        RECT 1786.950 552.650 1787.250 553.695 ;
        RECT 1787.855 552.650 1788.185 552.665 ;
        RECT 1786.950 552.350 1788.185 552.650 ;
        RECT 2316.870 552.650 2317.170 554.375 ;
        RECT 2317.775 552.650 2318.105 552.665 ;
        RECT 2316.870 552.350 2318.105 552.650 ;
        RECT 2510.070 552.650 2510.370 554.375 ;
        RECT 2656.350 553.345 2656.650 554.375 ;
        RECT 2656.335 553.015 2656.665 553.345 ;
        RECT 2752.935 553.015 2753.265 553.345 ;
        RECT 2510.975 552.650 2511.305 552.665 ;
        RECT 2510.070 552.350 2511.305 552.650 ;
        RECT 1787.855 552.335 1788.185 552.350 ;
        RECT 2317.775 552.335 2318.105 552.350 ;
        RECT 2510.975 552.335 2511.305 552.350 ;
        RECT 2752.950 551.985 2753.250 553.015 ;
        RECT 2752.935 551.655 2753.265 551.985 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 39.170 3203.380 39.490 3203.440 ;
        RECT 2339.170 3203.380 2339.490 3203.440 ;
        RECT 39.170 3203.240 2339.490 3203.380 ;
        RECT 39.170 3203.180 39.490 3203.240 ;
        RECT 2339.170 3203.180 2339.490 3203.240 ;
        RECT 16.630 1687.660 16.950 1687.720 ;
        RECT 39.170 1687.660 39.490 1687.720 ;
        RECT 16.630 1687.520 39.490 1687.660 ;
        RECT 16.630 1687.460 16.950 1687.520 ;
        RECT 39.170 1687.460 39.490 1687.520 ;
      LAYER via ;
        RECT 39.200 3203.180 39.460 3203.440 ;
        RECT 2339.200 3203.180 2339.460 3203.440 ;
        RECT 16.660 1687.460 16.920 1687.720 ;
        RECT 39.200 1687.460 39.460 1687.720 ;
      LAYER met2 ;
        RECT 39.200 3203.150 39.460 3203.470 ;
        RECT 2339.200 3203.150 2339.460 3203.470 ;
        RECT 39.260 1687.750 39.400 3203.150 ;
        RECT 2339.260 3200.000 2339.400 3203.150 ;
        RECT 2339.120 3196.000 2339.400 3200.000 ;
        RECT 16.660 1687.605 16.920 1687.750 ;
        RECT 16.650 1687.235 16.930 1687.605 ;
        RECT 39.200 1687.430 39.460 1687.750 ;
      LAYER via2 ;
        RECT 16.650 1687.280 16.930 1687.560 ;
      LAYER met3 ;
        RECT -4.800 1687.570 2.400 1688.020 ;
        RECT 16.625 1687.570 16.955 1687.585 ;
        RECT -4.800 1687.270 16.955 1687.570 ;
        RECT -4.800 1686.820 2.400 1687.270 ;
        RECT 16.625 1687.255 16.955 1687.270 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 38.710 3203.040 39.030 3203.100 ;
        RECT 2378.730 3203.040 2379.050 3203.100 ;
        RECT 38.710 3202.900 2379.050 3203.040 ;
        RECT 38.710 3202.840 39.030 3202.900 ;
        RECT 2378.730 3202.840 2379.050 3202.900 ;
        RECT 16.630 1474.820 16.950 1474.880 ;
        RECT 38.710 1474.820 39.030 1474.880 ;
        RECT 16.630 1474.680 39.030 1474.820 ;
        RECT 16.630 1474.620 16.950 1474.680 ;
        RECT 38.710 1474.620 39.030 1474.680 ;
      LAYER via ;
        RECT 38.740 3202.840 39.000 3203.100 ;
        RECT 2378.760 3202.840 2379.020 3203.100 ;
        RECT 16.660 1474.620 16.920 1474.880 ;
        RECT 38.740 1474.620 39.000 1474.880 ;
      LAYER met2 ;
        RECT 38.740 3202.810 39.000 3203.130 ;
        RECT 2378.760 3202.810 2379.020 3203.130 ;
        RECT 38.800 1474.910 38.940 3202.810 ;
        RECT 2378.820 3200.000 2378.960 3202.810 ;
        RECT 2378.680 3196.000 2378.960 3200.000 ;
        RECT 16.660 1474.590 16.920 1474.910 ;
        RECT 38.740 1474.590 39.000 1474.910 ;
        RECT 16.720 1472.045 16.860 1474.590 ;
        RECT 16.650 1471.675 16.930 1472.045 ;
      LAYER via2 ;
        RECT 16.650 1471.720 16.930 1472.000 ;
      LAYER met3 ;
        RECT -4.800 1472.010 2.400 1472.460 ;
        RECT 16.625 1472.010 16.955 1472.025 ;
        RECT -4.800 1471.710 16.955 1472.010 ;
        RECT -4.800 1471.260 2.400 1471.710 ;
        RECT 16.625 1471.695 16.955 1471.710 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2418.310 3211.795 2418.590 3212.165 ;
        RECT 2418.380 3200.000 2418.520 3211.795 ;
        RECT 2418.240 3196.000 2418.520 3200.000 ;
        RECT 15.730 1262.235 16.010 1262.605 ;
        RECT 15.800 1256.485 15.940 1262.235 ;
        RECT 15.730 1256.115 16.010 1256.485 ;
      LAYER via2 ;
        RECT 2418.310 3211.840 2418.590 3212.120 ;
        RECT 15.730 1262.280 16.010 1262.560 ;
        RECT 15.730 1256.160 16.010 1256.440 ;
      LAYER met3 ;
        RECT 1308.510 3212.130 1308.890 3212.140 ;
        RECT 2418.285 3212.130 2418.615 3212.145 ;
        RECT 1308.510 3211.830 2418.615 3212.130 ;
        RECT 1308.510 3211.820 1308.890 3211.830 ;
        RECT 2418.285 3211.815 2418.615 3211.830 ;
        RECT 15.705 1262.570 16.035 1262.585 ;
        RECT 1308.510 1262.570 1308.890 1262.580 ;
        RECT 15.705 1262.270 1169.930 1262.570 ;
        RECT 15.705 1262.255 16.035 1262.270 ;
        RECT 1169.630 1261.890 1169.930 1262.270 ;
        RECT 1172.390 1262.270 1308.890 1262.570 ;
        RECT 1172.390 1261.890 1172.690 1262.270 ;
        RECT 1308.510 1262.260 1308.890 1262.270 ;
        RECT 1169.630 1261.590 1172.690 1261.890 ;
        RECT -4.800 1256.450 2.400 1256.900 ;
        RECT 15.705 1256.450 16.035 1256.465 ;
        RECT -4.800 1256.150 16.035 1256.450 ;
        RECT -4.800 1255.700 2.400 1256.150 ;
        RECT 15.705 1256.135 16.035 1256.150 ;
      LAYER via3 ;
        RECT 1308.540 3211.820 1308.860 3212.140 ;
        RECT 1308.540 1262.260 1308.860 1262.580 ;
      LAYER met4 ;
        RECT 1308.535 3211.815 1308.865 3212.145 ;
        RECT 1308.550 1262.585 1308.850 3211.815 ;
        RECT 1308.535 1262.255 1308.865 1262.585 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2457.410 3211.115 2457.690 3211.485 ;
        RECT 2457.480 3200.000 2457.620 3211.115 ;
        RECT 2457.340 3196.000 2457.620 3200.000 ;
      LAYER via2 ;
        RECT 2457.410 3211.160 2457.690 3211.440 ;
      LAYER met3 ;
        RECT 1307.590 3211.450 1307.970 3211.460 ;
        RECT 2457.385 3211.450 2457.715 3211.465 ;
        RECT 1307.590 3211.150 2457.715 3211.450 ;
        RECT 1307.590 3211.140 1307.970 3211.150 ;
        RECT 2457.385 3211.135 2457.715 3211.150 ;
        RECT 1307.590 1041.570 1307.970 1041.580 ;
        RECT -4.800 1040.890 2.400 1041.340 ;
        RECT 3.070 1041.270 1307.970 1041.570 ;
        RECT 3.070 1040.890 3.370 1041.270 ;
        RECT 1307.590 1041.260 1307.970 1041.270 ;
        RECT -4.800 1040.590 3.370 1040.890 ;
        RECT -4.800 1040.140 2.400 1040.590 ;
      LAYER via3 ;
        RECT 1307.620 3211.140 1307.940 3211.460 ;
        RECT 1307.620 1041.260 1307.940 1041.580 ;
      LAYER met4 ;
        RECT 1307.615 3211.135 1307.945 3211.465 ;
        RECT 1307.630 1041.585 1307.930 3211.135 ;
        RECT 1307.615 1041.255 1307.945 1041.585 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 23.990 3202.700 24.310 3202.760 ;
        RECT 2496.950 3202.700 2497.270 3202.760 ;
        RECT 23.990 3202.560 2497.270 3202.700 ;
        RECT 23.990 3202.500 24.310 3202.560 ;
        RECT 2496.950 3202.500 2497.270 3202.560 ;
        RECT 13.870 825.760 14.190 825.820 ;
        RECT 23.990 825.760 24.310 825.820 ;
        RECT 13.870 825.620 24.310 825.760 ;
        RECT 13.870 825.560 14.190 825.620 ;
        RECT 23.990 825.560 24.310 825.620 ;
      LAYER via ;
        RECT 24.020 3202.500 24.280 3202.760 ;
        RECT 2496.980 3202.500 2497.240 3202.760 ;
        RECT 13.900 825.560 14.160 825.820 ;
        RECT 24.020 825.560 24.280 825.820 ;
      LAYER met2 ;
        RECT 24.020 3202.470 24.280 3202.790 ;
        RECT 2496.980 3202.470 2497.240 3202.790 ;
        RECT 24.080 825.850 24.220 3202.470 ;
        RECT 2497.040 3200.000 2497.180 3202.470 ;
        RECT 2496.900 3196.000 2497.180 3200.000 ;
        RECT 13.900 825.530 14.160 825.850 ;
        RECT 24.020 825.530 24.280 825.850 ;
        RECT 13.960 825.365 14.100 825.530 ;
        RECT 13.890 824.995 14.170 825.365 ;
      LAYER via2 ;
        RECT 13.890 825.040 14.170 825.320 ;
      LAYER met3 ;
        RECT -4.800 825.330 2.400 825.780 ;
        RECT 13.865 825.330 14.195 825.345 ;
        RECT -4.800 825.030 14.195 825.330 ;
        RECT -4.800 824.580 2.400 825.030 ;
        RECT 13.865 825.015 14.195 825.030 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 30.890 3202.360 31.210 3202.420 ;
        RECT 2536.510 3202.360 2536.830 3202.420 ;
        RECT 30.890 3202.220 2536.830 3202.360 ;
        RECT 30.890 3202.160 31.210 3202.220 ;
        RECT 2536.510 3202.160 2536.830 3202.220 ;
        RECT 14.790 611.220 15.110 611.280 ;
        RECT 30.890 611.220 31.210 611.280 ;
        RECT 14.790 611.080 31.210 611.220 ;
        RECT 14.790 611.020 15.110 611.080 ;
        RECT 30.890 611.020 31.210 611.080 ;
      LAYER via ;
        RECT 30.920 3202.160 31.180 3202.420 ;
        RECT 2536.540 3202.160 2536.800 3202.420 ;
        RECT 14.820 611.020 15.080 611.280 ;
        RECT 30.920 611.020 31.180 611.280 ;
      LAYER met2 ;
        RECT 30.920 3202.130 31.180 3202.450 ;
        RECT 2536.540 3202.130 2536.800 3202.450 ;
        RECT 30.980 611.310 31.120 3202.130 ;
        RECT 2536.600 3200.000 2536.740 3202.130 ;
        RECT 2536.460 3196.000 2536.740 3200.000 ;
        RECT 14.820 610.990 15.080 611.310 ;
        RECT 30.920 610.990 31.180 611.310 ;
        RECT 14.880 610.485 15.020 610.990 ;
        RECT 14.810 610.115 15.090 610.485 ;
      LAYER via2 ;
        RECT 14.810 610.160 15.090 610.440 ;
      LAYER met3 ;
        RECT -4.800 610.450 2.400 610.900 ;
        RECT 14.785 610.450 15.115 610.465 ;
        RECT -4.800 610.150 15.115 610.450 ;
        RECT -4.800 609.700 2.400 610.150 ;
        RECT 14.785 610.135 15.115 610.150 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 38.250 3202.020 38.570 3202.080 ;
        RECT 2576.070 3202.020 2576.390 3202.080 ;
        RECT 38.250 3201.880 2576.390 3202.020 ;
        RECT 38.250 3201.820 38.570 3201.880 ;
        RECT 2576.070 3201.820 2576.390 3201.880 ;
        RECT 16.630 396.000 16.950 396.060 ;
        RECT 38.250 396.000 38.570 396.060 ;
        RECT 16.630 395.860 38.570 396.000 ;
        RECT 16.630 395.800 16.950 395.860 ;
        RECT 38.250 395.800 38.570 395.860 ;
      LAYER via ;
        RECT 38.280 3201.820 38.540 3202.080 ;
        RECT 2576.100 3201.820 2576.360 3202.080 ;
        RECT 16.660 395.800 16.920 396.060 ;
        RECT 38.280 395.800 38.540 396.060 ;
      LAYER met2 ;
        RECT 38.280 3201.790 38.540 3202.110 ;
        RECT 2576.100 3201.790 2576.360 3202.110 ;
        RECT 38.340 396.090 38.480 3201.790 ;
        RECT 2576.160 3200.000 2576.300 3201.790 ;
        RECT 2576.020 3196.000 2576.300 3200.000 ;
        RECT 16.660 395.770 16.920 396.090 ;
        RECT 38.280 395.770 38.540 396.090 ;
        RECT 16.720 394.925 16.860 395.770 ;
        RECT 16.650 394.555 16.930 394.925 ;
      LAYER via2 ;
        RECT 16.650 394.600 16.930 394.880 ;
      LAYER met3 ;
        RECT -4.800 394.890 2.400 395.340 ;
        RECT 16.625 394.890 16.955 394.905 ;
        RECT -4.800 394.590 16.955 394.890 ;
        RECT -4.800 394.140 2.400 394.590 ;
        RECT 16.625 394.575 16.955 394.590 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 37.790 3201.680 38.110 3201.740 ;
        RECT 2615.630 3201.680 2615.950 3201.740 ;
        RECT 37.790 3201.540 2615.950 3201.680 ;
        RECT 37.790 3201.480 38.110 3201.540 ;
        RECT 2615.630 3201.480 2615.950 3201.540 ;
        RECT 17.550 179.420 17.870 179.480 ;
        RECT 37.790 179.420 38.110 179.480 ;
        RECT 17.550 179.280 38.110 179.420 ;
        RECT 17.550 179.220 17.870 179.280 ;
        RECT 37.790 179.220 38.110 179.280 ;
      LAYER via ;
        RECT 37.820 3201.480 38.080 3201.740 ;
        RECT 2615.660 3201.480 2615.920 3201.740 ;
        RECT 17.580 179.220 17.840 179.480 ;
        RECT 37.820 179.220 38.080 179.480 ;
      LAYER met2 ;
        RECT 37.820 3201.450 38.080 3201.770 ;
        RECT 2615.660 3201.450 2615.920 3201.770 ;
        RECT 37.880 179.510 38.020 3201.450 ;
        RECT 2615.720 3200.000 2615.860 3201.450 ;
        RECT 2615.580 3196.000 2615.860 3200.000 ;
        RECT 17.580 179.365 17.840 179.510 ;
        RECT 17.570 178.995 17.850 179.365 ;
        RECT 37.820 179.190 38.080 179.510 ;
      LAYER via2 ;
        RECT 17.570 179.040 17.850 179.320 ;
      LAYER met3 ;
        RECT -4.800 179.330 2.400 179.780 ;
        RECT 17.545 179.330 17.875 179.345 ;
        RECT -4.800 179.030 17.875 179.330 ;
        RECT -4.800 178.580 2.400 179.030 ;
        RECT 17.545 179.015 17.875 179.030 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2028.670 788.700 2028.990 788.760 ;
        RECT 2076.510 788.700 2076.830 788.760 ;
        RECT 2028.670 788.560 2076.830 788.700 ;
        RECT 2028.670 788.500 2028.990 788.560 ;
        RECT 2076.510 788.500 2076.830 788.560 ;
        RECT 2608.270 787.340 2608.590 787.400 ;
        RECT 2632.190 787.340 2632.510 787.400 ;
        RECT 2608.270 787.200 2632.510 787.340 ;
        RECT 2608.270 787.140 2608.590 787.200 ;
        RECT 2632.190 787.140 2632.510 787.200 ;
      LAYER via ;
        RECT 2028.700 788.500 2028.960 788.760 ;
        RECT 2076.540 788.500 2076.800 788.760 ;
        RECT 2608.300 787.140 2608.560 787.400 ;
        RECT 2632.220 787.140 2632.480 787.400 ;
      LAYER met2 ;
        RECT 1273.300 3196.410 1273.580 3200.000 ;
        RECT 1274.750 3196.410 1275.030 3196.525 ;
        RECT 1273.300 3196.270 1275.030 3196.410 ;
        RECT 1273.300 3196.000 1273.580 3196.270 ;
        RECT 1274.750 3196.155 1275.030 3196.270 ;
        RECT 1586.630 788.955 1586.910 789.325 ;
        RECT 2704.430 788.955 2704.710 789.325 ;
        RECT 1586.700 787.965 1586.840 788.955 ;
        RECT 2028.700 788.645 2028.960 788.790 ;
        RECT 2076.540 788.645 2076.800 788.790 ;
        RECT 2028.690 788.275 2028.970 788.645 ;
        RECT 2076.530 788.275 2076.810 788.645 ;
        RECT 1393.430 787.595 1393.710 787.965 ;
        RECT 1586.630 787.595 1586.910 787.965 ;
        RECT 1877.350 787.595 1877.630 787.965 ;
        RECT 2283.530 787.850 2283.810 787.965 ;
        RECT 2284.450 787.850 2284.730 787.965 ;
        RECT 2283.530 787.710 2284.730 787.850 ;
        RECT 2283.530 787.595 2283.810 787.710 ;
        RECT 2284.450 787.595 2284.730 787.710 ;
        RECT 2572.870 787.595 2573.150 787.965 ;
        RECT 2632.210 787.595 2632.490 787.965 ;
        RECT 1393.500 787.285 1393.640 787.595 ;
        RECT 1393.430 786.915 1393.710 787.285 ;
        RECT 1877.420 786.605 1877.560 787.595 ;
        RECT 1877.350 786.235 1877.630 786.605 ;
        RECT 2572.940 785.925 2573.080 787.595 ;
        RECT 2632.280 787.430 2632.420 787.595 ;
        RECT 2608.300 787.285 2608.560 787.430 ;
        RECT 2608.290 786.915 2608.570 787.285 ;
        RECT 2632.220 787.110 2632.480 787.430 ;
        RECT 2704.500 787.285 2704.640 788.955 ;
        RECT 2801.030 788.275 2801.310 788.645 ;
        RECT 2704.430 786.915 2704.710 787.285 ;
        RECT 2801.100 786.605 2801.240 788.275 ;
        RECT 2863.130 787.595 2863.410 787.965 ;
        RECT 2863.200 787.170 2863.340 787.595 ;
        RECT 2863.590 787.170 2863.870 787.285 ;
        RECT 2863.200 787.030 2863.870 787.170 ;
        RECT 2863.590 786.915 2863.870 787.030 ;
        RECT 2801.030 786.235 2801.310 786.605 ;
        RECT 2572.870 785.555 2573.150 785.925 ;
      LAYER via2 ;
        RECT 1274.750 3196.200 1275.030 3196.480 ;
        RECT 1586.630 789.000 1586.910 789.280 ;
        RECT 2704.430 789.000 2704.710 789.280 ;
        RECT 2028.690 788.320 2028.970 788.600 ;
        RECT 2076.530 788.320 2076.810 788.600 ;
        RECT 1393.430 787.640 1393.710 787.920 ;
        RECT 1586.630 787.640 1586.910 787.920 ;
        RECT 1877.350 787.640 1877.630 787.920 ;
        RECT 2283.530 787.640 2283.810 787.920 ;
        RECT 2284.450 787.640 2284.730 787.920 ;
        RECT 2572.870 787.640 2573.150 787.920 ;
        RECT 2632.210 787.640 2632.490 787.920 ;
        RECT 1393.430 786.960 1393.710 787.240 ;
        RECT 1877.350 786.280 1877.630 786.560 ;
        RECT 2608.290 786.960 2608.570 787.240 ;
        RECT 2801.030 788.320 2801.310 788.600 ;
        RECT 2704.430 786.960 2704.710 787.240 ;
        RECT 2863.130 787.640 2863.410 787.920 ;
        RECT 2863.590 786.960 2863.870 787.240 ;
        RECT 2801.030 786.280 2801.310 786.560 ;
        RECT 2572.870 785.600 2573.150 785.880 ;
      LAYER met3 ;
        RECT 1274.725 3196.490 1275.055 3196.505 ;
        RECT 1275.390 3196.490 1275.770 3196.500 ;
        RECT 1274.725 3196.190 1275.770 3196.490 ;
        RECT 1274.725 3196.175 1275.055 3196.190 ;
        RECT 1275.390 3196.180 1275.770 3196.190 ;
        RECT 2917.600 792.010 2924.800 792.460 ;
        RECT 2916.710 791.710 2924.800 792.010 ;
        RECT 1538.510 789.290 1538.890 789.300 ;
        RECT 1586.605 789.290 1586.935 789.305 ;
        RECT 1538.510 788.990 1586.935 789.290 ;
        RECT 1538.510 788.980 1538.890 788.990 ;
        RECT 1586.605 788.975 1586.935 788.990 ;
        RECT 1924.910 789.290 1925.290 789.300 ;
        RECT 2510.030 789.290 2510.410 789.300 ;
        RECT 1924.910 788.990 1932.610 789.290 ;
        RECT 1924.910 788.980 1925.290 788.990 ;
        RECT 1932.310 788.610 1932.610 788.990 ;
        RECT 2476.030 788.990 2510.410 789.290 ;
        RECT 2028.665 788.610 2028.995 788.625 ;
        RECT 1462.190 788.310 1463.410 788.610 ;
        RECT 1275.390 787.930 1275.770 787.940 ;
        RECT 1393.405 787.930 1393.735 787.945 ;
        RECT 1275.390 787.630 1393.735 787.930 ;
        RECT 1275.390 787.620 1275.770 787.630 ;
        RECT 1393.405 787.615 1393.735 787.630 ;
        RECT 1393.405 787.250 1393.735 787.265 ;
        RECT 1462.190 787.250 1462.490 788.310 ;
        RECT 1463.110 787.930 1463.410 788.310 ;
        RECT 1665.510 788.310 1667.650 788.610 ;
        RECT 1497.110 787.930 1497.490 787.940 ;
        RECT 1463.110 787.630 1497.490 787.930 ;
        RECT 1497.110 787.620 1497.490 787.630 ;
        RECT 1586.605 787.930 1586.935 787.945 ;
        RECT 1586.605 787.630 1617.970 787.930 ;
        RECT 1586.605 787.615 1586.935 787.630 ;
        RECT 1393.405 786.950 1462.490 787.250 ;
        RECT 1497.110 787.250 1497.490 787.260 ;
        RECT 1538.510 787.250 1538.890 787.260 ;
        RECT 1497.110 786.950 1538.890 787.250 ;
        RECT 1617.670 787.250 1617.970 787.630 ;
        RECT 1665.510 787.250 1665.810 788.310 ;
        RECT 1667.350 787.930 1667.650 788.310 ;
        RECT 1702.310 788.310 1704.450 788.610 ;
        RECT 1932.310 788.310 2028.995 788.610 ;
        RECT 1702.310 787.930 1702.610 788.310 ;
        RECT 1667.350 787.630 1702.610 787.930 ;
        RECT 1704.150 787.930 1704.450 788.310 ;
        RECT 2028.665 788.295 2028.995 788.310 ;
        RECT 2076.505 788.610 2076.835 788.625 ;
        RECT 2089.630 788.610 2091.770 788.780 ;
        RECT 2076.505 788.480 2138.690 788.610 ;
        RECT 2076.505 788.310 2089.930 788.480 ;
        RECT 2091.470 788.310 2138.690 788.480 ;
        RECT 2076.505 788.295 2076.835 788.310 ;
        RECT 1877.325 787.930 1877.655 787.945 ;
        RECT 1704.150 787.630 1877.655 787.930 ;
        RECT 1877.325 787.615 1877.655 787.630 ;
        RECT 1617.670 786.950 1665.810 787.250 ;
        RECT 2138.390 787.250 2138.690 788.310 ;
        RECT 2139.310 788.310 2187.450 788.610 ;
        RECT 2139.310 787.250 2139.610 788.310 ;
        RECT 2138.390 786.950 2139.610 787.250 ;
        RECT 2187.150 787.250 2187.450 788.310 ;
        RECT 2283.505 787.930 2283.835 787.945 ;
        RECT 2235.910 787.630 2283.835 787.930 ;
        RECT 2235.910 787.250 2236.210 787.630 ;
        RECT 2283.505 787.615 2283.835 787.630 ;
        RECT 2284.425 787.930 2284.755 787.945 ;
        RECT 2476.030 787.930 2476.330 788.990 ;
        RECT 2510.030 788.980 2510.410 788.990 ;
        RECT 2656.310 789.290 2656.690 789.300 ;
        RECT 2704.405 789.290 2704.735 789.305 ;
        RECT 2656.310 788.990 2704.735 789.290 ;
        RECT 2656.310 788.980 2656.690 788.990 ;
        RECT 2704.405 788.975 2704.735 788.990 ;
        RECT 2801.005 788.610 2801.335 788.625 ;
        RECT 2801.005 788.310 2815.810 788.610 ;
        RECT 2801.005 788.295 2801.335 788.310 ;
        RECT 2572.845 787.930 2573.175 787.945 ;
        RECT 2284.425 787.630 2331.890 787.930 ;
        RECT 2284.425 787.615 2284.755 787.630 ;
        RECT 2187.150 786.950 2236.210 787.250 ;
        RECT 2331.590 787.250 2331.890 787.630 ;
        RECT 2332.510 787.630 2379.730 787.930 ;
        RECT 2332.510 787.250 2332.810 787.630 ;
        RECT 2331.590 786.950 2332.810 787.250 ;
        RECT 2379.430 787.250 2379.730 787.630 ;
        RECT 2429.110 787.630 2476.330 787.930 ;
        RECT 2525.710 787.630 2573.175 787.930 ;
        RECT 2429.110 787.250 2429.410 787.630 ;
        RECT 2379.430 786.950 2429.410 787.250 ;
        RECT 2510.950 787.250 2511.330 787.260 ;
        RECT 2525.710 787.250 2526.010 787.630 ;
        RECT 2572.845 787.615 2573.175 787.630 ;
        RECT 2632.185 787.930 2632.515 787.945 ;
        RECT 2656.310 787.930 2656.690 787.940 ;
        RECT 2752.910 787.930 2753.290 787.940 ;
        RECT 2632.185 787.630 2656.690 787.930 ;
        RECT 2632.185 787.615 2632.515 787.630 ;
        RECT 2656.310 787.620 2656.690 787.630 ;
        RECT 2718.910 787.630 2753.290 787.930 ;
        RECT 2608.265 787.250 2608.595 787.265 ;
        RECT 2510.950 786.950 2526.010 787.250 ;
        RECT 2607.590 786.950 2608.595 787.250 ;
        RECT 1393.405 786.935 1393.735 786.950 ;
        RECT 1497.110 786.940 1497.490 786.950 ;
        RECT 1538.510 786.940 1538.890 786.950 ;
        RECT 2510.950 786.940 2511.330 786.950 ;
        RECT 1877.325 786.570 1877.655 786.585 ;
        RECT 1923.990 786.570 1924.370 786.580 ;
        RECT 1877.325 786.270 1924.370 786.570 ;
        RECT 1877.325 786.255 1877.655 786.270 ;
        RECT 1923.990 786.260 1924.370 786.270 ;
        RECT 2572.845 785.890 2573.175 785.905 ;
        RECT 2607.590 785.890 2607.890 786.950 ;
        RECT 2608.265 786.935 2608.595 786.950 ;
        RECT 2704.405 787.250 2704.735 787.265 ;
        RECT 2718.910 787.250 2719.210 787.630 ;
        RECT 2752.910 787.620 2753.290 787.630 ;
        RECT 2704.405 786.950 2719.210 787.250 ;
        RECT 2815.510 787.250 2815.810 788.310 ;
        RECT 2863.105 787.930 2863.435 787.945 ;
        RECT 2916.710 787.930 2917.010 791.710 ;
        RECT 2917.600 791.260 2924.800 791.710 ;
        RECT 2849.550 787.630 2863.435 787.930 ;
        RECT 2849.550 787.250 2849.850 787.630 ;
        RECT 2863.105 787.615 2863.435 787.630 ;
        RECT 2884.510 787.630 2917.010 787.930 ;
        RECT 2815.510 786.950 2849.850 787.250 ;
        RECT 2863.565 787.250 2863.895 787.265 ;
        RECT 2884.510 787.250 2884.810 787.630 ;
        RECT 2863.565 786.950 2884.810 787.250 ;
        RECT 2704.405 786.935 2704.735 786.950 ;
        RECT 2863.565 786.935 2863.895 786.950 ;
        RECT 2752.910 786.570 2753.290 786.580 ;
        RECT 2801.005 786.570 2801.335 786.585 ;
        RECT 2752.910 786.270 2801.335 786.570 ;
        RECT 2752.910 786.260 2753.290 786.270 ;
        RECT 2801.005 786.255 2801.335 786.270 ;
        RECT 2572.845 785.590 2607.890 785.890 ;
        RECT 2572.845 785.575 2573.175 785.590 ;
      LAYER via3 ;
        RECT 1275.420 3196.180 1275.740 3196.500 ;
        RECT 1538.540 788.980 1538.860 789.300 ;
        RECT 1924.940 788.980 1925.260 789.300 ;
        RECT 1275.420 787.620 1275.740 787.940 ;
        RECT 1497.140 787.620 1497.460 787.940 ;
        RECT 1497.140 786.940 1497.460 787.260 ;
        RECT 1538.540 786.940 1538.860 787.260 ;
        RECT 2510.060 788.980 2510.380 789.300 ;
        RECT 2656.340 788.980 2656.660 789.300 ;
        RECT 2510.980 786.940 2511.300 787.260 ;
        RECT 2656.340 787.620 2656.660 787.940 ;
        RECT 1924.020 786.260 1924.340 786.580 ;
        RECT 2752.940 787.620 2753.260 787.940 ;
        RECT 2752.940 786.260 2753.260 786.580 ;
      LAYER met4 ;
        RECT 1275.415 3196.175 1275.745 3196.505 ;
        RECT 1275.430 787.945 1275.730 3196.175 ;
        RECT 1538.535 788.975 1538.865 789.305 ;
        RECT 1924.935 788.975 1925.265 789.305 ;
        RECT 2510.055 788.975 2510.385 789.305 ;
        RECT 2656.335 788.975 2656.665 789.305 ;
        RECT 1275.415 787.615 1275.745 787.945 ;
        RECT 1497.135 787.615 1497.465 787.945 ;
        RECT 1497.150 787.265 1497.450 787.615 ;
        RECT 1538.550 787.265 1538.850 788.975 ;
        RECT 1497.135 786.935 1497.465 787.265 ;
        RECT 1538.535 786.935 1538.865 787.265 ;
        RECT 1924.950 787.250 1925.250 788.975 ;
        RECT 1924.030 786.950 1925.250 787.250 ;
        RECT 2510.070 787.250 2510.370 788.975 ;
        RECT 2656.350 787.945 2656.650 788.975 ;
        RECT 2656.335 787.615 2656.665 787.945 ;
        RECT 2752.935 787.615 2753.265 787.945 ;
        RECT 2510.975 787.250 2511.305 787.265 ;
        RECT 2510.070 786.950 2511.305 787.250 ;
        RECT 1924.030 786.585 1924.330 786.950 ;
        RECT 2510.975 786.935 2511.305 786.950 ;
        RECT 2752.950 786.585 2753.250 787.615 ;
        RECT 1924.015 786.255 1924.345 786.585 ;
        RECT 2752.935 786.255 2753.265 786.585 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1683.670 1021.940 1683.990 1022.000 ;
        RECT 1690.570 1021.940 1690.890 1022.000 ;
        RECT 1683.670 1021.800 1690.890 1021.940 ;
        RECT 1683.670 1021.740 1683.990 1021.800 ;
        RECT 1690.570 1021.740 1690.890 1021.800 ;
        RECT 1875.950 1021.940 1876.270 1022.000 ;
        RECT 1924.710 1021.940 1925.030 1022.000 ;
        RECT 1875.950 1021.800 1925.030 1021.940 ;
        RECT 1875.950 1021.740 1876.270 1021.800 ;
        RECT 1924.710 1021.740 1925.030 1021.800 ;
        RECT 2125.270 1021.940 2125.590 1022.000 ;
        RECT 2172.650 1021.940 2172.970 1022.000 ;
        RECT 2125.270 1021.800 2172.970 1021.940 ;
        RECT 2125.270 1021.740 2125.590 1021.800 ;
        RECT 2172.650 1021.740 2172.970 1021.800 ;
        RECT 2608.270 1021.940 2608.590 1022.000 ;
        RECT 2632.190 1021.940 2632.510 1022.000 ;
        RECT 2608.270 1021.800 2632.510 1021.940 ;
        RECT 2608.270 1021.740 2608.590 1021.800 ;
        RECT 2632.190 1021.740 2632.510 1021.800 ;
      LAYER via ;
        RECT 1683.700 1021.740 1683.960 1022.000 ;
        RECT 1690.600 1021.740 1690.860 1022.000 ;
        RECT 1875.980 1021.740 1876.240 1022.000 ;
        RECT 1924.740 1021.740 1925.000 1022.000 ;
        RECT 2125.300 1021.740 2125.560 1022.000 ;
        RECT 2172.680 1021.740 2172.940 1022.000 ;
        RECT 2608.300 1021.740 2608.560 1022.000 ;
        RECT 2632.220 1021.740 2632.480 1022.000 ;
      LAYER met2 ;
        RECT 1312.860 3196.410 1313.140 3200.000 ;
        RECT 1314.310 3196.410 1314.590 3196.525 ;
        RECT 1312.860 3196.270 1314.590 3196.410 ;
        RECT 1312.860 3196.000 1313.140 3196.270 ;
        RECT 1314.310 3196.155 1314.590 3196.270 ;
        RECT 1393.430 1042.595 1393.710 1042.965 ;
        RECT 1393.500 1023.245 1393.640 1042.595 ;
        RECT 1449.090 1023.555 1449.370 1023.925 ;
        RECT 1504.750 1023.555 1505.030 1023.925 ;
        RECT 2704.430 1023.555 2704.710 1023.925 ;
        RECT 1393.430 1022.875 1393.710 1023.245 ;
        RECT 1449.160 1022.565 1449.300 1023.555 ;
        RECT 1449.090 1022.195 1449.370 1022.565 ;
        RECT 1504.820 1021.885 1504.960 1023.555 ;
        RECT 2172.670 1022.875 2172.950 1023.245 ;
        RECT 1875.970 1022.195 1876.250 1022.565 ;
        RECT 1924.730 1022.195 1925.010 1022.565 ;
        RECT 2090.330 1022.195 2090.610 1022.565 ;
        RECT 1876.040 1022.030 1876.180 1022.195 ;
        RECT 1924.800 1022.030 1924.940 1022.195 ;
        RECT 1683.700 1021.885 1683.960 1022.030 ;
        RECT 1690.600 1021.885 1690.860 1022.030 ;
        RECT 1504.750 1021.515 1505.030 1021.885 ;
        RECT 1683.690 1021.515 1683.970 1021.885 ;
        RECT 1690.590 1021.515 1690.870 1021.885 ;
        RECT 1875.980 1021.710 1876.240 1022.030 ;
        RECT 1924.740 1021.710 1925.000 1022.030 ;
        RECT 2090.400 1020.525 2090.540 1022.195 ;
        RECT 2172.740 1022.030 2172.880 1022.875 ;
        RECT 2572.870 1022.195 2573.150 1022.565 ;
        RECT 2632.210 1022.195 2632.490 1022.565 ;
        RECT 2125.300 1021.885 2125.560 1022.030 ;
        RECT 2125.290 1021.515 2125.570 1021.885 ;
        RECT 2172.680 1021.710 2172.940 1022.030 ;
        RECT 2572.940 1020.525 2573.080 1022.195 ;
        RECT 2632.280 1022.030 2632.420 1022.195 ;
        RECT 2608.300 1021.885 2608.560 1022.030 ;
        RECT 2608.290 1021.515 2608.570 1021.885 ;
        RECT 2632.220 1021.710 2632.480 1022.030 ;
        RECT 2704.500 1021.885 2704.640 1023.555 ;
        RECT 2801.030 1022.875 2801.310 1023.245 ;
        RECT 2704.430 1021.515 2704.710 1021.885 ;
        RECT 2801.100 1021.205 2801.240 1022.875 ;
        RECT 2863.130 1022.195 2863.410 1022.565 ;
        RECT 2863.200 1021.770 2863.340 1022.195 ;
        RECT 2863.590 1021.770 2863.870 1021.885 ;
        RECT 2863.200 1021.630 2863.870 1021.770 ;
        RECT 2863.590 1021.515 2863.870 1021.630 ;
        RECT 2801.030 1020.835 2801.310 1021.205 ;
        RECT 2090.330 1020.155 2090.610 1020.525 ;
        RECT 2572.870 1020.155 2573.150 1020.525 ;
      LAYER via2 ;
        RECT 1314.310 3196.200 1314.590 3196.480 ;
        RECT 1393.430 1042.640 1393.710 1042.920 ;
        RECT 1449.090 1023.600 1449.370 1023.880 ;
        RECT 1504.750 1023.600 1505.030 1023.880 ;
        RECT 2704.430 1023.600 2704.710 1023.880 ;
        RECT 1393.430 1022.920 1393.710 1023.200 ;
        RECT 1449.090 1022.240 1449.370 1022.520 ;
        RECT 2172.670 1022.920 2172.950 1023.200 ;
        RECT 1875.970 1022.240 1876.250 1022.520 ;
        RECT 1924.730 1022.240 1925.010 1022.520 ;
        RECT 2090.330 1022.240 2090.610 1022.520 ;
        RECT 1504.750 1021.560 1505.030 1021.840 ;
        RECT 1683.690 1021.560 1683.970 1021.840 ;
        RECT 1690.590 1021.560 1690.870 1021.840 ;
        RECT 2572.870 1022.240 2573.150 1022.520 ;
        RECT 2632.210 1022.240 2632.490 1022.520 ;
        RECT 2125.290 1021.560 2125.570 1021.840 ;
        RECT 2608.290 1021.560 2608.570 1021.840 ;
        RECT 2801.030 1022.920 2801.310 1023.200 ;
        RECT 2704.430 1021.560 2704.710 1021.840 ;
        RECT 2863.130 1022.240 2863.410 1022.520 ;
        RECT 2863.590 1021.560 2863.870 1021.840 ;
        RECT 2801.030 1020.880 2801.310 1021.160 ;
        RECT 2090.330 1020.200 2090.610 1020.480 ;
        RECT 2572.870 1020.200 2573.150 1020.480 ;
      LAYER met3 ;
        RECT 1314.285 3196.490 1314.615 3196.505 ;
        RECT 1316.790 3196.490 1317.170 3196.500 ;
        RECT 1314.285 3196.190 1317.170 3196.490 ;
        RECT 1314.285 3196.175 1314.615 3196.190 ;
        RECT 1316.790 3196.180 1317.170 3196.190 ;
        RECT 1316.790 1042.930 1317.170 1042.940 ;
        RECT 1393.405 1042.930 1393.735 1042.945 ;
        RECT 1316.790 1042.630 1393.735 1042.930 ;
        RECT 1316.790 1042.620 1317.170 1042.630 ;
        RECT 1393.405 1042.615 1393.735 1042.630 ;
        RECT 2917.600 1026.610 2924.800 1027.060 ;
        RECT 2916.710 1026.310 2924.800 1026.610 ;
        RECT 1449.065 1023.890 1449.395 1023.905 ;
        RECT 1504.725 1023.890 1505.055 1023.905 ;
        RECT 1449.065 1023.590 1505.055 1023.890 ;
        RECT 1449.065 1023.575 1449.395 1023.590 ;
        RECT 1504.725 1023.575 1505.055 1023.590 ;
        RECT 1814.510 1023.890 1814.890 1023.900 ;
        RECT 1862.350 1023.890 1862.730 1023.900 ;
        RECT 2316.830 1023.890 2317.210 1023.900 ;
        RECT 2510.030 1023.890 2510.410 1023.900 ;
        RECT 1814.510 1023.590 1862.730 1023.890 ;
        RECT 1814.510 1023.580 1814.890 1023.590 ;
        RECT 1862.350 1023.580 1862.730 1023.590 ;
        RECT 2282.830 1023.590 2317.210 1023.890 ;
        RECT 1393.405 1023.210 1393.735 1023.225 ;
        RECT 2172.645 1023.210 2172.975 1023.225 ;
        RECT 1393.405 1022.910 1424.770 1023.210 ;
        RECT 1393.405 1022.895 1393.735 1022.910 ;
        RECT 1424.470 1022.530 1424.770 1022.910 ;
        RECT 1558.790 1022.910 1617.970 1023.210 ;
        RECT 1449.065 1022.530 1449.395 1022.545 ;
        RECT 1424.470 1022.230 1449.395 1022.530 ;
        RECT 1449.065 1022.215 1449.395 1022.230 ;
        RECT 1504.725 1021.850 1505.055 1021.865 ;
        RECT 1558.790 1021.850 1559.090 1022.910 ;
        RECT 1617.670 1022.530 1617.970 1022.910 ;
        RECT 1932.310 1022.910 1994.250 1023.210 ;
        RECT 1814.510 1022.530 1814.890 1022.540 ;
        RECT 1617.670 1022.230 1642.810 1022.530 ;
        RECT 1504.725 1021.550 1559.090 1021.850 ;
        RECT 1642.510 1021.850 1642.810 1022.230 ;
        RECT 1732.900 1022.230 1814.890 1022.530 ;
        RECT 1683.665 1021.850 1683.995 1021.865 ;
        RECT 1642.510 1021.550 1683.995 1021.850 ;
        RECT 1504.725 1021.535 1505.055 1021.550 ;
        RECT 1683.665 1021.535 1683.995 1021.550 ;
        RECT 1690.565 1021.850 1690.895 1021.865 ;
        RECT 1732.900 1021.850 1733.200 1022.230 ;
        RECT 1814.510 1022.220 1814.890 1022.230 ;
        RECT 1862.350 1022.530 1862.730 1022.540 ;
        RECT 1875.945 1022.530 1876.275 1022.545 ;
        RECT 1862.350 1022.230 1876.275 1022.530 ;
        RECT 1862.350 1022.220 1862.730 1022.230 ;
        RECT 1875.945 1022.215 1876.275 1022.230 ;
        RECT 1924.705 1022.530 1925.035 1022.545 ;
        RECT 1932.310 1022.530 1932.610 1022.910 ;
        RECT 1924.705 1022.230 1932.610 1022.530 ;
        RECT 1924.705 1022.215 1925.035 1022.230 ;
        RECT 1690.565 1021.550 1733.200 1021.850 ;
        RECT 1993.950 1021.850 1994.250 1022.910 ;
        RECT 2172.645 1022.910 2187.450 1023.210 ;
        RECT 2172.645 1022.895 2172.975 1022.910 ;
        RECT 2090.305 1022.530 2090.635 1022.545 ;
        RECT 2042.710 1022.230 2090.635 1022.530 ;
        RECT 2042.710 1021.850 2043.010 1022.230 ;
        RECT 2090.305 1022.215 2090.635 1022.230 ;
        RECT 2125.265 1021.850 2125.595 1021.865 ;
        RECT 1993.950 1021.550 2043.010 1021.850 ;
        RECT 2124.590 1021.550 2125.595 1021.850 ;
        RECT 2187.150 1021.850 2187.450 1022.910 ;
        RECT 2282.830 1022.530 2283.130 1023.590 ;
        RECT 2316.830 1023.580 2317.210 1023.590 ;
        RECT 2476.030 1023.590 2510.410 1023.890 ;
        RECT 2476.030 1022.530 2476.330 1023.590 ;
        RECT 2510.030 1023.580 2510.410 1023.590 ;
        RECT 2656.310 1023.890 2656.690 1023.900 ;
        RECT 2704.405 1023.890 2704.735 1023.905 ;
        RECT 2656.310 1023.590 2704.735 1023.890 ;
        RECT 2656.310 1023.580 2656.690 1023.590 ;
        RECT 2704.405 1023.575 2704.735 1023.590 ;
        RECT 2801.005 1023.210 2801.335 1023.225 ;
        RECT 2801.005 1022.910 2815.810 1023.210 ;
        RECT 2801.005 1022.895 2801.335 1022.910 ;
        RECT 2572.845 1022.530 2573.175 1022.545 ;
        RECT 2235.910 1022.230 2283.130 1022.530 ;
        RECT 2332.510 1022.230 2414.690 1022.530 ;
        RECT 2235.910 1021.850 2236.210 1022.230 ;
        RECT 2187.150 1021.550 2236.210 1021.850 ;
        RECT 2317.750 1021.850 2318.130 1021.860 ;
        RECT 2332.510 1021.850 2332.810 1022.230 ;
        RECT 2317.750 1021.550 2332.810 1021.850 ;
        RECT 2414.390 1021.850 2414.690 1022.230 ;
        RECT 2429.110 1022.230 2476.330 1022.530 ;
        RECT 2525.710 1022.230 2573.175 1022.530 ;
        RECT 2429.110 1021.850 2429.410 1022.230 ;
        RECT 2414.390 1021.550 2429.410 1021.850 ;
        RECT 2510.950 1021.850 2511.330 1021.860 ;
        RECT 2525.710 1021.850 2526.010 1022.230 ;
        RECT 2572.845 1022.215 2573.175 1022.230 ;
        RECT 2632.185 1022.530 2632.515 1022.545 ;
        RECT 2656.310 1022.530 2656.690 1022.540 ;
        RECT 2752.910 1022.530 2753.290 1022.540 ;
        RECT 2632.185 1022.230 2656.690 1022.530 ;
        RECT 2632.185 1022.215 2632.515 1022.230 ;
        RECT 2656.310 1022.220 2656.690 1022.230 ;
        RECT 2718.910 1022.230 2753.290 1022.530 ;
        RECT 2608.265 1021.850 2608.595 1021.865 ;
        RECT 2510.950 1021.550 2526.010 1021.850 ;
        RECT 2607.590 1021.550 2608.595 1021.850 ;
        RECT 1690.565 1021.535 1690.895 1021.550 ;
        RECT 2090.305 1020.490 2090.635 1020.505 ;
        RECT 2124.590 1020.490 2124.890 1021.550 ;
        RECT 2125.265 1021.535 2125.595 1021.550 ;
        RECT 2317.750 1021.540 2318.130 1021.550 ;
        RECT 2510.950 1021.540 2511.330 1021.550 ;
        RECT 2090.305 1020.190 2124.890 1020.490 ;
        RECT 2572.845 1020.490 2573.175 1020.505 ;
        RECT 2607.590 1020.490 2607.890 1021.550 ;
        RECT 2608.265 1021.535 2608.595 1021.550 ;
        RECT 2704.405 1021.850 2704.735 1021.865 ;
        RECT 2718.910 1021.850 2719.210 1022.230 ;
        RECT 2752.910 1022.220 2753.290 1022.230 ;
        RECT 2704.405 1021.550 2719.210 1021.850 ;
        RECT 2815.510 1021.850 2815.810 1022.910 ;
        RECT 2863.105 1022.530 2863.435 1022.545 ;
        RECT 2916.710 1022.530 2917.010 1026.310 ;
        RECT 2917.600 1025.860 2924.800 1026.310 ;
        RECT 2849.550 1022.230 2863.435 1022.530 ;
        RECT 2849.550 1021.850 2849.850 1022.230 ;
        RECT 2863.105 1022.215 2863.435 1022.230 ;
        RECT 2884.510 1022.230 2917.010 1022.530 ;
        RECT 2815.510 1021.550 2849.850 1021.850 ;
        RECT 2863.565 1021.850 2863.895 1021.865 ;
        RECT 2884.510 1021.850 2884.810 1022.230 ;
        RECT 2863.565 1021.550 2884.810 1021.850 ;
        RECT 2704.405 1021.535 2704.735 1021.550 ;
        RECT 2863.565 1021.535 2863.895 1021.550 ;
        RECT 2752.910 1021.170 2753.290 1021.180 ;
        RECT 2801.005 1021.170 2801.335 1021.185 ;
        RECT 2752.910 1020.870 2801.335 1021.170 ;
        RECT 2752.910 1020.860 2753.290 1020.870 ;
        RECT 2801.005 1020.855 2801.335 1020.870 ;
        RECT 2572.845 1020.190 2607.890 1020.490 ;
        RECT 2090.305 1020.175 2090.635 1020.190 ;
        RECT 2572.845 1020.175 2573.175 1020.190 ;
      LAYER via3 ;
        RECT 1316.820 3196.180 1317.140 3196.500 ;
        RECT 1316.820 1042.620 1317.140 1042.940 ;
        RECT 1814.540 1023.580 1814.860 1023.900 ;
        RECT 1862.380 1023.580 1862.700 1023.900 ;
        RECT 1814.540 1022.220 1814.860 1022.540 ;
        RECT 1862.380 1022.220 1862.700 1022.540 ;
        RECT 2316.860 1023.580 2317.180 1023.900 ;
        RECT 2510.060 1023.580 2510.380 1023.900 ;
        RECT 2656.340 1023.580 2656.660 1023.900 ;
        RECT 2317.780 1021.540 2318.100 1021.860 ;
        RECT 2510.980 1021.540 2511.300 1021.860 ;
        RECT 2656.340 1022.220 2656.660 1022.540 ;
        RECT 2752.940 1022.220 2753.260 1022.540 ;
        RECT 2752.940 1020.860 2753.260 1021.180 ;
      LAYER met4 ;
        RECT 1316.815 3196.175 1317.145 3196.505 ;
        RECT 1316.830 1042.945 1317.130 3196.175 ;
        RECT 1316.815 1042.615 1317.145 1042.945 ;
        RECT 1814.535 1023.575 1814.865 1023.905 ;
        RECT 1862.375 1023.575 1862.705 1023.905 ;
        RECT 2316.855 1023.575 2317.185 1023.905 ;
        RECT 2510.055 1023.575 2510.385 1023.905 ;
        RECT 2656.335 1023.575 2656.665 1023.905 ;
        RECT 1814.550 1022.545 1814.850 1023.575 ;
        RECT 1862.390 1022.545 1862.690 1023.575 ;
        RECT 1814.535 1022.215 1814.865 1022.545 ;
        RECT 1862.375 1022.215 1862.705 1022.545 ;
        RECT 2316.870 1021.850 2317.170 1023.575 ;
        RECT 2317.775 1021.850 2318.105 1021.865 ;
        RECT 2316.870 1021.550 2318.105 1021.850 ;
        RECT 2510.070 1021.850 2510.370 1023.575 ;
        RECT 2656.350 1022.545 2656.650 1023.575 ;
        RECT 2656.335 1022.215 2656.665 1022.545 ;
        RECT 2752.935 1022.215 2753.265 1022.545 ;
        RECT 2510.975 1021.850 2511.305 1021.865 ;
        RECT 2510.070 1021.550 2511.305 1021.850 ;
        RECT 2317.775 1021.535 2318.105 1021.550 ;
        RECT 2510.975 1021.535 2511.305 1021.550 ;
        RECT 2752.950 1021.185 2753.250 1022.215 ;
        RECT 2752.935 1020.855 2753.265 1021.185 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1352.470 3213.580 1352.790 3213.640 ;
        RECT 2902.210 3213.580 2902.530 3213.640 ;
        RECT 1352.470 3213.440 2902.530 3213.580 ;
        RECT 1352.470 3213.380 1352.790 3213.440 ;
        RECT 2902.210 3213.380 2902.530 3213.440 ;
      LAYER via ;
        RECT 1352.500 3213.380 1352.760 3213.640 ;
        RECT 2902.240 3213.380 2902.500 3213.640 ;
      LAYER met2 ;
        RECT 1352.500 3213.350 1352.760 3213.670 ;
        RECT 2902.240 3213.350 2902.500 3213.670 ;
        RECT 1352.560 3200.000 1352.700 3213.350 ;
        RECT 1352.420 3196.000 1352.700 3200.000 ;
        RECT 2902.300 1261.245 2902.440 3213.350 ;
        RECT 2902.230 1260.875 2902.510 1261.245 ;
      LAYER via2 ;
        RECT 2902.230 1260.920 2902.510 1261.200 ;
      LAYER met3 ;
        RECT 2902.205 1261.210 2902.535 1261.225 ;
        RECT 2917.600 1261.210 2924.800 1261.660 ;
        RECT 2902.205 1260.910 2924.800 1261.210 ;
        RECT 2902.205 1260.895 2902.535 1260.910 ;
        RECT 2917.600 1260.460 2924.800 1260.910 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1391.570 3204.060 1391.890 3204.120 ;
        RECT 2652.890 3204.060 2653.210 3204.120 ;
        RECT 1391.570 3203.920 2653.210 3204.060 ;
        RECT 1391.570 3203.860 1391.890 3203.920 ;
        RECT 2652.890 3203.860 2653.210 3203.920 ;
        RECT 2652.890 1497.260 2653.210 1497.320 ;
        RECT 2898.530 1497.260 2898.850 1497.320 ;
        RECT 2652.890 1497.120 2898.850 1497.260 ;
        RECT 2652.890 1497.060 2653.210 1497.120 ;
        RECT 2898.530 1497.060 2898.850 1497.120 ;
      LAYER via ;
        RECT 1391.600 3203.860 1391.860 3204.120 ;
        RECT 2652.920 3203.860 2653.180 3204.120 ;
        RECT 2652.920 1497.060 2653.180 1497.320 ;
        RECT 2898.560 1497.060 2898.820 1497.320 ;
      LAYER met2 ;
        RECT 1391.600 3203.830 1391.860 3204.150 ;
        RECT 2652.920 3203.830 2653.180 3204.150 ;
        RECT 1391.660 3200.000 1391.800 3203.830 ;
        RECT 1391.520 3196.000 1391.800 3200.000 ;
        RECT 2652.980 1497.350 2653.120 3203.830 ;
        RECT 2652.920 1497.030 2653.180 1497.350 ;
        RECT 2898.560 1497.030 2898.820 1497.350 ;
        RECT 2898.620 1495.845 2898.760 1497.030 ;
        RECT 2898.550 1495.475 2898.830 1495.845 ;
      LAYER via2 ;
        RECT 2898.550 1495.520 2898.830 1495.800 ;
      LAYER met3 ;
        RECT 2898.525 1495.810 2898.855 1495.825 ;
        RECT 2917.600 1495.810 2924.800 1496.260 ;
        RECT 2898.525 1495.510 2924.800 1495.810 ;
        RECT 2898.525 1495.495 2898.855 1495.510 ;
        RECT 2917.600 1495.060 2924.800 1495.510 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1431.130 3204.400 1431.450 3204.460 ;
        RECT 2647.370 3204.400 2647.690 3204.460 ;
        RECT 1431.130 3204.260 2647.690 3204.400 ;
        RECT 1431.130 3204.200 1431.450 3204.260 ;
        RECT 2647.370 3204.200 2647.690 3204.260 ;
        RECT 2648.290 1731.860 2648.610 1731.920 ;
        RECT 2900.830 1731.860 2901.150 1731.920 ;
        RECT 2648.290 1731.720 2901.150 1731.860 ;
        RECT 2648.290 1731.660 2648.610 1731.720 ;
        RECT 2900.830 1731.660 2901.150 1731.720 ;
      LAYER via ;
        RECT 1431.160 3204.200 1431.420 3204.460 ;
        RECT 2647.400 3204.200 2647.660 3204.460 ;
        RECT 2648.320 1731.660 2648.580 1731.920 ;
        RECT 2900.860 1731.660 2901.120 1731.920 ;
      LAYER met2 ;
        RECT 1431.160 3204.170 1431.420 3204.490 ;
        RECT 2647.400 3204.170 2647.660 3204.490 ;
        RECT 1431.220 3200.000 1431.360 3204.170 ;
        RECT 1431.080 3196.000 1431.360 3200.000 ;
        RECT 2647.460 1731.690 2647.600 3204.170 ;
        RECT 2648.320 1731.690 2648.580 1731.950 ;
        RECT 2647.460 1731.630 2648.580 1731.690 ;
        RECT 2900.860 1731.630 2901.120 1731.950 ;
        RECT 2647.460 1731.550 2648.520 1731.630 ;
        RECT 2900.920 1730.445 2901.060 1731.630 ;
        RECT 2900.850 1730.075 2901.130 1730.445 ;
      LAYER via2 ;
        RECT 2900.850 1730.120 2901.130 1730.400 ;
      LAYER met3 ;
        RECT 2900.825 1730.410 2901.155 1730.425 ;
        RECT 2917.600 1730.410 2924.800 1730.860 ;
        RECT 2900.825 1730.110 2924.800 1730.410 ;
        RECT 2900.825 1730.095 2901.155 1730.110 ;
        RECT 2917.600 1729.660 2924.800 1730.110 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1470.690 3204.740 1471.010 3204.800 ;
        RECT 2647.830 3204.740 2648.150 3204.800 ;
        RECT 1470.690 3204.600 2648.150 3204.740 ;
        RECT 1470.690 3204.540 1471.010 3204.600 ;
        RECT 2647.830 3204.540 2648.150 3204.600 ;
        RECT 2647.830 1966.460 2648.150 1966.520 ;
        RECT 2898.070 1966.460 2898.390 1966.520 ;
        RECT 2647.830 1966.320 2898.390 1966.460 ;
        RECT 2647.830 1966.260 2648.150 1966.320 ;
        RECT 2898.070 1966.260 2898.390 1966.320 ;
      LAYER via ;
        RECT 1470.720 3204.540 1470.980 3204.800 ;
        RECT 2647.860 3204.540 2648.120 3204.800 ;
        RECT 2647.860 1966.260 2648.120 1966.520 ;
        RECT 2898.100 1966.260 2898.360 1966.520 ;
      LAYER met2 ;
        RECT 1470.720 3204.510 1470.980 3204.830 ;
        RECT 2647.860 3204.510 2648.120 3204.830 ;
        RECT 1470.780 3200.000 1470.920 3204.510 ;
        RECT 1470.640 3196.000 1470.920 3200.000 ;
        RECT 2647.920 1966.550 2648.060 3204.510 ;
        RECT 2647.860 1966.230 2648.120 1966.550 ;
        RECT 2898.100 1966.230 2898.360 1966.550 ;
        RECT 2898.160 1965.045 2898.300 1966.230 ;
        RECT 2898.090 1964.675 2898.370 1965.045 ;
      LAYER via2 ;
        RECT 2898.090 1964.720 2898.370 1965.000 ;
      LAYER met3 ;
        RECT 2898.065 1965.010 2898.395 1965.025 ;
        RECT 2917.600 1965.010 2924.800 1965.460 ;
        RECT 2898.065 1964.710 2924.800 1965.010 ;
        RECT 2898.065 1964.695 2898.395 1964.710 ;
        RECT 2917.600 1964.260 2924.800 1964.710 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1510.250 3205.080 1510.570 3205.140 ;
        RECT 2654.270 3205.080 2654.590 3205.140 ;
        RECT 1510.250 3204.940 2654.590 3205.080 ;
        RECT 1510.250 3204.880 1510.570 3204.940 ;
        RECT 2654.270 3204.880 2654.590 3204.940 ;
        RECT 2654.270 2201.060 2654.590 2201.120 ;
        RECT 2900.830 2201.060 2901.150 2201.120 ;
        RECT 2654.270 2200.920 2901.150 2201.060 ;
        RECT 2654.270 2200.860 2654.590 2200.920 ;
        RECT 2900.830 2200.860 2901.150 2200.920 ;
      LAYER via ;
        RECT 1510.280 3204.880 1510.540 3205.140 ;
        RECT 2654.300 3204.880 2654.560 3205.140 ;
        RECT 2654.300 2200.860 2654.560 2201.120 ;
        RECT 2900.860 2200.860 2901.120 2201.120 ;
      LAYER met2 ;
        RECT 1510.280 3204.850 1510.540 3205.170 ;
        RECT 2654.300 3204.850 2654.560 3205.170 ;
        RECT 1510.340 3200.000 1510.480 3204.850 ;
        RECT 1510.200 3196.000 1510.480 3200.000 ;
        RECT 2654.360 2201.150 2654.500 3204.850 ;
        RECT 2654.300 2200.830 2654.560 2201.150 ;
        RECT 2900.860 2200.830 2901.120 2201.150 ;
        RECT 2900.920 2199.645 2901.060 2200.830 ;
        RECT 2900.850 2199.275 2901.130 2199.645 ;
      LAYER via2 ;
        RECT 2900.850 2199.320 2901.130 2199.600 ;
      LAYER met3 ;
        RECT 2900.825 2199.610 2901.155 2199.625 ;
        RECT 2917.600 2199.610 2924.800 2200.060 ;
        RECT 2900.825 2199.310 2924.800 2199.610 ;
        RECT 2900.825 2199.295 2901.155 2199.310 ;
        RECT 2917.600 2198.860 2924.800 2199.310 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1338.670 201.860 1338.990 201.920 ;
        RECT 1386.510 201.860 1386.830 201.920 ;
        RECT 1338.670 201.720 1386.830 201.860 ;
        RECT 1338.670 201.660 1338.990 201.720 ;
        RECT 1386.510 201.660 1386.830 201.720 ;
        RECT 2014.870 201.860 2015.190 201.920 ;
        RECT 2062.250 201.860 2062.570 201.920 ;
        RECT 2014.870 201.720 2062.570 201.860 ;
        RECT 2014.870 201.660 2015.190 201.720 ;
        RECT 2062.250 201.660 2062.570 201.720 ;
        RECT 1559.010 200.500 1559.330 200.560 ;
        RECT 1586.610 200.500 1586.930 200.560 ;
        RECT 1559.010 200.360 1586.930 200.500 ;
        RECT 1559.010 200.300 1559.330 200.360 ;
        RECT 1586.610 200.300 1586.930 200.360 ;
        RECT 2608.270 200.500 2608.590 200.560 ;
        RECT 2632.190 200.500 2632.510 200.560 ;
        RECT 2608.270 200.360 2632.510 200.500 ;
        RECT 2608.270 200.300 2608.590 200.360 ;
        RECT 2632.190 200.300 2632.510 200.360 ;
      LAYER via ;
        RECT 1338.700 201.660 1338.960 201.920 ;
        RECT 1386.540 201.660 1386.800 201.920 ;
        RECT 2014.900 201.660 2015.160 201.920 ;
        RECT 2062.280 201.660 2062.540 201.920 ;
        RECT 1559.040 200.300 1559.300 200.560 ;
        RECT 1586.640 200.300 1586.900 200.560 ;
        RECT 2608.300 200.300 2608.560 200.560 ;
        RECT 2632.220 200.300 2632.480 200.560 ;
      LAYER met2 ;
        RECT 1167.960 3196.410 1168.240 3200.000 ;
        RECT 1169.870 3196.410 1170.150 3196.525 ;
        RECT 1167.960 3196.270 1170.150 3196.410 ;
        RECT 1167.960 3196.000 1168.240 3196.270 ;
        RECT 1169.870 3196.155 1170.150 3196.270 ;
        RECT 1171.710 1682.475 1171.990 1682.845 ;
        RECT 1171.780 1635.925 1171.920 1682.475 ;
        RECT 1171.710 1635.555 1171.990 1635.925 ;
        RECT 1171.250 1515.195 1171.530 1515.565 ;
        RECT 1171.320 1498.565 1171.460 1515.195 ;
        RECT 1171.250 1498.195 1171.530 1498.565 ;
        RECT 1169.870 1309.835 1170.150 1310.205 ;
        RECT 1169.940 1263.285 1170.080 1309.835 ;
        RECT 1169.870 1262.915 1170.150 1263.285 ;
        RECT 1171.710 1034.435 1171.990 1034.805 ;
        RECT 1171.780 987.885 1171.920 1034.435 ;
        RECT 1171.710 987.515 1171.990 987.885 ;
        RECT 1172.630 937.195 1172.910 937.565 ;
        RECT 1172.700 890.645 1172.840 937.195 ;
        RECT 1172.630 890.275 1172.910 890.645 ;
        RECT 1171.710 693.075 1171.990 693.445 ;
        RECT 1171.780 609.125 1171.920 693.075 ;
        RECT 1171.710 608.755 1171.990 609.125 ;
        RECT 1173.550 606.715 1173.830 607.085 ;
        RECT 1173.620 564.925 1173.760 606.715 ;
        RECT 1173.550 564.555 1173.830 564.925 ;
        RECT 1200.230 219.115 1200.510 219.485 ;
        RECT 1200.300 201.125 1200.440 219.115 ;
        RECT 1749.010 202.115 1749.290 202.485 ;
        RECT 2062.270 202.115 2062.550 202.485 ;
        RECT 2069.630 202.115 2069.910 202.485 ;
        RECT 2704.430 202.115 2704.710 202.485 ;
        RECT 1338.700 201.805 1338.960 201.950 ;
        RECT 1386.540 201.805 1386.800 201.950 ;
        RECT 1338.690 201.435 1338.970 201.805 ;
        RECT 1386.530 201.435 1386.810 201.805 ;
        RECT 1393.430 201.435 1393.710 201.805 ;
        RECT 1200.230 200.755 1200.510 201.125 ;
        RECT 1393.500 200.445 1393.640 201.435 ;
        RECT 1749.080 201.125 1749.220 202.115 ;
        RECT 2062.340 201.950 2062.480 202.115 ;
        RECT 2014.900 201.805 2015.160 201.950 ;
        RECT 2014.890 201.435 2015.170 201.805 ;
        RECT 2062.280 201.630 2062.540 201.950 ;
        RECT 2069.700 201.125 2069.840 202.115 ;
        RECT 1586.630 200.755 1586.910 201.125 ;
        RECT 1634.010 200.755 1634.290 201.125 ;
        RECT 1705.310 200.755 1705.590 201.125 ;
        RECT 1749.010 200.755 1749.290 201.125 ;
        RECT 1917.830 200.755 1918.110 201.125 ;
        RECT 2069.630 200.755 2069.910 201.125 ;
        RECT 2283.530 201.010 2283.810 201.125 ;
        RECT 2284.450 201.010 2284.730 201.125 ;
        RECT 2283.530 200.870 2284.730 201.010 ;
        RECT 2283.530 200.755 2283.810 200.870 ;
        RECT 2284.450 200.755 2284.730 200.870 ;
        RECT 2572.870 200.755 2573.150 201.125 ;
        RECT 2632.210 200.755 2632.490 201.125 ;
        RECT 1586.700 200.590 1586.840 200.755 ;
        RECT 1559.040 200.445 1559.300 200.590 ;
        RECT 1393.430 200.075 1393.710 200.445 ;
        RECT 1559.030 200.075 1559.310 200.445 ;
        RECT 1586.640 200.270 1586.900 200.590 ;
        RECT 1634.080 200.330 1634.220 200.755 ;
        RECT 1634.930 200.330 1635.210 200.445 ;
        RECT 1634.080 200.190 1635.210 200.330 ;
        RECT 1634.930 200.075 1635.210 200.190 ;
        RECT 1705.380 199.085 1705.520 200.755 ;
        RECT 1917.900 200.445 1918.040 200.755 ;
        RECT 1917.830 200.075 1918.110 200.445 ;
        RECT 2572.940 199.085 2573.080 200.755 ;
        RECT 2632.280 200.590 2632.420 200.755 ;
        RECT 2608.300 200.445 2608.560 200.590 ;
        RECT 2608.290 200.075 2608.570 200.445 ;
        RECT 2632.220 200.270 2632.480 200.590 ;
        RECT 2704.500 200.445 2704.640 202.115 ;
        RECT 2801.030 201.435 2801.310 201.805 ;
        RECT 2704.430 200.075 2704.710 200.445 ;
        RECT 2801.100 199.765 2801.240 201.435 ;
        RECT 2863.130 200.755 2863.410 201.125 ;
        RECT 2863.200 200.330 2863.340 200.755 ;
        RECT 2863.590 200.330 2863.870 200.445 ;
        RECT 2863.200 200.190 2863.870 200.330 ;
        RECT 2863.590 200.075 2863.870 200.190 ;
        RECT 2801.030 199.395 2801.310 199.765 ;
        RECT 1705.310 198.715 1705.590 199.085 ;
        RECT 2572.870 198.715 2573.150 199.085 ;
      LAYER via2 ;
        RECT 1169.870 3196.200 1170.150 3196.480 ;
        RECT 1171.710 1682.520 1171.990 1682.800 ;
        RECT 1171.710 1635.600 1171.990 1635.880 ;
        RECT 1171.250 1515.240 1171.530 1515.520 ;
        RECT 1171.250 1498.240 1171.530 1498.520 ;
        RECT 1169.870 1309.880 1170.150 1310.160 ;
        RECT 1169.870 1262.960 1170.150 1263.240 ;
        RECT 1171.710 1034.480 1171.990 1034.760 ;
        RECT 1171.710 987.560 1171.990 987.840 ;
        RECT 1172.630 937.240 1172.910 937.520 ;
        RECT 1172.630 890.320 1172.910 890.600 ;
        RECT 1171.710 693.120 1171.990 693.400 ;
        RECT 1171.710 608.800 1171.990 609.080 ;
        RECT 1173.550 606.760 1173.830 607.040 ;
        RECT 1173.550 564.600 1173.830 564.880 ;
        RECT 1200.230 219.160 1200.510 219.440 ;
        RECT 1749.010 202.160 1749.290 202.440 ;
        RECT 2062.270 202.160 2062.550 202.440 ;
        RECT 2069.630 202.160 2069.910 202.440 ;
        RECT 2704.430 202.160 2704.710 202.440 ;
        RECT 1338.690 201.480 1338.970 201.760 ;
        RECT 1386.530 201.480 1386.810 201.760 ;
        RECT 1393.430 201.480 1393.710 201.760 ;
        RECT 1200.230 200.800 1200.510 201.080 ;
        RECT 2014.890 201.480 2015.170 201.760 ;
        RECT 1586.630 200.800 1586.910 201.080 ;
        RECT 1634.010 200.800 1634.290 201.080 ;
        RECT 1705.310 200.800 1705.590 201.080 ;
        RECT 1749.010 200.800 1749.290 201.080 ;
        RECT 1917.830 200.800 1918.110 201.080 ;
        RECT 2069.630 200.800 2069.910 201.080 ;
        RECT 2283.530 200.800 2283.810 201.080 ;
        RECT 2284.450 200.800 2284.730 201.080 ;
        RECT 2572.870 200.800 2573.150 201.080 ;
        RECT 2632.210 200.800 2632.490 201.080 ;
        RECT 1393.430 200.120 1393.710 200.400 ;
        RECT 1559.030 200.120 1559.310 200.400 ;
        RECT 1634.930 200.120 1635.210 200.400 ;
        RECT 1917.830 200.120 1918.110 200.400 ;
        RECT 2608.290 200.120 2608.570 200.400 ;
        RECT 2801.030 201.480 2801.310 201.760 ;
        RECT 2704.430 200.120 2704.710 200.400 ;
        RECT 2863.130 200.800 2863.410 201.080 ;
        RECT 2863.590 200.120 2863.870 200.400 ;
        RECT 2801.030 199.440 2801.310 199.720 ;
        RECT 1705.310 198.760 1705.590 199.040 ;
        RECT 2572.870 198.760 2573.150 199.040 ;
      LAYER met3 ;
        RECT 1169.845 3196.490 1170.175 3196.505 ;
        RECT 1172.350 3196.490 1172.730 3196.500 ;
        RECT 1169.845 3196.190 1172.730 3196.490 ;
        RECT 1169.845 3196.175 1170.175 3196.190 ;
        RECT 1172.350 3196.180 1172.730 3196.190 ;
        RECT 1171.430 1683.180 1171.810 1683.500 ;
        RECT 1171.470 1682.825 1171.770 1683.180 ;
        RECT 1171.470 1682.510 1172.015 1682.825 ;
        RECT 1171.685 1682.495 1172.015 1682.510 ;
        RECT 1171.685 1635.890 1172.015 1635.905 ;
        RECT 1173.270 1635.890 1173.650 1635.900 ;
        RECT 1171.685 1635.590 1173.650 1635.890 ;
        RECT 1171.685 1635.575 1172.015 1635.590 ;
        RECT 1173.270 1635.580 1173.650 1635.590 ;
        RECT 1173.270 1595.090 1173.650 1595.100 ;
        RECT 1171.470 1594.790 1173.650 1595.090 ;
        RECT 1171.470 1594.420 1171.770 1594.790 ;
        RECT 1173.270 1594.780 1173.650 1594.790 ;
        RECT 1171.430 1594.100 1171.810 1594.420 ;
        RECT 1171.225 1515.540 1171.555 1515.545 ;
        RECT 1171.225 1515.530 1171.810 1515.540 ;
        RECT 1171.000 1515.230 1171.810 1515.530 ;
        RECT 1171.225 1515.220 1171.810 1515.230 ;
        RECT 1171.225 1515.215 1171.555 1515.220 ;
        RECT 1171.225 1498.530 1171.555 1498.545 ;
        RECT 1171.225 1498.215 1171.770 1498.530 ;
        RECT 1171.470 1497.860 1171.770 1498.215 ;
        RECT 1171.430 1497.540 1171.810 1497.860 ;
        RECT 1171.430 1452.290 1171.810 1452.300 ;
        RECT 1173.270 1452.290 1173.650 1452.300 ;
        RECT 1171.430 1451.990 1173.650 1452.290 ;
        RECT 1171.430 1451.980 1171.810 1451.990 ;
        RECT 1173.270 1451.980 1173.650 1451.990 ;
        RECT 1172.350 1367.290 1172.730 1367.300 ;
        RECT 1170.550 1366.990 1172.730 1367.290 ;
        RECT 1170.550 1366.620 1170.850 1366.990 ;
        RECT 1172.350 1366.980 1172.730 1366.990 ;
        RECT 1170.510 1366.300 1170.890 1366.620 ;
        RECT 1170.510 1319.010 1170.890 1319.020 ;
        RECT 1169.630 1318.710 1170.890 1319.010 ;
        RECT 1169.630 1317.660 1169.930 1318.710 ;
        RECT 1170.510 1318.700 1170.890 1318.710 ;
        RECT 1169.590 1317.340 1169.970 1317.660 ;
        RECT 1169.590 1310.540 1169.970 1310.860 ;
        RECT 1169.630 1310.185 1169.930 1310.540 ;
        RECT 1169.630 1309.870 1170.175 1310.185 ;
        RECT 1169.845 1309.855 1170.175 1309.870 ;
        RECT 1169.845 1263.250 1170.175 1263.265 ;
        RECT 1170.510 1263.250 1170.890 1263.260 ;
        RECT 1169.845 1262.950 1170.890 1263.250 ;
        RECT 1169.845 1262.935 1170.175 1262.950 ;
        RECT 1170.510 1262.940 1170.890 1262.950 ;
        RECT 1170.510 1238.770 1170.890 1238.780 ;
        RECT 1172.350 1238.770 1172.730 1238.780 ;
        RECT 1170.510 1238.470 1172.730 1238.770 ;
        RECT 1170.510 1238.460 1170.890 1238.470 ;
        RECT 1172.350 1238.460 1172.730 1238.470 ;
        RECT 1172.350 1125.890 1172.730 1125.900 ;
        RECT 1171.470 1125.590 1172.730 1125.890 ;
        RECT 1171.470 1124.540 1171.770 1125.590 ;
        RECT 1172.350 1125.580 1172.730 1125.590 ;
        RECT 1171.430 1124.220 1171.810 1124.540 ;
        RECT 1171.685 1034.770 1172.015 1034.785 ;
        RECT 1172.350 1034.770 1172.730 1034.780 ;
        RECT 1171.685 1034.470 1172.730 1034.770 ;
        RECT 1171.685 1034.455 1172.015 1034.470 ;
        RECT 1172.350 1034.460 1172.730 1034.470 ;
        RECT 1171.685 987.850 1172.015 987.865 ;
        RECT 1171.470 987.535 1172.015 987.850 ;
        RECT 1171.470 987.180 1171.770 987.535 ;
        RECT 1171.430 986.860 1171.810 987.180 ;
        RECT 1171.430 938.890 1171.810 938.900 ;
        RECT 1172.350 938.890 1172.730 938.900 ;
        RECT 1171.430 938.590 1172.730 938.890 ;
        RECT 1171.430 938.580 1171.810 938.590 ;
        RECT 1172.350 938.580 1172.730 938.590 ;
        RECT 1172.605 937.540 1172.935 937.545 ;
        RECT 1172.350 937.530 1172.935 937.540 ;
        RECT 1172.150 937.230 1172.935 937.530 ;
        RECT 1172.350 937.220 1172.935 937.230 ;
        RECT 1172.605 937.215 1172.935 937.220 ;
        RECT 1172.605 890.610 1172.935 890.625 ;
        RECT 1173.270 890.610 1173.650 890.620 ;
        RECT 1172.605 890.310 1173.650 890.610 ;
        RECT 1172.605 890.295 1172.935 890.310 ;
        RECT 1173.270 890.300 1173.650 890.310 ;
        RECT 1171.430 821.250 1171.810 821.260 ;
        RECT 1173.270 821.250 1173.650 821.260 ;
        RECT 1171.430 820.950 1173.650 821.250 ;
        RECT 1171.430 820.940 1171.810 820.950 ;
        RECT 1173.270 820.940 1173.650 820.950 ;
        RECT 1171.430 772.970 1171.810 772.980 ;
        RECT 1172.350 772.970 1172.730 772.980 ;
        RECT 1171.430 772.670 1172.730 772.970 ;
        RECT 1171.430 772.660 1171.810 772.670 ;
        RECT 1172.350 772.660 1172.730 772.670 ;
        RECT 1171.430 724.690 1171.810 724.700 ;
        RECT 1172.350 724.690 1172.730 724.700 ;
        RECT 1171.430 724.390 1172.730 724.690 ;
        RECT 1171.430 724.380 1171.810 724.390 ;
        RECT 1172.350 724.380 1172.730 724.390 ;
        RECT 1171.685 693.420 1172.015 693.425 ;
        RECT 1171.430 693.410 1172.015 693.420 ;
        RECT 1171.230 693.110 1172.015 693.410 ;
        RECT 1171.430 693.100 1172.015 693.110 ;
        RECT 1171.685 693.095 1172.015 693.100 ;
        RECT 1171.685 609.090 1172.015 609.105 ;
        RECT 1171.685 608.790 1172.690 609.090 ;
        RECT 1171.685 608.775 1172.015 608.790 ;
        RECT 1172.390 608.420 1172.690 608.790 ;
        RECT 1172.350 608.100 1172.730 608.420 ;
        RECT 1173.525 607.060 1173.855 607.065 ;
        RECT 1173.270 607.050 1173.855 607.060 ;
        RECT 1173.070 606.750 1173.855 607.050 ;
        RECT 1173.270 606.740 1173.855 606.750 ;
        RECT 1173.525 606.735 1173.855 606.740 ;
        RECT 1173.525 564.900 1173.855 564.905 ;
        RECT 1173.270 564.890 1173.855 564.900 ;
        RECT 1173.270 564.590 1174.080 564.890 ;
        RECT 1173.270 564.580 1173.855 564.590 ;
        RECT 1173.525 564.575 1173.855 564.580 ;
        RECT 1171.430 483.290 1171.810 483.300 ;
        RECT 1172.350 483.290 1172.730 483.300 ;
        RECT 1171.430 482.990 1172.730 483.290 ;
        RECT 1171.430 482.980 1171.810 482.990 ;
        RECT 1172.350 482.980 1172.730 482.990 ;
        RECT 1172.350 449.290 1172.730 449.300 ;
        RECT 1171.470 448.990 1172.730 449.290 ;
        RECT 1171.470 447.940 1171.770 448.990 ;
        RECT 1172.350 448.980 1172.730 448.990 ;
        RECT 1171.430 447.620 1171.810 447.940 ;
        RECT 1171.430 403.730 1171.810 403.740 ;
        RECT 1173.270 403.730 1173.650 403.740 ;
        RECT 1171.430 403.430 1173.650 403.730 ;
        RECT 1171.430 403.420 1171.810 403.430 ;
        RECT 1173.270 403.420 1173.650 403.430 ;
        RECT 1172.350 379.250 1172.730 379.260 ;
        RECT 1173.270 379.250 1173.650 379.260 ;
        RECT 1172.350 378.950 1173.650 379.250 ;
        RECT 1172.350 378.940 1172.730 378.950 ;
        RECT 1173.270 378.940 1173.650 378.950 ;
        RECT 1170.510 219.450 1170.890 219.460 ;
        RECT 1200.205 219.450 1200.535 219.465 ;
        RECT 1170.510 219.150 1200.535 219.450 ;
        RECT 1170.510 219.140 1170.890 219.150 ;
        RECT 1200.205 219.135 1200.535 219.150 ;
        RECT 2917.600 205.170 2924.800 205.620 ;
        RECT 2916.710 204.870 2924.800 205.170 ;
        RECT 1290.110 202.450 1290.490 202.460 ;
        RECT 1272.670 202.150 1290.490 202.450 ;
        RECT 1200.205 201.090 1200.535 201.105 ;
        RECT 1272.670 201.090 1272.970 202.150 ;
        RECT 1290.110 202.140 1290.490 202.150 ;
        RECT 1748.985 202.450 1749.315 202.465 ;
        RECT 2062.245 202.450 2062.575 202.465 ;
        RECT 2069.605 202.450 2069.935 202.465 ;
        RECT 2656.310 202.450 2656.690 202.460 ;
        RECT 2704.405 202.450 2704.735 202.465 ;
        RECT 1748.985 202.150 1798.290 202.450 ;
        RECT 1748.985 202.135 1749.315 202.150 ;
        RECT 1338.665 201.770 1338.995 201.785 ;
        RECT 1200.205 200.790 1272.970 201.090 ;
        RECT 1337.990 201.470 1338.995 201.770 ;
        RECT 1200.205 200.775 1200.535 200.790 ;
        RECT 1290.110 200.410 1290.490 200.420 ;
        RECT 1337.990 200.410 1338.290 201.470 ;
        RECT 1338.665 201.455 1338.995 201.470 ;
        RECT 1386.505 201.770 1386.835 201.785 ;
        RECT 1393.405 201.770 1393.735 201.785 ;
        RECT 1386.505 201.470 1393.735 201.770 ;
        RECT 1386.505 201.455 1386.835 201.470 ;
        RECT 1393.405 201.455 1393.735 201.470 ;
        RECT 1465.870 201.470 1514.930 201.770 ;
        RECT 1290.110 200.110 1338.290 200.410 ;
        RECT 1393.405 200.410 1393.735 200.425 ;
        RECT 1465.870 200.410 1466.170 201.470 ;
        RECT 1393.405 200.110 1466.170 200.410 ;
        RECT 1514.630 200.410 1514.930 201.470 ;
        RECT 1586.605 201.090 1586.935 201.105 ;
        RECT 1633.985 201.090 1634.315 201.105 ;
        RECT 1586.605 200.790 1634.315 201.090 ;
        RECT 1586.605 200.775 1586.935 200.790 ;
        RECT 1633.985 200.775 1634.315 200.790 ;
        RECT 1705.285 201.090 1705.615 201.105 ;
        RECT 1748.985 201.090 1749.315 201.105 ;
        RECT 1705.285 200.790 1749.315 201.090 ;
        RECT 1705.285 200.775 1705.615 200.790 ;
        RECT 1748.985 200.775 1749.315 200.790 ;
        RECT 1559.005 200.410 1559.335 200.425 ;
        RECT 1514.630 200.110 1559.335 200.410 ;
        RECT 1290.110 200.100 1290.490 200.110 ;
        RECT 1393.405 200.095 1393.735 200.110 ;
        RECT 1559.005 200.095 1559.335 200.110 ;
        RECT 1634.905 200.410 1635.235 200.425 ;
        RECT 1676.510 200.410 1676.890 200.420 ;
        RECT 1634.905 200.110 1676.890 200.410 ;
        RECT 1797.990 200.410 1798.290 202.150 ;
        RECT 2062.245 202.150 2069.935 202.450 ;
        RECT 2062.245 202.135 2062.575 202.150 ;
        RECT 2069.605 202.135 2069.935 202.150 ;
        RECT 2463.150 202.150 2511.290 202.450 ;
        RECT 1918.470 201.770 1918.850 201.780 ;
        RECT 2014.865 201.770 2015.195 201.785 ;
        RECT 1918.470 201.470 2015.195 201.770 ;
        RECT 1918.470 201.460 1918.850 201.470 ;
        RECT 2014.865 201.455 2015.195 201.470 ;
        RECT 2124.590 201.470 2138.690 201.770 ;
        RECT 1917.805 201.090 1918.135 201.105 ;
        RECT 2069.605 201.090 2069.935 201.105 ;
        RECT 2124.590 201.090 2124.890 201.470 ;
        RECT 1917.805 200.790 1918.810 201.090 ;
        RECT 1917.805 200.775 1918.135 200.790 ;
        RECT 1917.805 200.410 1918.135 200.425 ;
        RECT 1918.510 200.420 1918.810 200.790 ;
        RECT 2069.605 200.790 2124.890 201.090 ;
        RECT 2069.605 200.775 2069.935 200.790 ;
        RECT 1797.990 200.110 1822.210 200.410 ;
        RECT 1634.905 200.095 1635.235 200.110 ;
        RECT 1676.510 200.100 1676.890 200.110 ;
        RECT 1821.910 199.730 1822.210 200.110 ;
        RECT 1869.750 200.110 1918.135 200.410 ;
        RECT 1869.750 199.730 1870.050 200.110 ;
        RECT 1917.805 200.095 1918.135 200.110 ;
        RECT 1918.470 200.100 1918.850 200.420 ;
        RECT 2138.390 200.410 2138.690 201.470 ;
        RECT 2139.310 201.470 2187.450 201.770 ;
        RECT 2139.310 200.410 2139.610 201.470 ;
        RECT 2138.390 200.110 2139.610 200.410 ;
        RECT 2187.150 200.410 2187.450 201.470 ;
        RECT 2283.505 201.090 2283.835 201.105 ;
        RECT 2235.910 200.790 2283.835 201.090 ;
        RECT 2235.910 200.410 2236.210 200.790 ;
        RECT 2283.505 200.775 2283.835 200.790 ;
        RECT 2284.425 201.090 2284.755 201.105 ;
        RECT 2463.150 201.090 2463.450 202.150 ;
        RECT 2510.990 201.780 2511.290 202.150 ;
        RECT 2656.310 202.150 2704.735 202.450 ;
        RECT 2656.310 202.140 2656.690 202.150 ;
        RECT 2704.405 202.135 2704.735 202.150 ;
        RECT 2510.950 201.460 2511.330 201.780 ;
        RECT 2801.005 201.770 2801.335 201.785 ;
        RECT 2801.005 201.470 2815.810 201.770 ;
        RECT 2801.005 201.455 2801.335 201.470 ;
        RECT 2572.845 201.090 2573.175 201.105 ;
        RECT 2284.425 200.790 2331.890 201.090 ;
        RECT 2284.425 200.775 2284.755 200.790 ;
        RECT 2187.150 200.110 2236.210 200.410 ;
        RECT 2331.590 200.410 2331.890 200.790 ;
        RECT 2332.510 200.790 2414.690 201.090 ;
        RECT 2332.510 200.410 2332.810 200.790 ;
        RECT 2331.590 200.110 2332.810 200.410 ;
        RECT 2414.390 200.410 2414.690 200.790 ;
        RECT 2429.110 200.790 2463.450 201.090 ;
        RECT 2525.710 200.790 2573.175 201.090 ;
        RECT 2429.110 200.410 2429.410 200.790 ;
        RECT 2414.390 200.110 2429.410 200.410 ;
        RECT 2510.950 200.410 2511.330 200.420 ;
        RECT 2525.710 200.410 2526.010 200.790 ;
        RECT 2572.845 200.775 2573.175 200.790 ;
        RECT 2632.185 201.090 2632.515 201.105 ;
        RECT 2656.310 201.090 2656.690 201.100 ;
        RECT 2752.910 201.090 2753.290 201.100 ;
        RECT 2632.185 200.790 2656.690 201.090 ;
        RECT 2632.185 200.775 2632.515 200.790 ;
        RECT 2656.310 200.780 2656.690 200.790 ;
        RECT 2718.910 200.790 2753.290 201.090 ;
        RECT 2608.265 200.410 2608.595 200.425 ;
        RECT 2510.950 200.110 2526.010 200.410 ;
        RECT 2607.590 200.110 2608.595 200.410 ;
        RECT 2510.950 200.100 2511.330 200.110 ;
        RECT 1821.910 199.430 1870.050 199.730 ;
        RECT 1676.510 199.050 1676.890 199.060 ;
        RECT 1705.285 199.050 1705.615 199.065 ;
        RECT 1676.510 198.750 1705.615 199.050 ;
        RECT 1676.510 198.740 1676.890 198.750 ;
        RECT 1705.285 198.735 1705.615 198.750 ;
        RECT 2572.845 199.050 2573.175 199.065 ;
        RECT 2607.590 199.050 2607.890 200.110 ;
        RECT 2608.265 200.095 2608.595 200.110 ;
        RECT 2704.405 200.410 2704.735 200.425 ;
        RECT 2718.910 200.410 2719.210 200.790 ;
        RECT 2752.910 200.780 2753.290 200.790 ;
        RECT 2704.405 200.110 2719.210 200.410 ;
        RECT 2815.510 200.410 2815.810 201.470 ;
        RECT 2863.105 201.090 2863.435 201.105 ;
        RECT 2916.710 201.090 2917.010 204.870 ;
        RECT 2917.600 204.420 2924.800 204.870 ;
        RECT 2849.550 200.790 2863.435 201.090 ;
        RECT 2849.550 200.410 2849.850 200.790 ;
        RECT 2863.105 200.775 2863.435 200.790 ;
        RECT 2884.510 200.790 2917.010 201.090 ;
        RECT 2815.510 200.110 2849.850 200.410 ;
        RECT 2863.565 200.410 2863.895 200.425 ;
        RECT 2884.510 200.410 2884.810 200.790 ;
        RECT 2863.565 200.110 2884.810 200.410 ;
        RECT 2704.405 200.095 2704.735 200.110 ;
        RECT 2863.565 200.095 2863.895 200.110 ;
        RECT 2752.910 199.730 2753.290 199.740 ;
        RECT 2801.005 199.730 2801.335 199.745 ;
        RECT 2752.910 199.430 2801.335 199.730 ;
        RECT 2752.910 199.420 2753.290 199.430 ;
        RECT 2801.005 199.415 2801.335 199.430 ;
        RECT 2572.845 198.750 2607.890 199.050 ;
        RECT 2572.845 198.735 2573.175 198.750 ;
      LAYER via3 ;
        RECT 1172.380 3196.180 1172.700 3196.500 ;
        RECT 1171.460 1683.180 1171.780 1683.500 ;
        RECT 1173.300 1635.580 1173.620 1635.900 ;
        RECT 1173.300 1594.780 1173.620 1595.100 ;
        RECT 1171.460 1594.100 1171.780 1594.420 ;
        RECT 1171.460 1515.220 1171.780 1515.540 ;
        RECT 1171.460 1497.540 1171.780 1497.860 ;
        RECT 1171.460 1451.980 1171.780 1452.300 ;
        RECT 1173.300 1451.980 1173.620 1452.300 ;
        RECT 1172.380 1366.980 1172.700 1367.300 ;
        RECT 1170.540 1366.300 1170.860 1366.620 ;
        RECT 1170.540 1318.700 1170.860 1319.020 ;
        RECT 1169.620 1317.340 1169.940 1317.660 ;
        RECT 1169.620 1310.540 1169.940 1310.860 ;
        RECT 1170.540 1262.940 1170.860 1263.260 ;
        RECT 1170.540 1238.460 1170.860 1238.780 ;
        RECT 1172.380 1238.460 1172.700 1238.780 ;
        RECT 1172.380 1125.580 1172.700 1125.900 ;
        RECT 1171.460 1124.220 1171.780 1124.540 ;
        RECT 1172.380 1034.460 1172.700 1034.780 ;
        RECT 1171.460 986.860 1171.780 987.180 ;
        RECT 1171.460 938.580 1171.780 938.900 ;
        RECT 1172.380 938.580 1172.700 938.900 ;
        RECT 1172.380 937.220 1172.700 937.540 ;
        RECT 1173.300 890.300 1173.620 890.620 ;
        RECT 1171.460 820.940 1171.780 821.260 ;
        RECT 1173.300 820.940 1173.620 821.260 ;
        RECT 1171.460 772.660 1171.780 772.980 ;
        RECT 1172.380 772.660 1172.700 772.980 ;
        RECT 1171.460 724.380 1171.780 724.700 ;
        RECT 1172.380 724.380 1172.700 724.700 ;
        RECT 1171.460 693.100 1171.780 693.420 ;
        RECT 1172.380 608.100 1172.700 608.420 ;
        RECT 1173.300 606.740 1173.620 607.060 ;
        RECT 1173.300 564.580 1173.620 564.900 ;
        RECT 1171.460 482.980 1171.780 483.300 ;
        RECT 1172.380 482.980 1172.700 483.300 ;
        RECT 1172.380 448.980 1172.700 449.300 ;
        RECT 1171.460 447.620 1171.780 447.940 ;
        RECT 1171.460 403.420 1171.780 403.740 ;
        RECT 1173.300 403.420 1173.620 403.740 ;
        RECT 1172.380 378.940 1172.700 379.260 ;
        RECT 1173.300 378.940 1173.620 379.260 ;
        RECT 1170.540 219.140 1170.860 219.460 ;
        RECT 1290.140 202.140 1290.460 202.460 ;
        RECT 1290.140 200.100 1290.460 200.420 ;
        RECT 1676.540 200.100 1676.860 200.420 ;
        RECT 1918.500 201.460 1918.820 201.780 ;
        RECT 1918.500 200.100 1918.820 200.420 ;
        RECT 2656.340 202.140 2656.660 202.460 ;
        RECT 2510.980 201.460 2511.300 201.780 ;
        RECT 2510.980 200.100 2511.300 200.420 ;
        RECT 2656.340 200.780 2656.660 201.100 ;
        RECT 1676.540 198.740 1676.860 199.060 ;
        RECT 2752.940 200.780 2753.260 201.100 ;
        RECT 2752.940 199.420 2753.260 199.740 ;
      LAYER met4 ;
        RECT 1172.375 3196.175 1172.705 3196.505 ;
        RECT 1172.390 2647.490 1172.690 3196.175 ;
        RECT 1171.950 2646.310 1173.130 2647.490 ;
        RECT 1177.470 2646.310 1178.650 2647.490 ;
        RECT 1177.910 2603.290 1178.210 2646.310 ;
        RECT 1171.950 2602.110 1173.130 2603.290 ;
        RECT 1177.470 2602.110 1178.650 2603.290 ;
        RECT 1172.390 2453.690 1172.690 2602.110 ;
        RECT 1167.350 2452.510 1168.530 2453.690 ;
        RECT 1171.950 2452.510 1173.130 2453.690 ;
        RECT 1167.790 2409.490 1168.090 2452.510 ;
        RECT 1167.350 2408.310 1168.530 2409.490 ;
        RECT 1171.950 2408.310 1173.130 2409.490 ;
        RECT 1172.390 1970.890 1172.690 2408.310 ;
        RECT 1171.950 1969.710 1173.130 1970.890 ;
        RECT 1177.470 1969.710 1178.650 1970.890 ;
        RECT 1177.910 1926.690 1178.210 1969.710 ;
        RECT 1171.950 1925.510 1173.130 1926.690 ;
        RECT 1177.470 1925.510 1178.650 1926.690 ;
        RECT 1172.390 1780.490 1172.690 1925.510 ;
        RECT 1167.350 1779.310 1168.530 1780.490 ;
        RECT 1171.950 1779.310 1173.130 1780.490 ;
        RECT 1167.790 1732.890 1168.090 1779.310 ;
        RECT 1167.350 1731.710 1168.530 1732.890 ;
        RECT 1171.950 1731.710 1173.130 1732.890 ;
        RECT 1172.390 1708.650 1172.690 1731.710 ;
        RECT 1170.550 1708.350 1172.690 1708.650 ;
        RECT 1170.550 1701.850 1170.850 1708.350 ;
        RECT 1170.550 1701.550 1171.770 1701.850 ;
        RECT 1171.470 1683.505 1171.770 1701.550 ;
        RECT 1171.455 1683.175 1171.785 1683.505 ;
        RECT 1173.295 1635.575 1173.625 1635.905 ;
        RECT 1173.310 1595.105 1173.610 1635.575 ;
        RECT 1173.295 1594.775 1173.625 1595.105 ;
        RECT 1171.455 1594.095 1171.785 1594.425 ;
        RECT 1171.470 1515.545 1171.770 1594.095 ;
        RECT 1171.455 1515.215 1171.785 1515.545 ;
        RECT 1171.455 1497.535 1171.785 1497.865 ;
        RECT 1171.470 1452.305 1171.770 1497.535 ;
        RECT 1171.455 1451.975 1171.785 1452.305 ;
        RECT 1173.295 1451.975 1173.625 1452.305 ;
        RECT 1173.310 1395.850 1173.610 1451.975 ;
        RECT 1172.390 1395.550 1173.610 1395.850 ;
        RECT 1172.390 1367.305 1172.690 1395.550 ;
        RECT 1172.375 1366.975 1172.705 1367.305 ;
        RECT 1170.535 1366.295 1170.865 1366.625 ;
        RECT 1170.550 1319.025 1170.850 1366.295 ;
        RECT 1170.535 1318.695 1170.865 1319.025 ;
        RECT 1169.615 1317.335 1169.945 1317.665 ;
        RECT 1169.630 1310.865 1169.930 1317.335 ;
        RECT 1169.615 1310.535 1169.945 1310.865 ;
        RECT 1170.535 1262.935 1170.865 1263.265 ;
        RECT 1170.550 1238.785 1170.850 1262.935 ;
        RECT 1170.535 1238.455 1170.865 1238.785 ;
        RECT 1172.375 1238.455 1172.705 1238.785 ;
        RECT 1172.390 1125.905 1172.690 1238.455 ;
        RECT 1172.375 1125.575 1172.705 1125.905 ;
        RECT 1171.455 1124.215 1171.785 1124.545 ;
        RECT 1171.470 1079.650 1171.770 1124.215 ;
        RECT 1171.470 1079.350 1172.690 1079.650 ;
        RECT 1172.390 1034.785 1172.690 1079.350 ;
        RECT 1172.375 1034.455 1172.705 1034.785 ;
        RECT 1171.455 986.855 1171.785 987.185 ;
        RECT 1171.470 938.905 1171.770 986.855 ;
        RECT 1171.455 938.575 1171.785 938.905 ;
        RECT 1172.375 938.575 1172.705 938.905 ;
        RECT 1172.390 937.545 1172.690 938.575 ;
        RECT 1172.375 937.215 1172.705 937.545 ;
        RECT 1173.295 890.295 1173.625 890.625 ;
        RECT 1173.310 821.265 1173.610 890.295 ;
        RECT 1171.455 820.935 1171.785 821.265 ;
        RECT 1173.295 820.935 1173.625 821.265 ;
        RECT 1171.470 772.985 1171.770 820.935 ;
        RECT 1171.455 772.655 1171.785 772.985 ;
        RECT 1172.375 772.655 1172.705 772.985 ;
        RECT 1172.390 724.705 1172.690 772.655 ;
        RECT 1171.455 724.375 1171.785 724.705 ;
        RECT 1172.375 724.375 1172.705 724.705 ;
        RECT 1171.470 693.425 1171.770 724.375 ;
        RECT 1171.455 693.095 1171.785 693.425 ;
        RECT 1172.375 608.095 1172.705 608.425 ;
        RECT 1172.390 607.050 1172.690 608.095 ;
        RECT 1173.295 607.050 1173.625 607.065 ;
        RECT 1172.390 606.750 1173.625 607.050 ;
        RECT 1173.295 606.735 1173.625 606.750 ;
        RECT 1173.295 564.575 1173.625 564.905 ;
        RECT 1173.310 542.450 1173.610 564.575 ;
        RECT 1171.470 542.150 1173.610 542.450 ;
        RECT 1171.470 483.305 1171.770 542.150 ;
        RECT 1171.455 482.975 1171.785 483.305 ;
        RECT 1172.375 482.975 1172.705 483.305 ;
        RECT 1172.390 449.305 1172.690 482.975 ;
        RECT 1172.375 448.975 1172.705 449.305 ;
        RECT 1171.455 447.615 1171.785 447.945 ;
        RECT 1171.470 403.745 1171.770 447.615 ;
        RECT 1171.455 403.415 1171.785 403.745 ;
        RECT 1173.295 403.415 1173.625 403.745 ;
        RECT 1173.310 379.265 1173.610 403.415 ;
        RECT 1172.375 378.935 1172.705 379.265 ;
        RECT 1173.295 378.935 1173.625 379.265 ;
        RECT 1172.390 256.850 1172.690 378.935 ;
        RECT 1170.550 256.550 1172.690 256.850 ;
        RECT 1170.550 219.465 1170.850 256.550 ;
        RECT 1170.535 219.135 1170.865 219.465 ;
        RECT 1290.135 202.135 1290.465 202.465 ;
        RECT 2656.335 202.135 2656.665 202.465 ;
        RECT 1290.150 200.425 1290.450 202.135 ;
        RECT 1918.495 201.455 1918.825 201.785 ;
        RECT 2510.975 201.455 2511.305 201.785 ;
        RECT 1918.510 200.425 1918.810 201.455 ;
        RECT 2510.990 200.425 2511.290 201.455 ;
        RECT 2656.350 201.105 2656.650 202.135 ;
        RECT 2656.335 200.775 2656.665 201.105 ;
        RECT 2752.935 200.775 2753.265 201.105 ;
        RECT 1290.135 200.095 1290.465 200.425 ;
        RECT 1676.535 200.095 1676.865 200.425 ;
        RECT 1918.495 200.095 1918.825 200.425 ;
        RECT 2510.975 200.095 2511.305 200.425 ;
        RECT 1676.550 199.065 1676.850 200.095 ;
        RECT 2752.950 199.745 2753.250 200.775 ;
        RECT 2752.935 199.415 2753.265 199.745 ;
        RECT 1676.535 198.735 1676.865 199.065 ;
      LAYER met5 ;
        RECT 1171.740 2646.100 1178.860 2647.700 ;
        RECT 1171.740 2601.900 1178.860 2603.500 ;
        RECT 1167.140 2452.300 1173.340 2453.900 ;
        RECT 1167.140 2408.100 1173.340 2409.700 ;
        RECT 1171.740 1969.500 1178.860 1971.100 ;
        RECT 1171.740 1925.300 1178.860 1926.900 ;
        RECT 1167.140 1779.100 1173.340 1780.700 ;
        RECT 1167.140 1731.500 1173.340 1733.100 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1562.690 3205.420 1563.010 3205.480 ;
        RECT 2655.650 3205.420 2655.970 3205.480 ;
        RECT 1562.690 3205.280 2655.970 3205.420 ;
        RECT 1562.690 3205.220 1563.010 3205.280 ;
        RECT 2655.650 3205.220 2655.970 3205.280 ;
        RECT 2655.650 2552.960 2655.970 2553.020 ;
        RECT 2900.370 2552.960 2900.690 2553.020 ;
        RECT 2655.650 2552.820 2900.690 2552.960 ;
        RECT 2655.650 2552.760 2655.970 2552.820 ;
        RECT 2900.370 2552.760 2900.690 2552.820 ;
      LAYER via ;
        RECT 1562.720 3205.220 1562.980 3205.480 ;
        RECT 2655.680 3205.220 2655.940 3205.480 ;
        RECT 2655.680 2552.760 2655.940 2553.020 ;
        RECT 2900.400 2552.760 2900.660 2553.020 ;
      LAYER met2 ;
        RECT 1562.720 3205.190 1562.980 3205.510 ;
        RECT 2655.680 3205.190 2655.940 3205.510 ;
        RECT 1562.780 3200.000 1562.920 3205.190 ;
        RECT 1562.640 3196.000 1562.920 3200.000 ;
        RECT 2655.740 2553.050 2655.880 3205.190 ;
        RECT 2655.680 2552.730 2655.940 2553.050 ;
        RECT 2900.400 2552.730 2900.660 2553.050 ;
        RECT 2900.460 2551.885 2900.600 2552.730 ;
        RECT 2900.390 2551.515 2900.670 2551.885 ;
      LAYER via2 ;
        RECT 2900.390 2551.560 2900.670 2551.840 ;
      LAYER met3 ;
        RECT 2900.365 2551.850 2900.695 2551.865 ;
        RECT 2917.600 2551.850 2924.800 2552.300 ;
        RECT 2900.365 2551.550 2924.800 2551.850 ;
        RECT 2900.365 2551.535 2900.695 2551.550 ;
        RECT 2917.600 2551.100 2924.800 2551.550 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1602.250 3205.760 1602.570 3205.820 ;
        RECT 2652.430 3205.760 2652.750 3205.820 ;
        RECT 1602.250 3205.620 2652.750 3205.760 ;
        RECT 1602.250 3205.560 1602.570 3205.620 ;
        RECT 2652.430 3205.560 2652.750 3205.620 ;
        RECT 2652.430 2787.560 2652.750 2787.620 ;
        RECT 2900.370 2787.560 2900.690 2787.620 ;
        RECT 2652.430 2787.420 2900.690 2787.560 ;
        RECT 2652.430 2787.360 2652.750 2787.420 ;
        RECT 2900.370 2787.360 2900.690 2787.420 ;
      LAYER via ;
        RECT 1602.280 3205.560 1602.540 3205.820 ;
        RECT 2652.460 3205.560 2652.720 3205.820 ;
        RECT 2652.460 2787.360 2652.720 2787.620 ;
        RECT 2900.400 2787.360 2900.660 2787.620 ;
      LAYER met2 ;
        RECT 1602.280 3205.530 1602.540 3205.850 ;
        RECT 2652.460 3205.530 2652.720 3205.850 ;
        RECT 1602.340 3200.000 1602.480 3205.530 ;
        RECT 1602.200 3196.000 1602.480 3200.000 ;
        RECT 2652.520 2787.650 2652.660 3205.530 ;
        RECT 2652.460 2787.330 2652.720 2787.650 ;
        RECT 2900.400 2787.330 2900.660 2787.650 ;
        RECT 2900.460 2786.485 2900.600 2787.330 ;
        RECT 2900.390 2786.115 2900.670 2786.485 ;
      LAYER via2 ;
        RECT 2900.390 2786.160 2900.670 2786.440 ;
      LAYER met3 ;
        RECT 2900.365 2786.450 2900.695 2786.465 ;
        RECT 2917.600 2786.450 2924.800 2786.900 ;
        RECT 2900.365 2786.150 2924.800 2786.450 ;
        RECT 2900.365 2786.135 2900.695 2786.150 ;
        RECT 2917.600 2785.700 2924.800 2786.150 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1642.270 3198.620 1642.590 3198.680 ;
        RECT 1690.110 3198.620 1690.430 3198.680 ;
        RECT 1642.270 3198.480 1690.430 3198.620 ;
        RECT 1642.270 3198.420 1642.590 3198.480 ;
        RECT 1690.110 3198.420 1690.430 3198.480 ;
        RECT 2651.510 3022.160 2651.830 3022.220 ;
        RECT 2900.370 3022.160 2900.690 3022.220 ;
        RECT 2651.510 3022.020 2900.690 3022.160 ;
        RECT 2651.510 3021.960 2651.830 3022.020 ;
        RECT 2900.370 3021.960 2900.690 3022.020 ;
      LAYER via ;
        RECT 1642.300 3198.420 1642.560 3198.680 ;
        RECT 1690.140 3198.420 1690.400 3198.680 ;
        RECT 2651.540 3021.960 2651.800 3022.220 ;
        RECT 2900.400 3021.960 2900.660 3022.220 ;
      LAYER met2 ;
        RECT 1641.760 3197.090 1642.040 3200.000 ;
        RECT 1642.300 3198.390 1642.560 3198.710 ;
        RECT 1690.140 3198.390 1690.400 3198.710 ;
        RECT 1642.360 3197.090 1642.500 3198.390 ;
        RECT 1641.760 3196.950 1642.500 3197.090 ;
        RECT 1641.760 3196.000 1642.040 3196.950 ;
        RECT 1690.200 3196.525 1690.340 3198.390 ;
        RECT 1990.510 3198.195 1990.790 3198.565 ;
        RECT 1990.580 3197.205 1990.720 3198.195 ;
        RECT 1990.510 3196.835 1990.790 3197.205 ;
        RECT 1690.130 3196.155 1690.410 3196.525 ;
        RECT 2651.530 3194.115 2651.810 3194.485 ;
        RECT 2651.600 3022.250 2651.740 3194.115 ;
        RECT 2651.540 3021.930 2651.800 3022.250 ;
        RECT 2900.400 3021.930 2900.660 3022.250 ;
        RECT 2900.460 3021.085 2900.600 3021.930 ;
        RECT 2900.390 3020.715 2900.670 3021.085 ;
      LAYER via2 ;
        RECT 1990.510 3198.240 1990.790 3198.520 ;
        RECT 1990.510 3196.880 1990.790 3197.160 ;
        RECT 1690.130 3196.200 1690.410 3196.480 ;
        RECT 2651.530 3194.160 2651.810 3194.440 ;
        RECT 2900.390 3020.760 2900.670 3021.040 ;
      LAYER met3 ;
        RECT 1990.485 3198.530 1990.815 3198.545 ;
        RECT 2014.150 3198.530 2014.530 3198.540 ;
        RECT 1990.485 3198.230 2014.530 3198.530 ;
        RECT 1990.485 3198.215 1990.815 3198.230 ;
        RECT 2014.150 3198.220 2014.530 3198.230 ;
        RECT 1924.910 3197.170 1925.290 3197.180 ;
        RECT 1990.485 3197.170 1990.815 3197.185 ;
        RECT 1924.910 3196.870 1990.815 3197.170 ;
        RECT 1924.910 3196.860 1925.290 3196.870 ;
        RECT 1990.485 3196.855 1990.815 3196.870 ;
        RECT 1690.105 3196.490 1690.435 3196.505 ;
        RECT 1713.310 3196.490 1713.690 3196.500 ;
        RECT 1690.105 3196.190 1713.690 3196.490 ;
        RECT 1690.105 3196.175 1690.435 3196.190 ;
        RECT 1713.310 3196.180 1713.690 3196.190 ;
        RECT 2014.150 3195.130 2014.530 3195.140 ;
        RECT 1812.710 3194.830 1824.970 3195.130 ;
        RECT 1713.310 3194.450 1713.690 3194.460 ;
        RECT 1812.710 3194.450 1813.010 3194.830 ;
        RECT 1713.310 3194.150 1813.010 3194.450 ;
        RECT 1824.670 3194.450 1824.970 3194.830 ;
        RECT 2014.150 3194.830 2015.410 3195.130 ;
        RECT 2014.150 3194.820 2014.530 3194.830 ;
        RECT 1922.150 3194.450 1922.530 3194.460 ;
        RECT 1824.670 3194.150 1922.530 3194.450 ;
        RECT 1713.310 3194.140 1713.690 3194.150 ;
        RECT 1922.150 3194.140 1922.530 3194.150 ;
        RECT 1923.990 3194.450 1924.370 3194.460 ;
        RECT 1924.910 3194.450 1925.290 3194.460 ;
        RECT 1923.990 3194.150 1925.290 3194.450 ;
        RECT 2015.110 3194.450 2015.410 3194.830 ;
        RECT 2041.750 3194.450 2042.130 3194.460 ;
        RECT 2015.110 3194.150 2042.130 3194.450 ;
        RECT 1923.990 3194.140 1924.370 3194.150 ;
        RECT 1924.910 3194.140 1925.290 3194.150 ;
        RECT 2041.750 3194.140 2042.130 3194.150 ;
        RECT 2042.670 3194.450 2043.050 3194.460 ;
        RECT 2187.110 3194.450 2187.490 3194.460 ;
        RECT 2042.670 3194.150 2044.850 3194.450 ;
        RECT 2042.670 3194.140 2043.050 3194.150 ;
        RECT 2044.550 3193.770 2044.850 3194.150 ;
        RECT 2109.870 3194.150 2187.490 3194.450 ;
        RECT 2109.870 3193.770 2110.170 3194.150 ;
        RECT 2187.110 3194.140 2187.490 3194.150 ;
        RECT 2188.950 3194.450 2189.330 3194.460 ;
        RECT 2651.505 3194.450 2651.835 3194.465 ;
        RECT 2188.950 3194.150 2651.835 3194.450 ;
        RECT 2188.950 3194.140 2189.330 3194.150 ;
        RECT 2651.505 3194.135 2651.835 3194.150 ;
        RECT 2044.550 3193.470 2110.170 3193.770 ;
        RECT 2900.365 3021.050 2900.695 3021.065 ;
        RECT 2917.600 3021.050 2924.800 3021.500 ;
        RECT 2900.365 3020.750 2924.800 3021.050 ;
        RECT 2900.365 3020.735 2900.695 3020.750 ;
        RECT 2917.600 3020.300 2924.800 3020.750 ;
      LAYER via3 ;
        RECT 2014.180 3198.220 2014.500 3198.540 ;
        RECT 1924.940 3196.860 1925.260 3197.180 ;
        RECT 1713.340 3196.180 1713.660 3196.500 ;
        RECT 1713.340 3194.140 1713.660 3194.460 ;
        RECT 2014.180 3194.820 2014.500 3195.140 ;
        RECT 1922.180 3194.140 1922.500 3194.460 ;
        RECT 1924.020 3194.140 1924.340 3194.460 ;
        RECT 1924.940 3194.140 1925.260 3194.460 ;
        RECT 2041.780 3194.140 2042.100 3194.460 ;
        RECT 2042.700 3194.140 2043.020 3194.460 ;
        RECT 2187.140 3194.140 2187.460 3194.460 ;
        RECT 2188.980 3194.140 2189.300 3194.460 ;
      LAYER met4 ;
        RECT 2014.175 3198.215 2014.505 3198.545 ;
        RECT 1924.935 3196.855 1925.265 3197.185 ;
        RECT 1713.335 3196.175 1713.665 3196.505 ;
        RECT 1713.350 3194.465 1713.650 3196.175 ;
        RECT 1924.950 3194.465 1925.250 3196.855 ;
        RECT 2014.190 3195.145 2014.490 3198.215 ;
        RECT 2014.175 3194.815 2014.505 3195.145 ;
        RECT 1713.335 3194.135 1713.665 3194.465 ;
        RECT 1922.175 3194.450 1922.505 3194.465 ;
        RECT 1924.015 3194.450 1924.345 3194.465 ;
        RECT 1922.175 3194.150 1924.345 3194.450 ;
        RECT 1922.175 3194.135 1922.505 3194.150 ;
        RECT 1924.015 3194.135 1924.345 3194.150 ;
        RECT 1924.935 3194.135 1925.265 3194.465 ;
        RECT 2041.775 3194.450 2042.105 3194.465 ;
        RECT 2042.695 3194.450 2043.025 3194.465 ;
        RECT 2041.775 3194.150 2043.025 3194.450 ;
        RECT 2041.775 3194.135 2042.105 3194.150 ;
        RECT 2042.695 3194.135 2043.025 3194.150 ;
        RECT 2187.135 3194.450 2187.465 3194.465 ;
        RECT 2188.975 3194.450 2189.305 3194.465 ;
        RECT 2187.135 3194.150 2189.305 3194.450 ;
        RECT 2187.135 3194.135 2187.465 3194.150 ;
        RECT 2188.975 3194.135 2189.305 3194.150 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1683.210 3250.300 1683.530 3250.360 ;
        RECT 2900.830 3250.300 2901.150 3250.360 ;
        RECT 1683.210 3250.160 2901.150 3250.300 ;
        RECT 1683.210 3250.100 1683.530 3250.160 ;
        RECT 2900.830 3250.100 2901.150 3250.160 ;
      LAYER via ;
        RECT 1683.240 3250.100 1683.500 3250.360 ;
        RECT 2900.860 3250.100 2901.120 3250.360 ;
      LAYER met2 ;
        RECT 2900.850 3255.315 2901.130 3255.685 ;
        RECT 2900.920 3250.390 2901.060 3255.315 ;
        RECT 1683.240 3250.070 1683.500 3250.390 ;
        RECT 2900.860 3250.070 2901.120 3250.390 ;
        RECT 1681.320 3199.810 1681.600 3200.000 ;
        RECT 1683.300 3199.810 1683.440 3250.070 ;
        RECT 1681.320 3199.670 1683.440 3199.810 ;
        RECT 1681.320 3196.000 1681.600 3199.670 ;
      LAYER via2 ;
        RECT 2900.850 3255.360 2901.130 3255.640 ;
      LAYER met3 ;
        RECT 2900.825 3255.650 2901.155 3255.665 ;
        RECT 2917.600 3255.650 2924.800 3256.100 ;
        RECT 2900.825 3255.350 2924.800 3255.650 ;
        RECT 2900.825 3255.335 2901.155 3255.350 ;
        RECT 2917.600 3254.900 2924.800 3255.350 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1724.610 3484.900 1724.930 3484.960 ;
        RECT 2900.830 3484.900 2901.150 3484.960 ;
        RECT 1724.610 3484.760 2901.150 3484.900 ;
        RECT 1724.610 3484.700 1724.930 3484.760 ;
        RECT 2900.830 3484.700 2901.150 3484.760 ;
      LAYER via ;
        RECT 1724.640 3484.700 1724.900 3484.960 ;
        RECT 2900.860 3484.700 2901.120 3484.960 ;
      LAYER met2 ;
        RECT 2900.850 3489.915 2901.130 3490.285 ;
        RECT 2900.920 3484.990 2901.060 3489.915 ;
        RECT 1724.640 3484.670 1724.900 3484.990 ;
        RECT 2900.860 3484.670 2901.120 3484.990 ;
        RECT 1724.700 3200.490 1724.840 3484.670 ;
        RECT 1722.860 3200.350 1724.840 3200.490 ;
        RECT 1720.880 3199.810 1721.160 3200.000 ;
        RECT 1722.860 3199.810 1723.000 3200.350 ;
        RECT 1720.880 3199.670 1723.000 3199.810 ;
        RECT 1720.880 3196.000 1721.160 3199.670 ;
      LAYER via2 ;
        RECT 2900.850 3489.960 2901.130 3490.240 ;
      LAYER met3 ;
        RECT 2900.825 3490.250 2901.155 3490.265 ;
        RECT 2917.600 3490.250 2924.800 3490.700 ;
        RECT 2900.825 3489.950 2924.800 3490.250 ;
        RECT 2900.825 3489.935 2901.155 3489.950 ;
        RECT 2917.600 3489.500 2924.800 3489.950 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1766.010 3501.220 1766.330 3501.280 ;
        RECT 2635.870 3501.220 2636.190 3501.280 ;
        RECT 1766.010 3501.080 2636.190 3501.220 ;
        RECT 1766.010 3501.020 1766.330 3501.080 ;
        RECT 2635.870 3501.020 2636.190 3501.080 ;
      LAYER via ;
        RECT 1766.040 3501.020 1766.300 3501.280 ;
        RECT 2635.900 3501.020 2636.160 3501.280 ;
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
        RECT 2635.960 3501.310 2636.100 3517.600 ;
        RECT 1766.040 3500.990 1766.300 3501.310 ;
        RECT 2635.900 3500.990 2636.160 3501.310 ;
        RECT 1766.100 3200.490 1766.240 3500.990 ;
        RECT 1762.880 3200.350 1766.240 3200.490 ;
        RECT 1759.980 3199.810 1760.260 3200.000 ;
        RECT 1762.880 3199.810 1763.020 3200.350 ;
        RECT 1759.980 3199.670 1763.020 3199.810 ;
        RECT 1759.980 3196.000 1760.260 3199.670 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1800.510 3500.200 1800.830 3500.260 ;
        RECT 2311.570 3500.200 2311.890 3500.260 ;
        RECT 1800.510 3500.060 2311.890 3500.200 ;
        RECT 1800.510 3500.000 1800.830 3500.060 ;
        RECT 2311.570 3500.000 2311.890 3500.060 ;
      LAYER via ;
        RECT 1800.540 3500.000 1800.800 3500.260 ;
        RECT 2311.600 3500.000 2311.860 3500.260 ;
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
        RECT 2311.660 3500.290 2311.800 3517.600 ;
        RECT 1800.540 3499.970 1800.800 3500.290 ;
        RECT 2311.600 3499.970 2311.860 3500.290 ;
        RECT 1799.540 3199.810 1799.820 3200.000 ;
        RECT 1800.600 3199.810 1800.740 3499.970 ;
        RECT 1799.540 3199.670 1800.740 3199.810 ;
        RECT 1799.540 3196.000 1799.820 3199.670 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1841.910 3498.500 1842.230 3498.560 ;
        RECT 1987.270 3498.500 1987.590 3498.560 ;
        RECT 1841.910 3498.360 1987.590 3498.500 ;
        RECT 1841.910 3498.300 1842.230 3498.360 ;
        RECT 1987.270 3498.300 1987.590 3498.360 ;
      LAYER via ;
        RECT 1841.940 3498.300 1842.200 3498.560 ;
        RECT 1987.300 3498.300 1987.560 3498.560 ;
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
        RECT 1987.360 3498.590 1987.500 3517.600 ;
        RECT 1841.940 3498.270 1842.200 3498.590 ;
        RECT 1987.300 3498.270 1987.560 3498.590 ;
        RECT 1839.100 3199.130 1839.380 3200.000 ;
        RECT 1842.000 3199.130 1842.140 3498.270 ;
        RECT 1839.100 3198.990 1842.140 3199.130 ;
        RECT 1839.100 3196.000 1839.380 3198.990 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1662.510 3499.520 1662.830 3499.580 ;
        RECT 1876.870 3499.520 1877.190 3499.580 ;
        RECT 1662.510 3499.380 1877.190 3499.520 ;
        RECT 1662.510 3499.320 1662.830 3499.380 ;
        RECT 1876.870 3499.320 1877.190 3499.380 ;
      LAYER via ;
        RECT 1662.540 3499.320 1662.800 3499.580 ;
        RECT 1876.900 3499.320 1877.160 3499.580 ;
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
        RECT 1662.600 3499.610 1662.740 3517.600 ;
        RECT 1662.540 3499.290 1662.800 3499.610 ;
        RECT 1876.900 3499.290 1877.160 3499.610 ;
        RECT 1876.960 3199.810 1877.100 3499.290 ;
        RECT 1878.660 3199.810 1878.940 3200.000 ;
        RECT 1876.960 3199.670 1878.940 3199.810 ;
        RECT 1878.660 3196.000 1878.940 3199.670 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1338.210 3500.880 1338.530 3500.940 ;
        RECT 1918.270 3500.880 1918.590 3500.940 ;
        RECT 1338.210 3500.740 1918.590 3500.880 ;
        RECT 1338.210 3500.680 1338.530 3500.740 ;
        RECT 1918.270 3500.680 1918.590 3500.740 ;
      LAYER via ;
        RECT 1338.240 3500.680 1338.500 3500.940 ;
        RECT 1918.300 3500.680 1918.560 3500.940 ;
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
        RECT 1338.300 3500.970 1338.440 3517.600 ;
        RECT 1338.240 3500.650 1338.500 3500.970 ;
        RECT 1918.300 3500.650 1918.560 3500.970 ;
        RECT 1918.360 3200.000 1918.500 3500.650 ;
        RECT 1918.220 3196.000 1918.500 3200.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1828.110 436.120 1828.430 436.180 ;
        RECT 1869.510 436.120 1869.830 436.180 ;
        RECT 1828.110 435.980 1869.830 436.120 ;
        RECT 1828.110 435.920 1828.430 435.980 ;
        RECT 1869.510 435.920 1869.830 435.980 ;
        RECT 1338.670 435.780 1338.990 435.840 ;
        RECT 1368.570 435.780 1368.890 435.840 ;
        RECT 1338.670 435.640 1368.890 435.780 ;
        RECT 1338.670 435.580 1338.990 435.640 ;
        RECT 1368.570 435.580 1368.890 435.640 ;
        RECT 1642.730 435.780 1643.050 435.840 ;
        RECT 1690.110 435.780 1690.430 435.840 ;
        RECT 1642.730 435.640 1690.430 435.780 ;
        RECT 1642.730 435.580 1643.050 435.640 ;
        RECT 1690.110 435.580 1690.430 435.640 ;
        RECT 1703.910 435.780 1704.230 435.840 ;
        RECT 1772.910 435.780 1773.230 435.840 ;
        RECT 1703.910 435.640 1773.230 435.780 ;
        RECT 1703.910 435.580 1704.230 435.640 ;
        RECT 1772.910 435.580 1773.230 435.640 ;
        RECT 2076.970 435.440 2077.290 435.500 ;
        RECT 2123.890 435.440 2124.210 435.500 ;
        RECT 2076.970 435.300 2124.210 435.440 ;
        RECT 2076.970 435.240 2077.290 435.300 ;
        RECT 2123.890 435.240 2124.210 435.300 ;
        RECT 2379.650 435.440 2379.970 435.500 ;
        RECT 2380.570 435.440 2380.890 435.500 ;
        RECT 2379.650 435.300 2380.890 435.440 ;
        RECT 2379.650 435.240 2379.970 435.300 ;
        RECT 2380.570 435.240 2380.890 435.300 ;
        RECT 2863.110 435.440 2863.430 435.500 ;
        RECT 2883.810 435.440 2884.130 435.500 ;
        RECT 2863.110 435.300 2884.130 435.440 ;
        RECT 2863.110 435.240 2863.430 435.300 ;
        RECT 2883.810 435.240 2884.130 435.300 ;
        RECT 2125.270 435.100 2125.590 435.160 ;
        RECT 2172.650 435.100 2172.970 435.160 ;
        RECT 2125.270 434.960 2172.970 435.100 ;
        RECT 2125.270 434.900 2125.590 434.960 ;
        RECT 2172.650 434.900 2172.970 434.960 ;
      LAYER via ;
        RECT 1828.140 435.920 1828.400 436.180 ;
        RECT 1869.540 435.920 1869.800 436.180 ;
        RECT 1338.700 435.580 1338.960 435.840 ;
        RECT 1368.600 435.580 1368.860 435.840 ;
        RECT 1642.760 435.580 1643.020 435.840 ;
        RECT 1690.140 435.580 1690.400 435.840 ;
        RECT 1703.940 435.580 1704.200 435.840 ;
        RECT 1772.940 435.580 1773.200 435.840 ;
        RECT 2077.000 435.240 2077.260 435.500 ;
        RECT 2123.920 435.240 2124.180 435.500 ;
        RECT 2379.680 435.240 2379.940 435.500 ;
        RECT 2380.600 435.240 2380.860 435.500 ;
        RECT 2863.140 435.240 2863.400 435.500 ;
        RECT 2883.840 435.240 2884.100 435.500 ;
        RECT 2125.300 434.900 2125.560 435.160 ;
        RECT 2172.680 434.900 2172.940 435.160 ;
      LAYER met2 ;
        RECT 1207.520 3196.410 1207.800 3200.000 ;
        RECT 1209.430 3196.410 1209.710 3196.525 ;
        RECT 1207.520 3196.270 1209.710 3196.410 ;
        RECT 1207.520 3196.000 1207.800 3196.270 ;
        RECT 1209.430 3196.155 1209.710 3196.270 ;
        RECT 2801.030 437.395 2801.310 437.765 ;
        RECT 1607.330 436.715 1607.610 437.085 ;
        RECT 2680.510 436.715 2680.790 437.085 ;
        RECT 1338.700 435.725 1338.960 435.870 ;
        RECT 1368.600 435.725 1368.860 435.870 ;
        RECT 1607.400 435.725 1607.540 436.715 ;
        RECT 1690.130 436.035 1690.410 436.405 ;
        RECT 1703.930 436.035 1704.210 436.405 ;
        RECT 1772.930 436.035 1773.210 436.405 ;
        RECT 1828.130 436.035 1828.410 436.405 ;
        RECT 1690.200 435.870 1690.340 436.035 ;
        RECT 1704.000 435.870 1704.140 436.035 ;
        RECT 1773.000 435.870 1773.140 436.035 ;
        RECT 1828.140 435.890 1828.400 436.035 ;
        RECT 1869.540 435.890 1869.800 436.210 ;
        RECT 1924.730 436.035 1925.010 436.405 ;
        RECT 2172.670 436.035 2172.950 436.405 ;
        RECT 1642.760 435.725 1643.020 435.870 ;
        RECT 1296.830 435.355 1297.110 435.725 ;
        RECT 1338.690 435.355 1338.970 435.725 ;
        RECT 1368.590 435.355 1368.870 435.725 ;
        RECT 1607.330 435.355 1607.610 435.725 ;
        RECT 1642.750 435.355 1643.030 435.725 ;
        RECT 1690.140 435.550 1690.400 435.870 ;
        RECT 1703.940 435.550 1704.200 435.870 ;
        RECT 1772.940 435.550 1773.200 435.870 ;
        RECT 1869.600 435.725 1869.740 435.890 ;
        RECT 1869.530 435.355 1869.810 435.725 ;
        RECT 1289.930 434.675 1290.210 435.045 ;
        RECT 1290.000 434.365 1290.140 434.675 ;
        RECT 1296.900 434.365 1297.040 435.355 ;
        RECT 1924.800 434.365 1924.940 436.035 ;
        RECT 2076.990 435.355 2077.270 435.725 ;
        RECT 2077.000 435.210 2077.260 435.355 ;
        RECT 2123.920 435.210 2124.180 435.530 ;
        RECT 2123.980 434.930 2124.120 435.210 ;
        RECT 2172.740 435.190 2172.880 436.035 ;
        RECT 2379.670 435.355 2379.950 435.725 ;
        RECT 2380.590 435.355 2380.870 435.725 ;
        RECT 2379.680 435.210 2379.940 435.355 ;
        RECT 2380.600 435.210 2380.860 435.355 ;
        RECT 2125.300 435.045 2125.560 435.190 ;
        RECT 2124.370 434.930 2124.650 435.045 ;
        RECT 2123.980 434.790 2124.650 434.930 ;
        RECT 2124.370 434.675 2124.650 434.790 ;
        RECT 2125.290 434.675 2125.570 435.045 ;
        RECT 2172.680 434.870 2172.940 435.190 ;
        RECT 2680.580 435.045 2680.720 436.715 ;
        RECT 2801.100 436.405 2801.240 437.395 ;
        RECT 2801.030 436.035 2801.310 436.405 ;
        RECT 2863.130 435.355 2863.410 435.725 ;
        RECT 2883.830 435.355 2884.110 435.725 ;
        RECT 2863.140 435.210 2863.400 435.355 ;
        RECT 2883.840 435.210 2884.100 435.355 ;
        RECT 2625.310 434.675 2625.590 435.045 ;
        RECT 2680.510 434.675 2680.790 435.045 ;
        RECT 1289.930 433.995 1290.210 434.365 ;
        RECT 1296.830 433.995 1297.110 434.365 ;
        RECT 1924.730 433.995 1925.010 434.365 ;
        RECT 2625.380 433.685 2625.520 434.675 ;
        RECT 2625.310 433.315 2625.590 433.685 ;
      LAYER via2 ;
        RECT 1209.430 3196.200 1209.710 3196.480 ;
        RECT 2801.030 437.440 2801.310 437.720 ;
        RECT 1607.330 436.760 1607.610 437.040 ;
        RECT 2680.510 436.760 2680.790 437.040 ;
        RECT 1690.130 436.080 1690.410 436.360 ;
        RECT 1703.930 436.080 1704.210 436.360 ;
        RECT 1772.930 436.080 1773.210 436.360 ;
        RECT 1828.130 436.080 1828.410 436.360 ;
        RECT 1924.730 436.080 1925.010 436.360 ;
        RECT 2172.670 436.080 2172.950 436.360 ;
        RECT 1296.830 435.400 1297.110 435.680 ;
        RECT 1338.690 435.400 1338.970 435.680 ;
        RECT 1368.590 435.400 1368.870 435.680 ;
        RECT 1607.330 435.400 1607.610 435.680 ;
        RECT 1642.750 435.400 1643.030 435.680 ;
        RECT 1869.530 435.400 1869.810 435.680 ;
        RECT 1289.930 434.720 1290.210 435.000 ;
        RECT 2076.990 435.400 2077.270 435.680 ;
        RECT 2379.670 435.400 2379.950 435.680 ;
        RECT 2380.590 435.400 2380.870 435.680 ;
        RECT 2124.370 434.720 2124.650 435.000 ;
        RECT 2125.290 434.720 2125.570 435.000 ;
        RECT 2801.030 436.080 2801.310 436.360 ;
        RECT 2863.130 435.400 2863.410 435.680 ;
        RECT 2883.830 435.400 2884.110 435.680 ;
        RECT 2625.310 434.720 2625.590 435.000 ;
        RECT 2680.510 434.720 2680.790 435.000 ;
        RECT 1289.930 434.040 1290.210 434.320 ;
        RECT 1296.830 434.040 1297.110 434.320 ;
        RECT 1924.730 434.040 1925.010 434.320 ;
        RECT 2625.310 433.360 2625.590 433.640 ;
      LAYER met3 ;
        RECT 1209.405 3196.490 1209.735 3196.505 ;
        RECT 1213.750 3196.490 1214.130 3196.500 ;
        RECT 1209.405 3196.190 1214.130 3196.490 ;
        RECT 1209.405 3196.175 1209.735 3196.190 ;
        RECT 1213.750 3196.180 1214.130 3196.190 ;
        RECT 2917.600 439.770 2924.800 440.220 ;
        RECT 2916.710 439.470 2924.800 439.770 ;
        RECT 2752.910 437.730 2753.290 437.740 ;
        RECT 2801.005 437.730 2801.335 437.745 ;
        RECT 2752.910 437.430 2801.335 437.730 ;
        RECT 2752.910 437.420 2753.290 437.430 ;
        RECT 2801.005 437.415 2801.335 437.430 ;
        RECT 1497.110 437.050 1497.490 437.060 ;
        RECT 1461.270 436.750 1497.490 437.050 ;
        RECT 1213.750 435.690 1214.130 435.700 ;
        RECT 1296.805 435.690 1297.135 435.705 ;
        RECT 1338.665 435.690 1338.995 435.705 ;
        RECT 1213.750 435.390 1242.610 435.690 ;
        RECT 1213.750 435.380 1214.130 435.390 ;
        RECT 1242.310 435.010 1242.610 435.390 ;
        RECT 1296.805 435.390 1338.995 435.690 ;
        RECT 1296.805 435.375 1297.135 435.390 ;
        RECT 1338.665 435.375 1338.995 435.390 ;
        RECT 1368.565 435.690 1368.895 435.705 ;
        RECT 1461.270 435.690 1461.570 436.750 ;
        RECT 1497.110 436.740 1497.490 436.750 ;
        RECT 1587.270 437.050 1587.650 437.060 ;
        RECT 1607.305 437.050 1607.635 437.065 ;
        RECT 2680.485 437.050 2680.815 437.065 ;
        RECT 1587.270 436.750 1607.635 437.050 ;
        RECT 1587.270 436.740 1587.650 436.750 ;
        RECT 1607.305 436.735 1607.635 436.750 ;
        RECT 2282.830 436.750 2318.090 437.050 ;
        RECT 1690.105 436.370 1690.435 436.385 ;
        RECT 1703.905 436.370 1704.235 436.385 ;
        RECT 1690.105 436.070 1704.235 436.370 ;
        RECT 1690.105 436.055 1690.435 436.070 ;
        RECT 1703.905 436.055 1704.235 436.070 ;
        RECT 1772.905 436.370 1773.235 436.385 ;
        RECT 1828.105 436.370 1828.435 436.385 ;
        RECT 1924.705 436.380 1925.035 436.385 ;
        RECT 1924.705 436.370 1925.290 436.380 ;
        RECT 1772.905 436.070 1828.435 436.370 ;
        RECT 1924.500 436.070 1925.290 436.370 ;
        RECT 1772.905 436.055 1773.235 436.070 ;
        RECT 1828.105 436.055 1828.435 436.070 ;
        RECT 1924.705 436.060 1925.290 436.070 ;
        RECT 1925.830 436.370 1926.210 436.380 ;
        RECT 2172.645 436.370 2172.975 436.385 ;
        RECT 1925.830 436.070 1994.250 436.370 ;
        RECT 1925.830 436.060 1926.210 436.070 ;
        RECT 1924.705 436.055 1925.035 436.060 ;
        RECT 1368.565 435.390 1461.570 435.690 ;
        RECT 1497.110 435.690 1497.490 435.700 ;
        RECT 1587.270 435.690 1587.650 435.700 ;
        RECT 1497.110 435.390 1587.650 435.690 ;
        RECT 1368.565 435.375 1368.895 435.390 ;
        RECT 1497.110 435.380 1497.490 435.390 ;
        RECT 1587.270 435.380 1587.650 435.390 ;
        RECT 1607.305 435.690 1607.635 435.705 ;
        RECT 1642.725 435.690 1643.055 435.705 ;
        RECT 1607.305 435.390 1643.055 435.690 ;
        RECT 1607.305 435.375 1607.635 435.390 ;
        RECT 1642.725 435.375 1643.055 435.390 ;
        RECT 1869.505 435.690 1869.835 435.705 ;
        RECT 1877.070 435.690 1877.450 435.700 ;
        RECT 1869.505 435.390 1877.450 435.690 ;
        RECT 1869.505 435.375 1869.835 435.390 ;
        RECT 1877.070 435.380 1877.450 435.390 ;
        RECT 1289.905 435.010 1290.235 435.025 ;
        RECT 1242.310 434.710 1290.235 435.010 ;
        RECT 1993.950 435.010 1994.250 436.070 ;
        RECT 2172.645 436.070 2187.450 436.370 ;
        RECT 2172.645 436.055 2172.975 436.070 ;
        RECT 2076.965 435.690 2077.295 435.705 ;
        RECT 2042.710 435.390 2077.295 435.690 ;
        RECT 2042.710 435.010 2043.010 435.390 ;
        RECT 2076.965 435.375 2077.295 435.390 ;
        RECT 1993.950 434.710 2043.010 435.010 ;
        RECT 2124.345 435.010 2124.675 435.025 ;
        RECT 2125.265 435.010 2125.595 435.025 ;
        RECT 2124.345 434.710 2125.595 435.010 ;
        RECT 2187.150 435.010 2187.450 436.070 ;
        RECT 2282.830 435.690 2283.130 436.750 ;
        RECT 2317.790 436.380 2318.090 436.750 ;
        RECT 2463.150 436.750 2511.290 437.050 ;
        RECT 2317.750 436.060 2318.130 436.380 ;
        RECT 2379.645 435.690 2379.975 435.705 ;
        RECT 2235.910 435.390 2283.130 435.690 ;
        RECT 2332.510 435.390 2379.975 435.690 ;
        RECT 2235.910 435.010 2236.210 435.390 ;
        RECT 2187.150 434.710 2236.210 435.010 ;
        RECT 2317.750 435.010 2318.130 435.020 ;
        RECT 2332.510 435.010 2332.810 435.390 ;
        RECT 2379.645 435.375 2379.975 435.390 ;
        RECT 2380.565 435.690 2380.895 435.705 ;
        RECT 2463.150 435.690 2463.450 436.750 ;
        RECT 2510.990 436.380 2511.290 436.750 ;
        RECT 2656.350 436.750 2680.815 437.050 ;
        RECT 2510.950 436.060 2511.330 436.380 ;
        RECT 2656.350 435.690 2656.650 436.750 ;
        RECT 2680.485 436.735 2680.815 436.750 ;
        RECT 2801.005 436.370 2801.335 436.385 ;
        RECT 2801.005 436.070 2815.810 436.370 ;
        RECT 2801.005 436.055 2801.335 436.070 ;
        RECT 2752.910 435.690 2753.290 435.700 ;
        RECT 2380.565 435.390 2414.690 435.690 ;
        RECT 2380.565 435.375 2380.895 435.390 ;
        RECT 2317.750 434.710 2332.810 435.010 ;
        RECT 2414.390 435.010 2414.690 435.390 ;
        RECT 2429.110 435.390 2463.450 435.690 ;
        RECT 2525.710 435.390 2583.970 435.690 ;
        RECT 2429.110 435.010 2429.410 435.390 ;
        RECT 2414.390 434.710 2429.410 435.010 ;
        RECT 2510.950 435.010 2511.330 435.020 ;
        RECT 2525.710 435.010 2526.010 435.390 ;
        RECT 2510.950 434.710 2526.010 435.010 ;
        RECT 2583.670 435.010 2583.970 435.390 ;
        RECT 2648.990 435.390 2656.650 435.690 ;
        RECT 2718.910 435.390 2753.290 435.690 ;
        RECT 2601.110 435.010 2601.490 435.020 ;
        RECT 2583.670 434.710 2601.490 435.010 ;
        RECT 1289.905 434.695 1290.235 434.710 ;
        RECT 2124.345 434.695 2124.675 434.710 ;
        RECT 2125.265 434.695 2125.595 434.710 ;
        RECT 2317.750 434.700 2318.130 434.710 ;
        RECT 2510.950 434.700 2511.330 434.710 ;
        RECT 2601.110 434.700 2601.490 434.710 ;
        RECT 2625.285 435.010 2625.615 435.025 ;
        RECT 2648.990 435.010 2649.290 435.390 ;
        RECT 2625.285 434.710 2649.290 435.010 ;
        RECT 2680.485 435.010 2680.815 435.025 ;
        RECT 2718.910 435.010 2719.210 435.390 ;
        RECT 2752.910 435.380 2753.290 435.390 ;
        RECT 2680.485 434.710 2719.210 435.010 ;
        RECT 2815.510 435.010 2815.810 436.070 ;
        RECT 2863.105 435.690 2863.435 435.705 ;
        RECT 2849.550 435.390 2863.435 435.690 ;
        RECT 2849.550 435.010 2849.850 435.390 ;
        RECT 2863.105 435.375 2863.435 435.390 ;
        RECT 2883.805 435.690 2884.135 435.705 ;
        RECT 2916.710 435.690 2917.010 439.470 ;
        RECT 2917.600 439.020 2924.800 439.470 ;
        RECT 2883.805 435.390 2917.010 435.690 ;
        RECT 2883.805 435.375 2884.135 435.390 ;
        RECT 2815.510 434.710 2849.850 435.010 ;
        RECT 2625.285 434.695 2625.615 434.710 ;
        RECT 2680.485 434.695 2680.815 434.710 ;
        RECT 1289.905 434.330 1290.235 434.345 ;
        RECT 1296.805 434.330 1297.135 434.345 ;
        RECT 1289.905 434.030 1297.135 434.330 ;
        RECT 1289.905 434.015 1290.235 434.030 ;
        RECT 1296.805 434.015 1297.135 434.030 ;
        RECT 1877.070 434.330 1877.450 434.340 ;
        RECT 1924.705 434.330 1925.035 434.345 ;
        RECT 1877.070 434.030 1925.035 434.330 ;
        RECT 1877.070 434.020 1877.450 434.030 ;
        RECT 1924.705 434.015 1925.035 434.030 ;
        RECT 2601.110 433.650 2601.490 433.660 ;
        RECT 2625.285 433.650 2625.615 433.665 ;
        RECT 2601.110 433.350 2625.615 433.650 ;
        RECT 2601.110 433.340 2601.490 433.350 ;
        RECT 2625.285 433.335 2625.615 433.350 ;
      LAYER via3 ;
        RECT 1213.780 3196.180 1214.100 3196.500 ;
        RECT 2752.940 437.420 2753.260 437.740 ;
        RECT 1213.780 435.380 1214.100 435.700 ;
        RECT 1497.140 436.740 1497.460 437.060 ;
        RECT 1587.300 436.740 1587.620 437.060 ;
        RECT 1924.940 436.060 1925.260 436.380 ;
        RECT 1925.860 436.060 1926.180 436.380 ;
        RECT 1497.140 435.380 1497.460 435.700 ;
        RECT 1587.300 435.380 1587.620 435.700 ;
        RECT 1877.100 435.380 1877.420 435.700 ;
        RECT 2317.780 436.060 2318.100 436.380 ;
        RECT 2317.780 434.700 2318.100 435.020 ;
        RECT 2510.980 436.060 2511.300 436.380 ;
        RECT 2510.980 434.700 2511.300 435.020 ;
        RECT 2601.140 434.700 2601.460 435.020 ;
        RECT 2752.940 435.380 2753.260 435.700 ;
        RECT 1877.100 434.020 1877.420 434.340 ;
        RECT 2601.140 433.340 2601.460 433.660 ;
      LAYER met4 ;
        RECT 1213.775 3196.175 1214.105 3196.505 ;
        RECT 1213.790 435.705 1214.090 3196.175 ;
        RECT 2752.935 437.415 2753.265 437.745 ;
        RECT 1497.135 436.735 1497.465 437.065 ;
        RECT 1587.295 436.735 1587.625 437.065 ;
        RECT 1924.950 436.750 1926.170 437.050 ;
        RECT 1497.150 435.705 1497.450 436.735 ;
        RECT 1587.310 435.705 1587.610 436.735 ;
        RECT 1924.950 436.385 1925.250 436.750 ;
        RECT 1925.870 436.385 1926.170 436.750 ;
        RECT 1924.935 436.055 1925.265 436.385 ;
        RECT 1925.855 436.055 1926.185 436.385 ;
        RECT 2317.775 436.055 2318.105 436.385 ;
        RECT 2510.975 436.055 2511.305 436.385 ;
        RECT 1213.775 435.375 1214.105 435.705 ;
        RECT 1497.135 435.375 1497.465 435.705 ;
        RECT 1587.295 435.375 1587.625 435.705 ;
        RECT 1877.095 435.375 1877.425 435.705 ;
        RECT 1877.110 434.345 1877.410 435.375 ;
        RECT 2317.790 435.025 2318.090 436.055 ;
        RECT 2510.990 435.025 2511.290 436.055 ;
        RECT 2752.950 435.705 2753.250 437.415 ;
        RECT 2752.935 435.375 2753.265 435.705 ;
        RECT 2317.775 434.695 2318.105 435.025 ;
        RECT 2510.975 434.695 2511.305 435.025 ;
        RECT 2601.135 434.695 2601.465 435.025 ;
        RECT 1877.095 434.015 1877.425 434.345 ;
        RECT 2601.150 433.665 2601.450 434.695 ;
        RECT 2601.135 433.335 2601.465 433.665 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1013.910 3504.280 1014.230 3504.340 ;
        RECT 1952.770 3504.280 1953.090 3504.340 ;
        RECT 1013.910 3504.140 1953.090 3504.280 ;
        RECT 1013.910 3504.080 1014.230 3504.140 ;
        RECT 1952.770 3504.080 1953.090 3504.140 ;
      LAYER via ;
        RECT 1013.940 3504.080 1014.200 3504.340 ;
        RECT 1952.800 3504.080 1953.060 3504.340 ;
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
        RECT 1014.000 3504.370 1014.140 3517.600 ;
        RECT 1013.940 3504.050 1014.200 3504.370 ;
        RECT 1952.800 3504.050 1953.060 3504.370 ;
        RECT 1952.860 3199.130 1953.000 3504.050 ;
        RECT 1957.320 3199.130 1957.600 3200.000 ;
        RECT 1952.860 3198.990 1957.600 3199.130 ;
        RECT 1957.320 3196.000 1957.600 3198.990 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 689.150 3503.260 689.470 3503.320 ;
        RECT 1994.170 3503.260 1994.490 3503.320 ;
        RECT 689.150 3503.120 1994.490 3503.260 ;
        RECT 689.150 3503.060 689.470 3503.120 ;
        RECT 1994.170 3503.060 1994.490 3503.120 ;
      LAYER via ;
        RECT 689.180 3503.060 689.440 3503.320 ;
        RECT 1994.200 3503.060 1994.460 3503.320 ;
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
        RECT 689.240 3503.350 689.380 3517.600 ;
        RECT 689.180 3503.030 689.440 3503.350 ;
        RECT 1994.200 3503.030 1994.460 3503.350 ;
        RECT 1994.260 3200.490 1994.400 3503.030 ;
        RECT 1994.260 3200.350 1995.780 3200.490 ;
        RECT 1995.640 3199.810 1995.780 3200.350 ;
        RECT 1996.880 3199.810 1997.160 3200.000 ;
        RECT 1995.640 3199.670 1997.160 3199.810 ;
        RECT 1996.880 3196.000 1997.160 3199.670 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 364.850 3502.240 365.170 3502.300 ;
        RECT 2035.570 3502.240 2035.890 3502.300 ;
        RECT 364.850 3502.100 2035.890 3502.240 ;
        RECT 364.850 3502.040 365.170 3502.100 ;
        RECT 2035.570 3502.040 2035.890 3502.100 ;
      LAYER via ;
        RECT 364.880 3502.040 365.140 3502.300 ;
        RECT 2035.600 3502.040 2035.860 3502.300 ;
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
        RECT 364.940 3502.330 365.080 3517.600 ;
        RECT 364.880 3502.010 365.140 3502.330 ;
        RECT 2035.600 3502.010 2035.860 3502.330 ;
        RECT 2035.660 3199.810 2035.800 3502.010 ;
        RECT 2036.440 3199.810 2036.720 3200.000 ;
        RECT 2035.660 3199.670 2036.720 3199.810 ;
        RECT 2036.440 3196.000 2036.720 3199.670 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
        RECT 40.640 3501.845 40.780 3517.600 ;
        RECT 40.570 3501.475 40.850 3501.845 ;
        RECT 2070.090 3501.475 2070.370 3501.845 ;
        RECT 2070.160 3199.130 2070.300 3501.475 ;
        RECT 2076.000 3199.130 2076.280 3200.000 ;
        RECT 2070.160 3198.990 2076.280 3199.130 ;
        RECT 2076.000 3196.000 2076.280 3198.990 ;
      LAYER via2 ;
        RECT 40.570 3501.520 40.850 3501.800 ;
        RECT 2070.090 3501.520 2070.370 3501.800 ;
      LAYER met3 ;
        RECT 40.545 3501.810 40.875 3501.825 ;
        RECT 2070.065 3501.810 2070.395 3501.825 ;
        RECT 40.545 3501.510 2070.395 3501.810 ;
        RECT 40.545 3501.495 40.875 3501.510 ;
        RECT 2070.065 3501.495 2070.395 3501.510 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.250 3263.900 15.570 3263.960 ;
        RECT 2111.470 3263.900 2111.790 3263.960 ;
        RECT 15.250 3263.760 2111.790 3263.900 ;
        RECT 15.250 3263.700 15.570 3263.760 ;
        RECT 2111.470 3263.700 2111.790 3263.760 ;
      LAYER via ;
        RECT 15.280 3263.700 15.540 3263.960 ;
        RECT 2111.500 3263.700 2111.760 3263.960 ;
      LAYER met2 ;
        RECT 15.270 3267.555 15.550 3267.925 ;
        RECT 15.340 3263.990 15.480 3267.555 ;
        RECT 15.280 3263.670 15.540 3263.990 ;
        RECT 2111.500 3263.670 2111.760 3263.990 ;
        RECT 2111.560 3199.130 2111.700 3263.670 ;
        RECT 2115.560 3199.130 2115.840 3200.000 ;
        RECT 2111.560 3198.990 2115.840 3199.130 ;
        RECT 2115.560 3196.000 2115.840 3198.990 ;
      LAYER via2 ;
        RECT 15.270 3267.600 15.550 3267.880 ;
      LAYER met3 ;
        RECT -4.800 3267.890 2.400 3268.340 ;
        RECT 15.245 3267.890 15.575 3267.905 ;
        RECT -4.800 3267.590 15.575 3267.890 ;
        RECT -4.800 3267.140 2.400 3267.590 ;
        RECT 15.245 3267.575 15.575 3267.590 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 2980.340 16.030 2980.400 ;
        RECT 40.550 2980.340 40.870 2980.400 ;
        RECT 15.710 2980.200 40.870 2980.340 ;
        RECT 15.710 2980.140 16.030 2980.200 ;
        RECT 40.550 2980.140 40.870 2980.200 ;
      LAYER via ;
        RECT 15.740 2980.140 16.000 2980.400 ;
        RECT 40.580 2980.140 40.840 2980.400 ;
      LAYER met2 ;
        RECT 2100.910 3198.195 2101.190 3198.565 ;
        RECT 2100.980 3196.525 2101.120 3198.195 ;
        RECT 2100.910 3196.155 2101.190 3196.525 ;
        RECT 2153.810 3196.410 2154.090 3196.525 ;
        RECT 2155.120 3196.410 2155.400 3200.000 ;
        RECT 2153.810 3196.270 2155.400 3196.410 ;
        RECT 2153.810 3196.155 2154.090 3196.270 ;
        RECT 2155.120 3196.000 2155.400 3196.270 ;
        RECT 40.570 3194.115 40.850 3194.485 ;
        RECT 87.030 3194.115 87.310 3194.485 ;
        RECT 130.730 3194.115 131.010 3194.485 ;
        RECT 183.630 3194.115 183.910 3194.485 ;
        RECT 227.330 3194.115 227.610 3194.485 ;
        RECT 280.230 3194.115 280.510 3194.485 ;
        RECT 323.930 3194.115 324.210 3194.485 ;
        RECT 376.830 3194.115 377.110 3194.485 ;
        RECT 420.530 3194.115 420.810 3194.485 ;
        RECT 473.430 3194.115 473.710 3194.485 ;
        RECT 517.130 3194.115 517.410 3194.485 ;
        RECT 570.030 3194.115 570.310 3194.485 ;
        RECT 613.730 3194.115 614.010 3194.485 ;
        RECT 666.630 3194.115 666.910 3194.485 ;
        RECT 710.330 3194.115 710.610 3194.485 ;
        RECT 763.230 3194.115 763.510 3194.485 ;
        RECT 806.930 3194.115 807.210 3194.485 ;
        RECT 859.830 3194.115 860.110 3194.485 ;
        RECT 903.530 3194.115 903.810 3194.485 ;
        RECT 956.430 3194.115 956.710 3194.485 ;
        RECT 1000.130 3194.115 1000.410 3194.485 ;
        RECT 1053.030 3194.115 1053.310 3194.485 ;
        RECT 1099.950 3194.115 1100.230 3194.485 ;
        RECT 40.640 2980.430 40.780 3194.115 ;
        RECT 87.100 3190.405 87.240 3194.115 ;
        RECT 130.800 3190.405 130.940 3194.115 ;
        RECT 183.700 3190.405 183.840 3194.115 ;
        RECT 227.400 3190.405 227.540 3194.115 ;
        RECT 280.300 3190.405 280.440 3194.115 ;
        RECT 324.000 3190.405 324.140 3194.115 ;
        RECT 376.900 3190.405 377.040 3194.115 ;
        RECT 420.600 3190.405 420.740 3194.115 ;
        RECT 473.500 3190.405 473.640 3194.115 ;
        RECT 517.200 3190.405 517.340 3194.115 ;
        RECT 570.100 3190.405 570.240 3194.115 ;
        RECT 613.800 3190.405 613.940 3194.115 ;
        RECT 666.700 3190.405 666.840 3194.115 ;
        RECT 710.400 3190.405 710.540 3194.115 ;
        RECT 763.300 3190.405 763.440 3194.115 ;
        RECT 807.000 3190.405 807.140 3194.115 ;
        RECT 859.900 3190.405 860.040 3194.115 ;
        RECT 903.600 3190.405 903.740 3194.115 ;
        RECT 956.500 3190.405 956.640 3194.115 ;
        RECT 1000.200 3190.405 1000.340 3194.115 ;
        RECT 1053.100 3190.405 1053.240 3194.115 ;
        RECT 1100.020 3190.405 1100.160 3194.115 ;
        RECT 87.030 3190.035 87.310 3190.405 ;
        RECT 130.730 3190.035 131.010 3190.405 ;
        RECT 183.630 3190.035 183.910 3190.405 ;
        RECT 227.330 3190.035 227.610 3190.405 ;
        RECT 280.230 3190.035 280.510 3190.405 ;
        RECT 323.930 3190.035 324.210 3190.405 ;
        RECT 376.830 3190.035 377.110 3190.405 ;
        RECT 420.530 3190.035 420.810 3190.405 ;
        RECT 473.430 3190.035 473.710 3190.405 ;
        RECT 517.130 3190.035 517.410 3190.405 ;
        RECT 570.030 3190.035 570.310 3190.405 ;
        RECT 613.730 3190.035 614.010 3190.405 ;
        RECT 666.630 3190.035 666.910 3190.405 ;
        RECT 710.330 3190.035 710.610 3190.405 ;
        RECT 763.230 3190.035 763.510 3190.405 ;
        RECT 806.930 3190.035 807.210 3190.405 ;
        RECT 859.830 3190.035 860.110 3190.405 ;
        RECT 903.530 3190.035 903.810 3190.405 ;
        RECT 956.430 3190.035 956.710 3190.405 ;
        RECT 1000.130 3190.035 1000.410 3190.405 ;
        RECT 1053.030 3190.035 1053.310 3190.405 ;
        RECT 1099.950 3190.035 1100.230 3190.405 ;
        RECT 15.740 2980.285 16.000 2980.430 ;
        RECT 15.730 2979.915 16.010 2980.285 ;
        RECT 40.580 2980.110 40.840 2980.430 ;
      LAYER via2 ;
        RECT 2100.910 3198.240 2101.190 3198.520 ;
        RECT 2100.910 3196.200 2101.190 3196.480 ;
        RECT 2153.810 3196.200 2154.090 3196.480 ;
        RECT 40.570 3194.160 40.850 3194.440 ;
        RECT 87.030 3194.160 87.310 3194.440 ;
        RECT 130.730 3194.160 131.010 3194.440 ;
        RECT 183.630 3194.160 183.910 3194.440 ;
        RECT 227.330 3194.160 227.610 3194.440 ;
        RECT 280.230 3194.160 280.510 3194.440 ;
        RECT 323.930 3194.160 324.210 3194.440 ;
        RECT 376.830 3194.160 377.110 3194.440 ;
        RECT 420.530 3194.160 420.810 3194.440 ;
        RECT 473.430 3194.160 473.710 3194.440 ;
        RECT 517.130 3194.160 517.410 3194.440 ;
        RECT 570.030 3194.160 570.310 3194.440 ;
        RECT 613.730 3194.160 614.010 3194.440 ;
        RECT 666.630 3194.160 666.910 3194.440 ;
        RECT 710.330 3194.160 710.610 3194.440 ;
        RECT 763.230 3194.160 763.510 3194.440 ;
        RECT 806.930 3194.160 807.210 3194.440 ;
        RECT 859.830 3194.160 860.110 3194.440 ;
        RECT 903.530 3194.160 903.810 3194.440 ;
        RECT 956.430 3194.160 956.710 3194.440 ;
        RECT 1000.130 3194.160 1000.410 3194.440 ;
        RECT 1053.030 3194.160 1053.310 3194.440 ;
        RECT 1099.950 3194.160 1100.230 3194.440 ;
        RECT 87.030 3190.080 87.310 3190.360 ;
        RECT 130.730 3190.080 131.010 3190.360 ;
        RECT 183.630 3190.080 183.910 3190.360 ;
        RECT 227.330 3190.080 227.610 3190.360 ;
        RECT 280.230 3190.080 280.510 3190.360 ;
        RECT 323.930 3190.080 324.210 3190.360 ;
        RECT 376.830 3190.080 377.110 3190.360 ;
        RECT 420.530 3190.080 420.810 3190.360 ;
        RECT 473.430 3190.080 473.710 3190.360 ;
        RECT 517.130 3190.080 517.410 3190.360 ;
        RECT 570.030 3190.080 570.310 3190.360 ;
        RECT 613.730 3190.080 614.010 3190.360 ;
        RECT 666.630 3190.080 666.910 3190.360 ;
        RECT 710.330 3190.080 710.610 3190.360 ;
        RECT 763.230 3190.080 763.510 3190.360 ;
        RECT 806.930 3190.080 807.210 3190.360 ;
        RECT 859.830 3190.080 860.110 3190.360 ;
        RECT 903.530 3190.080 903.810 3190.360 ;
        RECT 956.430 3190.080 956.710 3190.360 ;
        RECT 1000.130 3190.080 1000.410 3190.360 ;
        RECT 1053.030 3190.080 1053.310 3190.360 ;
        RECT 1099.950 3190.080 1100.230 3190.360 ;
        RECT 15.730 2979.960 16.010 2980.240 ;
      LAYER met3 ;
        RECT 2100.885 3198.530 2101.215 3198.545 ;
        RECT 2076.750 3198.230 2101.215 3198.530 ;
        RECT 2043.590 3196.490 2043.970 3196.500 ;
        RECT 2076.750 3196.490 2077.050 3198.230 ;
        RECT 2100.885 3198.215 2101.215 3198.230 ;
        RECT 2043.590 3196.190 2077.050 3196.490 ;
        RECT 2100.885 3196.490 2101.215 3196.505 ;
        RECT 2153.785 3196.490 2154.115 3196.505 ;
        RECT 2100.885 3196.190 2154.115 3196.490 ;
        RECT 2043.590 3196.180 2043.970 3196.190 ;
        RECT 2100.885 3196.175 2101.215 3196.190 ;
        RECT 2153.785 3196.175 2154.115 3196.190 ;
        RECT 1288.270 3195.130 1288.650 3195.140 ;
        RECT 1385.790 3195.130 1386.170 3195.140 ;
        RECT 1434.550 3195.130 1434.930 3195.140 ;
        RECT 1775.870 3195.130 1776.250 3195.140 ;
        RECT 1811.750 3195.130 1812.130 3195.140 ;
        RECT 1288.270 3194.830 1290.450 3195.130 ;
        RECT 1288.270 3194.820 1288.650 3194.830 ;
        RECT 40.545 3194.450 40.875 3194.465 ;
        RECT 87.005 3194.450 87.335 3194.465 ;
        RECT 40.545 3194.150 87.335 3194.450 ;
        RECT 40.545 3194.135 40.875 3194.150 ;
        RECT 87.005 3194.135 87.335 3194.150 ;
        RECT 130.705 3194.450 131.035 3194.465 ;
        RECT 183.605 3194.450 183.935 3194.465 ;
        RECT 130.705 3194.150 183.935 3194.450 ;
        RECT 130.705 3194.135 131.035 3194.150 ;
        RECT 183.605 3194.135 183.935 3194.150 ;
        RECT 227.305 3194.450 227.635 3194.465 ;
        RECT 280.205 3194.450 280.535 3194.465 ;
        RECT 227.305 3194.150 280.535 3194.450 ;
        RECT 227.305 3194.135 227.635 3194.150 ;
        RECT 280.205 3194.135 280.535 3194.150 ;
        RECT 323.905 3194.450 324.235 3194.465 ;
        RECT 376.805 3194.450 377.135 3194.465 ;
        RECT 323.905 3194.150 377.135 3194.450 ;
        RECT 323.905 3194.135 324.235 3194.150 ;
        RECT 376.805 3194.135 377.135 3194.150 ;
        RECT 420.505 3194.450 420.835 3194.465 ;
        RECT 473.405 3194.450 473.735 3194.465 ;
        RECT 420.505 3194.150 473.735 3194.450 ;
        RECT 420.505 3194.135 420.835 3194.150 ;
        RECT 473.405 3194.135 473.735 3194.150 ;
        RECT 517.105 3194.450 517.435 3194.465 ;
        RECT 570.005 3194.450 570.335 3194.465 ;
        RECT 517.105 3194.150 570.335 3194.450 ;
        RECT 517.105 3194.135 517.435 3194.150 ;
        RECT 570.005 3194.135 570.335 3194.150 ;
        RECT 613.705 3194.450 614.035 3194.465 ;
        RECT 666.605 3194.450 666.935 3194.465 ;
        RECT 613.705 3194.150 666.935 3194.450 ;
        RECT 613.705 3194.135 614.035 3194.150 ;
        RECT 666.605 3194.135 666.935 3194.150 ;
        RECT 710.305 3194.450 710.635 3194.465 ;
        RECT 763.205 3194.450 763.535 3194.465 ;
        RECT 710.305 3194.150 763.535 3194.450 ;
        RECT 710.305 3194.135 710.635 3194.150 ;
        RECT 763.205 3194.135 763.535 3194.150 ;
        RECT 806.905 3194.450 807.235 3194.465 ;
        RECT 859.805 3194.450 860.135 3194.465 ;
        RECT 806.905 3194.150 860.135 3194.450 ;
        RECT 806.905 3194.135 807.235 3194.150 ;
        RECT 859.805 3194.135 860.135 3194.150 ;
        RECT 903.505 3194.450 903.835 3194.465 ;
        RECT 956.405 3194.450 956.735 3194.465 ;
        RECT 903.505 3194.150 956.735 3194.450 ;
        RECT 903.505 3194.135 903.835 3194.150 ;
        RECT 956.405 3194.135 956.735 3194.150 ;
        RECT 1000.105 3194.450 1000.435 3194.465 ;
        RECT 1053.005 3194.450 1053.335 3194.465 ;
        RECT 1000.105 3194.150 1053.335 3194.450 ;
        RECT 1000.105 3194.135 1000.435 3194.150 ;
        RECT 1053.005 3194.135 1053.335 3194.150 ;
        RECT 1099.925 3194.450 1100.255 3194.465 ;
        RECT 1149.350 3194.450 1149.730 3194.460 ;
        RECT 1099.925 3194.150 1149.730 3194.450 ;
        RECT 1290.150 3194.450 1290.450 3194.830 ;
        RECT 1385.790 3194.830 1387.050 3195.130 ;
        RECT 1385.790 3194.820 1386.170 3194.830 ;
        RECT 1386.750 3194.460 1387.050 3194.830 ;
        RECT 1434.550 3194.830 1580.250 3195.130 ;
        RECT 1434.550 3194.820 1434.930 3194.830 ;
        RECT 1338.870 3194.450 1339.250 3194.460 ;
        RECT 1290.150 3194.150 1339.250 3194.450 ;
        RECT 1099.925 3194.135 1100.255 3194.150 ;
        RECT 1149.350 3194.140 1149.730 3194.150 ;
        RECT 1338.870 3194.140 1339.250 3194.150 ;
        RECT 1386.710 3194.140 1387.090 3194.460 ;
        RECT 1579.950 3194.450 1580.250 3194.830 ;
        RECT 1775.870 3194.830 1812.130 3195.130 ;
        RECT 1775.870 3194.820 1776.250 3194.830 ;
        RECT 1811.750 3194.820 1812.130 3194.830 ;
        RECT 1872.470 3195.130 1872.850 3195.140 ;
        RECT 1872.470 3194.830 1923.410 3195.130 ;
        RECT 1872.470 3194.820 1872.850 3194.830 ;
        RECT 1579.950 3194.150 1680.530 3194.450 ;
        RECT 1680.230 3193.770 1680.530 3194.150 ;
        RECT 1775.870 3193.770 1776.250 3193.780 ;
        RECT 1680.230 3193.470 1776.250 3193.770 ;
        RECT 1775.870 3193.460 1776.250 3193.470 ;
        RECT 1811.750 3193.770 1812.130 3193.780 ;
        RECT 1872.470 3193.770 1872.850 3193.780 ;
        RECT 1811.750 3193.470 1872.850 3193.770 ;
        RECT 1923.110 3193.770 1923.410 3194.830 ;
        RECT 2043.590 3193.770 2043.970 3193.780 ;
        RECT 1923.110 3193.470 2043.970 3193.770 ;
        RECT 1811.750 3193.460 1812.130 3193.470 ;
        RECT 1872.470 3193.460 1872.850 3193.470 ;
        RECT 2043.590 3193.460 2043.970 3193.470 ;
        RECT 87.005 3190.370 87.335 3190.385 ;
        RECT 130.705 3190.370 131.035 3190.385 ;
        RECT 87.005 3190.070 131.035 3190.370 ;
        RECT 87.005 3190.055 87.335 3190.070 ;
        RECT 130.705 3190.055 131.035 3190.070 ;
        RECT 183.605 3190.370 183.935 3190.385 ;
        RECT 227.305 3190.370 227.635 3190.385 ;
        RECT 183.605 3190.070 227.635 3190.370 ;
        RECT 183.605 3190.055 183.935 3190.070 ;
        RECT 227.305 3190.055 227.635 3190.070 ;
        RECT 280.205 3190.370 280.535 3190.385 ;
        RECT 323.905 3190.370 324.235 3190.385 ;
        RECT 280.205 3190.070 324.235 3190.370 ;
        RECT 280.205 3190.055 280.535 3190.070 ;
        RECT 323.905 3190.055 324.235 3190.070 ;
        RECT 376.805 3190.370 377.135 3190.385 ;
        RECT 420.505 3190.370 420.835 3190.385 ;
        RECT 376.805 3190.070 420.835 3190.370 ;
        RECT 376.805 3190.055 377.135 3190.070 ;
        RECT 420.505 3190.055 420.835 3190.070 ;
        RECT 473.405 3190.370 473.735 3190.385 ;
        RECT 517.105 3190.370 517.435 3190.385 ;
        RECT 473.405 3190.070 517.435 3190.370 ;
        RECT 473.405 3190.055 473.735 3190.070 ;
        RECT 517.105 3190.055 517.435 3190.070 ;
        RECT 570.005 3190.370 570.335 3190.385 ;
        RECT 613.705 3190.370 614.035 3190.385 ;
        RECT 570.005 3190.070 614.035 3190.370 ;
        RECT 570.005 3190.055 570.335 3190.070 ;
        RECT 613.705 3190.055 614.035 3190.070 ;
        RECT 666.605 3190.370 666.935 3190.385 ;
        RECT 710.305 3190.370 710.635 3190.385 ;
        RECT 666.605 3190.070 710.635 3190.370 ;
        RECT 666.605 3190.055 666.935 3190.070 ;
        RECT 710.305 3190.055 710.635 3190.070 ;
        RECT 763.205 3190.370 763.535 3190.385 ;
        RECT 806.905 3190.370 807.235 3190.385 ;
        RECT 763.205 3190.070 807.235 3190.370 ;
        RECT 763.205 3190.055 763.535 3190.070 ;
        RECT 806.905 3190.055 807.235 3190.070 ;
        RECT 859.805 3190.370 860.135 3190.385 ;
        RECT 903.505 3190.370 903.835 3190.385 ;
        RECT 859.805 3190.070 903.835 3190.370 ;
        RECT 859.805 3190.055 860.135 3190.070 ;
        RECT 903.505 3190.055 903.835 3190.070 ;
        RECT 956.405 3190.370 956.735 3190.385 ;
        RECT 1000.105 3190.370 1000.435 3190.385 ;
        RECT 956.405 3190.070 1000.435 3190.370 ;
        RECT 956.405 3190.055 956.735 3190.070 ;
        RECT 1000.105 3190.055 1000.435 3190.070 ;
        RECT 1053.005 3190.370 1053.335 3190.385 ;
        RECT 1099.925 3190.370 1100.255 3190.385 ;
        RECT 1053.005 3190.070 1100.255 3190.370 ;
        RECT 1053.005 3190.055 1053.335 3190.070 ;
        RECT 1099.925 3190.055 1100.255 3190.070 ;
        RECT 1149.350 3190.370 1149.730 3190.380 ;
        RECT 1288.270 3190.370 1288.650 3190.380 ;
        RECT 1149.350 3190.070 1288.650 3190.370 ;
        RECT 1149.350 3190.060 1149.730 3190.070 ;
        RECT 1288.270 3190.060 1288.650 3190.070 ;
        RECT 1338.870 3189.690 1339.250 3189.700 ;
        RECT 1385.790 3189.690 1386.170 3189.700 ;
        RECT 1338.870 3189.390 1386.170 3189.690 ;
        RECT 1338.870 3189.380 1339.250 3189.390 ;
        RECT 1385.790 3189.380 1386.170 3189.390 ;
        RECT 1386.710 3189.010 1387.090 3189.020 ;
        RECT 1434.550 3189.010 1434.930 3189.020 ;
        RECT 1386.710 3188.710 1434.930 3189.010 ;
        RECT 1386.710 3188.700 1387.090 3188.710 ;
        RECT 1434.550 3188.700 1434.930 3188.710 ;
        RECT -4.800 2980.250 2.400 2980.700 ;
        RECT 15.705 2980.250 16.035 2980.265 ;
        RECT -4.800 2979.950 16.035 2980.250 ;
        RECT -4.800 2979.500 2.400 2979.950 ;
        RECT 15.705 2979.935 16.035 2979.950 ;
      LAYER via3 ;
        RECT 2043.620 3196.180 2043.940 3196.500 ;
        RECT 1288.300 3194.820 1288.620 3195.140 ;
        RECT 1149.380 3194.140 1149.700 3194.460 ;
        RECT 1385.820 3194.820 1386.140 3195.140 ;
        RECT 1434.580 3194.820 1434.900 3195.140 ;
        RECT 1338.900 3194.140 1339.220 3194.460 ;
        RECT 1386.740 3194.140 1387.060 3194.460 ;
        RECT 1775.900 3194.820 1776.220 3195.140 ;
        RECT 1811.780 3194.820 1812.100 3195.140 ;
        RECT 1872.500 3194.820 1872.820 3195.140 ;
        RECT 1775.900 3193.460 1776.220 3193.780 ;
        RECT 1811.780 3193.460 1812.100 3193.780 ;
        RECT 1872.500 3193.460 1872.820 3193.780 ;
        RECT 2043.620 3193.460 2043.940 3193.780 ;
        RECT 1149.380 3190.060 1149.700 3190.380 ;
        RECT 1288.300 3190.060 1288.620 3190.380 ;
        RECT 1338.900 3189.380 1339.220 3189.700 ;
        RECT 1385.820 3189.380 1386.140 3189.700 ;
        RECT 1386.740 3188.700 1387.060 3189.020 ;
        RECT 1434.580 3188.700 1434.900 3189.020 ;
      LAYER met4 ;
        RECT 2043.615 3196.175 2043.945 3196.505 ;
        RECT 1288.295 3194.815 1288.625 3195.145 ;
        RECT 1385.815 3194.815 1386.145 3195.145 ;
        RECT 1434.575 3194.815 1434.905 3195.145 ;
        RECT 1775.895 3194.815 1776.225 3195.145 ;
        RECT 1811.775 3194.815 1812.105 3195.145 ;
        RECT 1872.495 3194.815 1872.825 3195.145 ;
        RECT 1149.375 3194.135 1149.705 3194.465 ;
        RECT 1149.390 3190.385 1149.690 3194.135 ;
        RECT 1288.310 3190.385 1288.610 3194.815 ;
        RECT 1338.895 3194.135 1339.225 3194.465 ;
        RECT 1149.375 3190.055 1149.705 3190.385 ;
        RECT 1288.295 3190.055 1288.625 3190.385 ;
        RECT 1338.910 3189.705 1339.210 3194.135 ;
        RECT 1385.830 3189.705 1386.130 3194.815 ;
        RECT 1386.735 3194.135 1387.065 3194.465 ;
        RECT 1338.895 3189.375 1339.225 3189.705 ;
        RECT 1385.815 3189.375 1386.145 3189.705 ;
        RECT 1386.750 3189.025 1387.050 3194.135 ;
        RECT 1434.590 3189.025 1434.890 3194.815 ;
        RECT 1775.910 3193.785 1776.210 3194.815 ;
        RECT 1811.790 3193.785 1812.090 3194.815 ;
        RECT 1872.510 3193.785 1872.810 3194.815 ;
        RECT 2043.630 3193.785 2043.930 3196.175 ;
        RECT 1775.895 3193.455 1776.225 3193.785 ;
        RECT 1811.775 3193.455 1812.105 3193.785 ;
        RECT 1872.495 3193.455 1872.825 3193.785 ;
        RECT 2043.615 3193.455 2043.945 3193.785 ;
        RECT 1386.735 3188.695 1387.065 3189.025 ;
        RECT 1434.575 3188.695 1434.905 3189.025 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.170 3212.560 16.490 3212.620 ;
        RECT 2194.270 3212.560 2194.590 3212.620 ;
        RECT 16.170 3212.420 2194.590 3212.560 ;
        RECT 16.170 3212.360 16.490 3212.420 ;
        RECT 2194.270 3212.360 2194.590 3212.420 ;
      LAYER via ;
        RECT 16.200 3212.360 16.460 3212.620 ;
        RECT 2194.300 3212.360 2194.560 3212.620 ;
      LAYER met2 ;
        RECT 16.200 3212.330 16.460 3212.650 ;
        RECT 2194.300 3212.330 2194.560 3212.650 ;
        RECT 16.260 2693.325 16.400 3212.330 ;
        RECT 2194.360 3200.000 2194.500 3212.330 ;
        RECT 2194.220 3196.000 2194.500 3200.000 ;
        RECT 16.190 2692.955 16.470 2693.325 ;
      LAYER via2 ;
        RECT 16.190 2693.000 16.470 2693.280 ;
      LAYER met3 ;
        RECT -4.800 2693.290 2.400 2693.740 ;
        RECT 16.165 2693.290 16.495 2693.305 ;
        RECT -4.800 2692.990 16.495 2693.290 ;
        RECT -4.800 2692.540 2.400 2692.990 ;
        RECT 16.165 2692.975 16.495 2692.990 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 40.090 3212.220 40.410 3212.280 ;
        RECT 2233.830 3212.220 2234.150 3212.280 ;
        RECT 40.090 3212.080 2234.150 3212.220 ;
        RECT 40.090 3212.020 40.410 3212.080 ;
        RECT 2233.830 3212.020 2234.150 3212.080 ;
        RECT 16.170 2406.420 16.490 2406.480 ;
        RECT 40.090 2406.420 40.410 2406.480 ;
        RECT 16.170 2406.280 40.410 2406.420 ;
        RECT 16.170 2406.220 16.490 2406.280 ;
        RECT 40.090 2406.220 40.410 2406.280 ;
      LAYER via ;
        RECT 40.120 3212.020 40.380 3212.280 ;
        RECT 2233.860 3212.020 2234.120 3212.280 ;
        RECT 16.200 2406.220 16.460 2406.480 ;
        RECT 40.120 2406.220 40.380 2406.480 ;
      LAYER met2 ;
        RECT 40.120 3211.990 40.380 3212.310 ;
        RECT 2233.860 3211.990 2234.120 3212.310 ;
        RECT 40.180 2406.510 40.320 3211.990 ;
        RECT 2233.920 3200.000 2234.060 3211.990 ;
        RECT 2233.780 3196.000 2234.060 3200.000 ;
        RECT 16.200 2406.190 16.460 2406.510 ;
        RECT 40.120 2406.190 40.380 2406.510 ;
        RECT 16.260 2405.685 16.400 2406.190 ;
        RECT 16.190 2405.315 16.470 2405.685 ;
      LAYER via2 ;
        RECT 16.190 2405.360 16.470 2405.640 ;
      LAYER met3 ;
        RECT -4.800 2405.650 2.400 2406.100 ;
        RECT 16.165 2405.650 16.495 2405.665 ;
        RECT -4.800 2405.350 16.495 2405.650 ;
        RECT -4.800 2404.900 2.400 2405.350 ;
        RECT 16.165 2405.335 16.495 2405.350 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 39.630 3211.540 39.950 3211.600 ;
        RECT 2273.390 3211.540 2273.710 3211.600 ;
        RECT 39.630 3211.400 2273.710 3211.540 ;
        RECT 39.630 3211.340 39.950 3211.400 ;
        RECT 2273.390 3211.340 2273.710 3211.400 ;
        RECT 16.170 2121.500 16.490 2121.560 ;
        RECT 39.630 2121.500 39.950 2121.560 ;
        RECT 16.170 2121.360 39.950 2121.500 ;
        RECT 16.170 2121.300 16.490 2121.360 ;
        RECT 39.630 2121.300 39.950 2121.360 ;
      LAYER via ;
        RECT 39.660 3211.340 39.920 3211.600 ;
        RECT 2273.420 3211.340 2273.680 3211.600 ;
        RECT 16.200 2121.300 16.460 2121.560 ;
        RECT 39.660 2121.300 39.920 2121.560 ;
      LAYER met2 ;
        RECT 39.660 3211.310 39.920 3211.630 ;
        RECT 2273.420 3211.310 2273.680 3211.630 ;
        RECT 39.720 2121.590 39.860 3211.310 ;
        RECT 2273.480 3200.000 2273.620 3211.310 ;
        RECT 2273.340 3196.000 2273.620 3200.000 ;
        RECT 16.200 2121.270 16.460 2121.590 ;
        RECT 39.660 2121.270 39.920 2121.590 ;
        RECT 16.260 2118.725 16.400 2121.270 ;
        RECT 16.190 2118.355 16.470 2118.725 ;
      LAYER via2 ;
        RECT 16.190 2118.400 16.470 2118.680 ;
      LAYER met3 ;
        RECT -4.800 2118.690 2.400 2119.140 ;
        RECT 16.165 2118.690 16.495 2118.705 ;
        RECT -4.800 2118.390 16.495 2118.690 ;
        RECT -4.800 2117.940 2.400 2118.390 ;
        RECT 16.165 2118.375 16.495 2118.390 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 13.870 1833.860 14.190 1833.920 ;
        RECT 25.370 1833.860 25.690 1833.920 ;
        RECT 13.870 1833.720 25.690 1833.860 ;
        RECT 13.870 1833.660 14.190 1833.720 ;
        RECT 25.370 1833.660 25.690 1833.720 ;
      LAYER via ;
        RECT 13.900 1833.660 14.160 1833.920 ;
        RECT 25.400 1833.660 25.660 1833.920 ;
      LAYER met2 ;
        RECT 2311.590 3196.410 2311.870 3196.525 ;
        RECT 2312.900 3196.410 2313.180 3200.000 ;
        RECT 2311.590 3196.270 2313.180 3196.410 ;
        RECT 2311.590 3196.155 2311.870 3196.270 ;
        RECT 2312.900 3196.000 2313.180 3196.270 ;
        RECT 25.390 3192.755 25.670 3193.125 ;
        RECT 25.460 1833.950 25.600 3192.755 ;
        RECT 13.900 1833.630 14.160 1833.950 ;
        RECT 25.400 1833.630 25.660 1833.950 ;
        RECT 13.960 1831.085 14.100 1833.630 ;
        RECT 13.890 1830.715 14.170 1831.085 ;
      LAYER via2 ;
        RECT 2311.590 3196.200 2311.870 3196.480 ;
        RECT 25.390 3192.800 25.670 3193.080 ;
        RECT 13.890 1830.760 14.170 1831.040 ;
      LAYER met3 ;
        RECT 2311.565 3196.500 2311.895 3196.505 ;
        RECT 2311.310 3196.490 2311.895 3196.500 ;
        RECT 2311.110 3196.190 2311.895 3196.490 ;
        RECT 2311.310 3196.180 2311.895 3196.190 ;
        RECT 2311.565 3196.175 2311.895 3196.180 ;
        RECT 1666.390 3195.810 1666.770 3195.820 ;
        RECT 1682.030 3195.810 1682.410 3195.820 ;
        RECT 1666.390 3195.510 1682.410 3195.810 ;
        RECT 1666.390 3195.500 1666.770 3195.510 ;
        RECT 1682.030 3195.500 1682.410 3195.510 ;
        RECT 25.365 3193.090 25.695 3193.105 ;
        RECT 1666.390 3193.090 1666.770 3193.100 ;
        RECT 25.365 3192.790 1666.770 3193.090 ;
        RECT 25.365 3192.775 25.695 3192.790 ;
        RECT 1666.390 3192.780 1666.770 3192.790 ;
        RECT 1682.030 3193.090 1682.410 3193.100 ;
        RECT 2311.310 3193.090 2311.690 3193.100 ;
        RECT 1682.030 3192.790 1822.210 3193.090 ;
        RECT 1682.030 3192.780 1682.410 3192.790 ;
        RECT 1821.910 3192.410 1822.210 3192.790 ;
        RECT 1823.750 3192.790 2311.690 3193.090 ;
        RECT 1823.750 3192.410 1824.050 3192.790 ;
        RECT 2311.310 3192.780 2311.690 3192.790 ;
        RECT 1821.910 3192.110 1824.050 3192.410 ;
        RECT -4.800 1831.050 2.400 1831.500 ;
        RECT 13.865 1831.050 14.195 1831.065 ;
        RECT -4.800 1830.750 14.195 1831.050 ;
        RECT -4.800 1830.300 2.400 1830.750 ;
        RECT 13.865 1830.735 14.195 1830.750 ;
      LAYER via3 ;
        RECT 2311.340 3196.180 2311.660 3196.500 ;
        RECT 1666.420 3195.500 1666.740 3195.820 ;
        RECT 1682.060 3195.500 1682.380 3195.820 ;
        RECT 1666.420 3192.780 1666.740 3193.100 ;
        RECT 1682.060 3192.780 1682.380 3193.100 ;
        RECT 2311.340 3192.780 2311.660 3193.100 ;
      LAYER met4 ;
        RECT 2311.335 3196.175 2311.665 3196.505 ;
        RECT 1666.415 3195.495 1666.745 3195.825 ;
        RECT 1682.055 3195.495 1682.385 3195.825 ;
        RECT 1666.430 3193.105 1666.730 3195.495 ;
        RECT 1682.070 3193.105 1682.370 3195.495 ;
        RECT 2311.350 3193.105 2311.650 3196.175 ;
        RECT 1666.415 3192.775 1666.745 3193.105 ;
        RECT 1682.055 3192.775 1682.385 3193.105 ;
        RECT 2311.335 3192.775 2311.665 3193.105 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1490.010 670.720 1490.330 670.780 ;
        RECT 1507.950 670.720 1508.270 670.780 ;
        RECT 1490.010 670.580 1508.270 670.720 ;
        RECT 1490.010 670.520 1490.330 670.580 ;
        RECT 1507.950 670.520 1508.270 670.580 ;
        RECT 1918.270 670.380 1918.590 670.440 ;
        RECT 1926.090 670.380 1926.410 670.440 ;
        RECT 1918.270 670.240 1926.410 670.380 ;
        RECT 1918.270 670.180 1918.590 670.240 ;
        RECT 1926.090 670.180 1926.410 670.240 ;
        RECT 2608.270 669.700 2608.590 669.760 ;
        RECT 2632.190 669.700 2632.510 669.760 ;
        RECT 2608.270 669.560 2632.510 669.700 ;
        RECT 2608.270 669.500 2608.590 669.560 ;
        RECT 2632.190 669.500 2632.510 669.560 ;
      LAYER via ;
        RECT 1490.040 670.520 1490.300 670.780 ;
        RECT 1507.980 670.520 1508.240 670.780 ;
        RECT 1918.300 670.180 1918.560 670.440 ;
        RECT 1926.120 670.180 1926.380 670.440 ;
        RECT 2608.300 669.500 2608.560 669.760 ;
        RECT 2632.220 669.500 2632.480 669.760 ;
      LAYER met2 ;
        RECT 1245.770 3196.410 1246.050 3196.525 ;
        RECT 1247.080 3196.410 1247.360 3200.000 ;
        RECT 1245.770 3196.270 1247.360 3196.410 ;
        RECT 1245.770 3196.155 1246.050 3196.270 ;
        RECT 1247.080 3196.000 1247.360 3196.270 ;
        RECT 1669.430 671.995 1669.710 672.365 ;
        RECT 1338.690 670.635 1338.970 671.005 ;
        RECT 1393.430 670.635 1393.710 671.005 ;
        RECT 1476.230 670.635 1476.510 671.005 ;
        RECT 1490.030 670.635 1490.310 671.005 ;
        RECT 1507.970 670.635 1508.250 671.005 ;
        RECT 1338.760 670.325 1338.900 670.635 ;
        RECT 1338.690 669.955 1338.970 670.325 ;
        RECT 1393.500 669.645 1393.640 670.635 ;
        RECT 1393.430 669.275 1393.710 669.645 ;
        RECT 1476.300 668.285 1476.440 670.635 ;
        RECT 1490.040 670.490 1490.300 670.635 ;
        RECT 1507.980 670.490 1508.240 670.635 ;
        RECT 1669.500 670.325 1669.640 671.995 ;
        RECT 2014.430 671.315 2014.710 671.685 ;
        RECT 2028.230 671.570 2028.510 671.685 ;
        RECT 2028.230 671.430 2028.900 671.570 ;
        RECT 2028.230 671.315 2028.510 671.430 ;
        RECT 1926.110 670.635 1926.390 671.005 ;
        RECT 1926.180 670.470 1926.320 670.635 ;
        RECT 1918.300 670.325 1918.560 670.470 ;
        RECT 1537.870 670.210 1538.150 670.325 ;
        RECT 1538.790 670.210 1539.070 670.325 ;
        RECT 1537.870 670.070 1539.070 670.210 ;
        RECT 1537.870 669.955 1538.150 670.070 ;
        RECT 1538.790 669.955 1539.070 670.070 ;
        RECT 1669.430 669.955 1669.710 670.325 ;
        RECT 1690.130 670.210 1690.410 670.325 ;
        RECT 1690.130 670.070 1690.800 670.210 ;
        RECT 1690.130 669.955 1690.410 670.070 ;
        RECT 1476.230 667.915 1476.510 668.285 ;
        RECT 1690.660 667.605 1690.800 670.070 ;
        RECT 1918.290 669.955 1918.570 670.325 ;
        RECT 1926.120 670.150 1926.380 670.470 ;
        RECT 2014.500 669.645 2014.640 671.315 ;
        RECT 2028.760 671.005 2028.900 671.430 ;
        RECT 2089.410 671.315 2089.690 671.685 ;
        RECT 2704.430 671.315 2704.710 671.685 ;
        RECT 2028.690 670.635 2028.970 671.005 ;
        RECT 2089.480 670.890 2089.620 671.315 ;
        RECT 2091.250 670.890 2091.530 671.005 ;
        RECT 2089.480 670.750 2091.530 670.890 ;
        RECT 2091.250 670.635 2091.530 670.750 ;
        RECT 2283.530 670.210 2283.810 670.325 ;
        RECT 2284.450 670.210 2284.730 670.325 ;
        RECT 2283.530 670.070 2284.730 670.210 ;
        RECT 2283.530 669.955 2283.810 670.070 ;
        RECT 2284.450 669.955 2284.730 670.070 ;
        RECT 2572.870 669.955 2573.150 670.325 ;
        RECT 2632.210 669.955 2632.490 670.325 ;
        RECT 2014.430 669.275 2014.710 669.645 ;
        RECT 2572.940 668.285 2573.080 669.955 ;
        RECT 2632.280 669.790 2632.420 669.955 ;
        RECT 2608.300 669.645 2608.560 669.790 ;
        RECT 2608.290 669.275 2608.570 669.645 ;
        RECT 2632.220 669.470 2632.480 669.790 ;
        RECT 2704.500 669.645 2704.640 671.315 ;
        RECT 2801.030 670.635 2801.310 671.005 ;
        RECT 2704.430 669.275 2704.710 669.645 ;
        RECT 2801.100 668.965 2801.240 670.635 ;
        RECT 2863.130 669.955 2863.410 670.325 ;
        RECT 2863.200 669.530 2863.340 669.955 ;
        RECT 2863.590 669.530 2863.870 669.645 ;
        RECT 2863.200 669.390 2863.870 669.530 ;
        RECT 2863.590 669.275 2863.870 669.390 ;
        RECT 2801.030 668.595 2801.310 668.965 ;
        RECT 2572.870 667.915 2573.150 668.285 ;
        RECT 1690.590 667.235 1690.870 667.605 ;
      LAYER via2 ;
        RECT 1245.770 3196.200 1246.050 3196.480 ;
        RECT 1669.430 672.040 1669.710 672.320 ;
        RECT 1338.690 670.680 1338.970 670.960 ;
        RECT 1393.430 670.680 1393.710 670.960 ;
        RECT 1476.230 670.680 1476.510 670.960 ;
        RECT 1490.030 670.680 1490.310 670.960 ;
        RECT 1507.970 670.680 1508.250 670.960 ;
        RECT 1338.690 670.000 1338.970 670.280 ;
        RECT 1393.430 669.320 1393.710 669.600 ;
        RECT 2014.430 671.360 2014.710 671.640 ;
        RECT 2028.230 671.360 2028.510 671.640 ;
        RECT 1926.110 670.680 1926.390 670.960 ;
        RECT 1537.870 670.000 1538.150 670.280 ;
        RECT 1538.790 670.000 1539.070 670.280 ;
        RECT 1669.430 670.000 1669.710 670.280 ;
        RECT 1690.130 670.000 1690.410 670.280 ;
        RECT 1476.230 667.960 1476.510 668.240 ;
        RECT 1918.290 670.000 1918.570 670.280 ;
        RECT 2089.410 671.360 2089.690 671.640 ;
        RECT 2704.430 671.360 2704.710 671.640 ;
        RECT 2028.690 670.680 2028.970 670.960 ;
        RECT 2091.250 670.680 2091.530 670.960 ;
        RECT 2283.530 670.000 2283.810 670.280 ;
        RECT 2284.450 670.000 2284.730 670.280 ;
        RECT 2572.870 670.000 2573.150 670.280 ;
        RECT 2632.210 670.000 2632.490 670.280 ;
        RECT 2014.430 669.320 2014.710 669.600 ;
        RECT 2608.290 669.320 2608.570 669.600 ;
        RECT 2801.030 670.680 2801.310 670.960 ;
        RECT 2704.430 669.320 2704.710 669.600 ;
        RECT 2863.130 670.000 2863.410 670.280 ;
        RECT 2863.590 669.320 2863.870 669.600 ;
        RECT 2801.030 668.640 2801.310 668.920 ;
        RECT 2572.870 667.960 2573.150 668.240 ;
        RECT 1690.590 667.280 1690.870 667.560 ;
      LAYER met3 ;
        RECT 1245.030 3196.490 1245.410 3196.500 ;
        RECT 1245.745 3196.490 1246.075 3196.505 ;
        RECT 1245.030 3196.190 1246.075 3196.490 ;
        RECT 1245.030 3196.180 1245.410 3196.190 ;
        RECT 1245.745 3196.175 1246.075 3196.190 ;
        RECT 2917.600 674.370 2924.800 674.820 ;
        RECT 2916.710 674.070 2924.800 674.370 ;
        RECT 1621.310 672.330 1621.690 672.340 ;
        RECT 1669.405 672.330 1669.735 672.345 ;
        RECT 1621.310 672.030 1669.735 672.330 ;
        RECT 1621.310 672.020 1621.690 672.030 ;
        RECT 1669.405 672.015 1669.735 672.030 ;
        RECT 2014.405 671.650 2014.735 671.665 ;
        RECT 2028.205 671.650 2028.535 671.665 ;
        RECT 2089.385 671.650 2089.715 671.665 ;
        RECT 2656.310 671.650 2656.690 671.660 ;
        RECT 2704.405 671.650 2704.735 671.665 ;
        RECT 2014.405 671.350 2028.535 671.650 ;
        RECT 2014.405 671.335 2014.735 671.350 ;
        RECT 2028.205 671.335 2028.535 671.350 ;
        RECT 2076.750 671.350 2089.715 671.650 ;
        RECT 1338.665 670.970 1338.995 670.985 ;
        RECT 1393.405 670.970 1393.735 670.985 ;
        RECT 1338.665 670.670 1393.735 670.970 ;
        RECT 1338.665 670.655 1338.995 670.670 ;
        RECT 1393.405 670.655 1393.735 670.670 ;
        RECT 1476.205 670.970 1476.535 670.985 ;
        RECT 1490.005 670.970 1490.335 670.985 ;
        RECT 1476.205 670.670 1490.335 670.970 ;
        RECT 1476.205 670.655 1476.535 670.670 ;
        RECT 1490.005 670.655 1490.335 670.670 ;
        RECT 1507.945 670.970 1508.275 670.985 ;
        RECT 1621.310 670.970 1621.690 670.980 ;
        RECT 1926.085 670.970 1926.415 670.985 ;
        RECT 1966.310 670.970 1966.690 670.980 ;
        RECT 1507.945 670.670 1532.410 670.970 ;
        RECT 1507.945 670.655 1508.275 670.670 ;
        RECT 1338.665 670.290 1338.995 670.305 ;
        RECT 1268.990 669.990 1338.995 670.290 ;
        RECT 1532.110 670.290 1532.410 670.670 ;
        RECT 1618.590 670.670 1621.690 670.970 ;
        RECT 1537.845 670.290 1538.175 670.305 ;
        RECT 1532.110 669.990 1538.175 670.290 ;
        RECT 1245.030 669.610 1245.410 669.620 ;
        RECT 1268.990 669.610 1269.290 669.990 ;
        RECT 1338.665 669.975 1338.995 669.990 ;
        RECT 1537.845 669.975 1538.175 669.990 ;
        RECT 1538.765 670.290 1539.095 670.305 ;
        RECT 1593.710 670.290 1594.090 670.300 ;
        RECT 1538.765 669.990 1594.090 670.290 ;
        RECT 1538.765 669.975 1539.095 669.990 ;
        RECT 1593.710 669.980 1594.090 669.990 ;
        RECT 1245.030 669.310 1269.290 669.610 ;
        RECT 1393.405 669.610 1393.735 669.625 ;
        RECT 1428.110 669.610 1428.490 669.620 ;
        RECT 1393.405 669.310 1428.490 669.610 ;
        RECT 1245.030 669.300 1245.410 669.310 ;
        RECT 1393.405 669.295 1393.735 669.310 ;
        RECT 1428.110 669.300 1428.490 669.310 ;
        RECT 1593.710 668.930 1594.090 668.940 ;
        RECT 1618.590 668.930 1618.890 670.670 ;
        RECT 1621.310 670.660 1621.690 670.670 ;
        RECT 1835.710 670.670 1877.410 670.970 ;
        RECT 1669.405 670.290 1669.735 670.305 ;
        RECT 1690.105 670.290 1690.435 670.305 ;
        RECT 1669.405 669.990 1690.435 670.290 ;
        RECT 1669.405 669.975 1669.735 669.990 ;
        RECT 1690.105 669.975 1690.435 669.990 ;
        RECT 1786.910 669.610 1787.290 669.620 ;
        RECT 1835.710 669.610 1836.010 670.670 ;
        RECT 1877.110 670.290 1877.410 670.670 ;
        RECT 1926.085 670.670 1966.690 670.970 ;
        RECT 1926.085 670.655 1926.415 670.670 ;
        RECT 1966.310 670.660 1966.690 670.670 ;
        RECT 2028.665 670.970 2028.995 670.985 ;
        RECT 2076.750 670.970 2077.050 671.350 ;
        RECT 2089.385 671.335 2089.715 671.350 ;
        RECT 2463.150 671.350 2511.290 671.650 ;
        RECT 2028.665 670.670 2077.050 670.970 ;
        RECT 2091.225 670.970 2091.555 670.985 ;
        RECT 2091.225 670.670 2138.690 670.970 ;
        RECT 2028.665 670.655 2028.995 670.670 ;
        RECT 2091.225 670.655 2091.555 670.670 ;
        RECT 1918.265 670.290 1918.595 670.305 ;
        RECT 1877.110 669.990 1918.595 670.290 ;
        RECT 1918.265 669.975 1918.595 669.990 ;
        RECT 1786.910 669.310 1836.010 669.610 ;
        RECT 1966.310 669.610 1966.690 669.620 ;
        RECT 2014.405 669.610 2014.735 669.625 ;
        RECT 1966.310 669.310 2014.735 669.610 ;
        RECT 2138.390 669.610 2138.690 670.670 ;
        RECT 2139.310 670.670 2187.450 670.970 ;
        RECT 2139.310 669.610 2139.610 670.670 ;
        RECT 2138.390 669.310 2139.610 669.610 ;
        RECT 2187.150 669.610 2187.450 670.670 ;
        RECT 2283.505 670.290 2283.835 670.305 ;
        RECT 2235.910 669.990 2283.835 670.290 ;
        RECT 2235.910 669.610 2236.210 669.990 ;
        RECT 2283.505 669.975 2283.835 669.990 ;
        RECT 2284.425 670.290 2284.755 670.305 ;
        RECT 2366.510 670.290 2366.890 670.300 ;
        RECT 2463.150 670.290 2463.450 671.350 ;
        RECT 2510.990 670.980 2511.290 671.350 ;
        RECT 2656.310 671.350 2704.735 671.650 ;
        RECT 2656.310 671.340 2656.690 671.350 ;
        RECT 2704.405 671.335 2704.735 671.350 ;
        RECT 2510.950 670.660 2511.330 670.980 ;
        RECT 2801.005 670.970 2801.335 670.985 ;
        RECT 2801.005 670.670 2815.810 670.970 ;
        RECT 2801.005 670.655 2801.335 670.670 ;
        RECT 2572.845 670.290 2573.175 670.305 ;
        RECT 2284.425 669.990 2331.890 670.290 ;
        RECT 2284.425 669.975 2284.755 669.990 ;
        RECT 2187.150 669.310 2236.210 669.610 ;
        RECT 2331.590 669.610 2331.890 669.990 ;
        RECT 2332.510 669.990 2366.890 670.290 ;
        RECT 2332.510 669.610 2332.810 669.990 ;
        RECT 2366.510 669.980 2366.890 669.990 ;
        RECT 2429.110 669.990 2463.450 670.290 ;
        RECT 2525.710 669.990 2573.175 670.290 ;
        RECT 2429.110 669.610 2429.410 669.990 ;
        RECT 2331.590 669.310 2332.810 669.610 ;
        RECT 2414.390 669.310 2429.410 669.610 ;
        RECT 2510.950 669.610 2511.330 669.620 ;
        RECT 2525.710 669.610 2526.010 669.990 ;
        RECT 2572.845 669.975 2573.175 669.990 ;
        RECT 2632.185 670.290 2632.515 670.305 ;
        RECT 2656.310 670.290 2656.690 670.300 ;
        RECT 2752.910 670.290 2753.290 670.300 ;
        RECT 2632.185 669.990 2656.690 670.290 ;
        RECT 2632.185 669.975 2632.515 669.990 ;
        RECT 2656.310 669.980 2656.690 669.990 ;
        RECT 2718.910 669.990 2753.290 670.290 ;
        RECT 2608.265 669.610 2608.595 669.625 ;
        RECT 2510.950 669.310 2526.010 669.610 ;
        RECT 2607.590 669.310 2608.595 669.610 ;
        RECT 1786.910 669.300 1787.290 669.310 ;
        RECT 1966.310 669.300 1966.690 669.310 ;
        RECT 2014.405 669.295 2014.735 669.310 ;
        RECT 1593.710 668.630 1618.890 668.930 ;
        RECT 1593.710 668.620 1594.090 668.630 ;
        RECT 1428.110 668.250 1428.490 668.260 ;
        RECT 1476.205 668.250 1476.535 668.265 ;
        RECT 1786.910 668.250 1787.290 668.260 ;
        RECT 1428.110 667.950 1476.535 668.250 ;
        RECT 1428.110 667.940 1428.490 667.950 ;
        RECT 1476.205 667.935 1476.535 667.950 ;
        RECT 1740.030 667.950 1787.290 668.250 ;
        RECT 1690.565 667.570 1690.895 667.585 ;
        RECT 1740.030 667.570 1740.330 667.950 ;
        RECT 1786.910 667.940 1787.290 667.950 ;
        RECT 2366.510 668.250 2366.890 668.260 ;
        RECT 2414.390 668.250 2414.690 669.310 ;
        RECT 2510.950 669.300 2511.330 669.310 ;
        RECT 2366.510 667.950 2414.690 668.250 ;
        RECT 2572.845 668.250 2573.175 668.265 ;
        RECT 2607.590 668.250 2607.890 669.310 ;
        RECT 2608.265 669.295 2608.595 669.310 ;
        RECT 2704.405 669.610 2704.735 669.625 ;
        RECT 2718.910 669.610 2719.210 669.990 ;
        RECT 2752.910 669.980 2753.290 669.990 ;
        RECT 2704.405 669.310 2719.210 669.610 ;
        RECT 2815.510 669.610 2815.810 670.670 ;
        RECT 2863.105 670.290 2863.435 670.305 ;
        RECT 2916.710 670.290 2917.010 674.070 ;
        RECT 2917.600 673.620 2924.800 674.070 ;
        RECT 2849.550 669.990 2863.435 670.290 ;
        RECT 2849.550 669.610 2849.850 669.990 ;
        RECT 2863.105 669.975 2863.435 669.990 ;
        RECT 2884.510 669.990 2917.010 670.290 ;
        RECT 2815.510 669.310 2849.850 669.610 ;
        RECT 2863.565 669.610 2863.895 669.625 ;
        RECT 2884.510 669.610 2884.810 669.990 ;
        RECT 2863.565 669.310 2884.810 669.610 ;
        RECT 2704.405 669.295 2704.735 669.310 ;
        RECT 2863.565 669.295 2863.895 669.310 ;
        RECT 2752.910 668.930 2753.290 668.940 ;
        RECT 2801.005 668.930 2801.335 668.945 ;
        RECT 2752.910 668.630 2801.335 668.930 ;
        RECT 2752.910 668.620 2753.290 668.630 ;
        RECT 2801.005 668.615 2801.335 668.630 ;
        RECT 2572.845 667.950 2607.890 668.250 ;
        RECT 2366.510 667.940 2366.890 667.950 ;
        RECT 2572.845 667.935 2573.175 667.950 ;
        RECT 1690.565 667.270 1740.330 667.570 ;
        RECT 1690.565 667.255 1690.895 667.270 ;
      LAYER via3 ;
        RECT 1245.060 3196.180 1245.380 3196.500 ;
        RECT 1621.340 672.020 1621.660 672.340 ;
        RECT 1245.060 669.300 1245.380 669.620 ;
        RECT 1593.740 669.980 1594.060 670.300 ;
        RECT 1428.140 669.300 1428.460 669.620 ;
        RECT 1593.740 668.620 1594.060 668.940 ;
        RECT 1621.340 670.660 1621.660 670.980 ;
        RECT 1786.940 669.300 1787.260 669.620 ;
        RECT 1966.340 670.660 1966.660 670.980 ;
        RECT 1966.340 669.300 1966.660 669.620 ;
        RECT 2366.540 669.980 2366.860 670.300 ;
        RECT 2656.340 671.340 2656.660 671.660 ;
        RECT 2510.980 670.660 2511.300 670.980 ;
        RECT 1428.140 667.940 1428.460 668.260 ;
        RECT 1786.940 667.940 1787.260 668.260 ;
        RECT 2366.540 667.940 2366.860 668.260 ;
        RECT 2510.980 669.300 2511.300 669.620 ;
        RECT 2656.340 669.980 2656.660 670.300 ;
        RECT 2752.940 669.980 2753.260 670.300 ;
        RECT 2752.940 668.620 2753.260 668.940 ;
      LAYER met4 ;
        RECT 1245.055 3196.175 1245.385 3196.505 ;
        RECT 1245.070 669.625 1245.370 3196.175 ;
        RECT 1621.335 672.015 1621.665 672.345 ;
        RECT 1621.350 670.985 1621.650 672.015 ;
        RECT 2656.335 671.335 2656.665 671.665 ;
        RECT 1621.335 670.655 1621.665 670.985 ;
        RECT 1966.335 670.655 1966.665 670.985 ;
        RECT 2510.975 670.655 2511.305 670.985 ;
        RECT 1593.735 669.975 1594.065 670.305 ;
        RECT 1245.055 669.295 1245.385 669.625 ;
        RECT 1428.135 669.295 1428.465 669.625 ;
        RECT 1428.150 668.265 1428.450 669.295 ;
        RECT 1593.750 668.945 1594.050 669.975 ;
        RECT 1966.350 669.625 1966.650 670.655 ;
        RECT 2366.535 669.975 2366.865 670.305 ;
        RECT 1786.935 669.295 1787.265 669.625 ;
        RECT 1966.335 669.295 1966.665 669.625 ;
        RECT 1593.735 668.615 1594.065 668.945 ;
        RECT 1786.950 668.265 1787.250 669.295 ;
        RECT 2366.550 668.265 2366.850 669.975 ;
        RECT 2510.990 669.625 2511.290 670.655 ;
        RECT 2656.350 670.305 2656.650 671.335 ;
        RECT 2656.335 669.975 2656.665 670.305 ;
        RECT 2752.935 669.975 2753.265 670.305 ;
        RECT 2510.975 669.295 2511.305 669.625 ;
        RECT 2752.950 668.945 2753.250 669.975 ;
        RECT 2752.935 668.615 2753.265 668.945 ;
        RECT 1428.135 667.935 1428.465 668.265 ;
        RECT 1786.935 667.935 1787.265 668.265 ;
        RECT 2366.535 667.935 2366.865 668.265 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 24.910 3210.520 25.230 3210.580 ;
        RECT 2352.510 3210.520 2352.830 3210.580 ;
        RECT 24.910 3210.380 2352.830 3210.520 ;
        RECT 24.910 3210.320 25.230 3210.380 ;
        RECT 2352.510 3210.320 2352.830 3210.380 ;
        RECT 13.870 1544.180 14.190 1544.240 ;
        RECT 24.910 1544.180 25.230 1544.240 ;
        RECT 13.870 1544.040 25.230 1544.180 ;
        RECT 13.870 1543.980 14.190 1544.040 ;
        RECT 24.910 1543.980 25.230 1544.040 ;
      LAYER via ;
        RECT 24.940 3210.320 25.200 3210.580 ;
        RECT 2352.540 3210.320 2352.800 3210.580 ;
        RECT 13.900 1543.980 14.160 1544.240 ;
        RECT 24.940 1543.980 25.200 1544.240 ;
      LAYER met2 ;
        RECT 24.940 3210.290 25.200 3210.610 ;
        RECT 2352.540 3210.290 2352.800 3210.610 ;
        RECT 25.000 1544.270 25.140 3210.290 ;
        RECT 2352.600 3200.000 2352.740 3210.290 ;
        RECT 2352.460 3196.000 2352.740 3200.000 ;
        RECT 13.900 1544.125 14.160 1544.270 ;
        RECT 13.890 1543.755 14.170 1544.125 ;
        RECT 24.940 1543.950 25.200 1544.270 ;
      LAYER via2 ;
        RECT 13.890 1543.800 14.170 1544.080 ;
      LAYER met3 ;
        RECT -4.800 1544.090 2.400 1544.540 ;
        RECT 13.865 1544.090 14.195 1544.105 ;
        RECT -4.800 1543.790 14.195 1544.090 ;
        RECT -4.800 1543.340 2.400 1543.790 ;
        RECT 13.865 1543.775 14.195 1543.790 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2391.630 3212.475 2391.910 3212.845 ;
        RECT 2391.700 3200.000 2391.840 3212.475 ;
        RECT 2391.560 3196.000 2391.840 3200.000 ;
      LAYER via2 ;
        RECT 2391.630 3212.520 2391.910 3212.800 ;
      LAYER met3 ;
        RECT 1309.430 3212.810 1309.810 3212.820 ;
        RECT 2391.605 3212.810 2391.935 3212.825 ;
        RECT 1309.430 3212.510 2391.935 3212.810 ;
        RECT 1309.430 3212.500 1309.810 3212.510 ;
        RECT 2391.605 3212.495 2391.935 3212.510 ;
        RECT 1309.430 1331.250 1309.810 1331.260 ;
        RECT 3.070 1330.950 1309.810 1331.250 ;
        RECT -4.800 1328.530 2.400 1328.980 ;
        RECT 3.070 1328.530 3.370 1330.950 ;
        RECT 1309.430 1330.940 1309.810 1330.950 ;
        RECT -4.800 1328.230 3.370 1328.530 ;
        RECT -4.800 1327.780 2.400 1328.230 ;
      LAYER via3 ;
        RECT 1309.460 3212.500 1309.780 3212.820 ;
        RECT 1309.460 1330.940 1309.780 1331.260 ;
      LAYER met4 ;
        RECT 1309.455 3212.495 1309.785 3212.825 ;
        RECT 1309.470 1331.265 1309.770 3212.495 ;
        RECT 1309.455 1330.935 1309.785 1331.265 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 20.310 3209.840 20.630 3209.900 ;
        RECT 2431.170 3209.840 2431.490 3209.900 ;
        RECT 20.310 3209.700 2431.490 3209.840 ;
        RECT 20.310 3209.640 20.630 3209.700 ;
        RECT 2431.170 3209.640 2431.490 3209.700 ;
      LAYER via ;
        RECT 20.340 3209.640 20.600 3209.900 ;
        RECT 2431.200 3209.640 2431.460 3209.900 ;
      LAYER met2 ;
        RECT 20.340 3209.610 20.600 3209.930 ;
        RECT 2431.200 3209.610 2431.460 3209.930 ;
        RECT 20.400 1113.005 20.540 3209.610 ;
        RECT 2431.260 3200.000 2431.400 3209.610 ;
        RECT 2431.120 3196.000 2431.400 3200.000 ;
        RECT 20.330 1112.635 20.610 1113.005 ;
      LAYER via2 ;
        RECT 20.330 1112.680 20.610 1112.960 ;
      LAYER met3 ;
        RECT -4.800 1112.970 2.400 1113.420 ;
        RECT 20.305 1112.970 20.635 1112.985 ;
        RECT -4.800 1112.670 20.635 1112.970 ;
        RECT -4.800 1112.220 2.400 1112.670 ;
        RECT 20.305 1112.655 20.635 1112.670 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2470.750 3210.435 2471.030 3210.805 ;
        RECT 2470.820 3200.000 2470.960 3210.435 ;
        RECT 2470.680 3196.000 2470.960 3200.000 ;
        RECT 16.650 903.195 16.930 903.565 ;
        RECT 16.720 897.445 16.860 903.195 ;
        RECT 16.650 897.075 16.930 897.445 ;
      LAYER via2 ;
        RECT 2470.750 3210.480 2471.030 3210.760 ;
        RECT 16.650 903.240 16.930 903.520 ;
        RECT 16.650 897.120 16.930 897.400 ;
      LAYER met3 ;
        RECT 1293.790 3210.770 1294.170 3210.780 ;
        RECT 2470.725 3210.770 2471.055 3210.785 ;
        RECT 1293.790 3210.470 2471.055 3210.770 ;
        RECT 1293.790 3210.460 1294.170 3210.470 ;
        RECT 2470.725 3210.455 2471.055 3210.470 ;
        RECT 16.625 903.530 16.955 903.545 ;
        RECT 1293.790 903.530 1294.170 903.540 ;
        RECT 16.625 903.230 1294.170 903.530 ;
        RECT 16.625 903.215 16.955 903.230 ;
        RECT 1293.790 903.220 1294.170 903.230 ;
        RECT -4.800 897.410 2.400 897.860 ;
        RECT 16.625 897.410 16.955 897.425 ;
        RECT -4.800 897.110 16.955 897.410 ;
        RECT -4.800 896.660 2.400 897.110 ;
        RECT 16.625 897.095 16.955 897.110 ;
      LAYER via3 ;
        RECT 1293.820 3210.460 1294.140 3210.780 ;
        RECT 1293.820 903.220 1294.140 903.540 ;
      LAYER met4 ;
        RECT 1293.815 3210.455 1294.145 3210.785 ;
        RECT 1293.830 903.545 1294.130 3210.455 ;
        RECT 1293.815 903.215 1294.145 903.545 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 19.390 3209.160 19.710 3209.220 ;
        RECT 2510.290 3209.160 2510.610 3209.220 ;
        RECT 19.390 3209.020 2510.610 3209.160 ;
        RECT 19.390 3208.960 19.710 3209.020 ;
        RECT 2510.290 3208.960 2510.610 3209.020 ;
      LAYER via ;
        RECT 19.420 3208.960 19.680 3209.220 ;
        RECT 2510.320 3208.960 2510.580 3209.220 ;
      LAYER met2 ;
        RECT 19.420 3208.930 19.680 3209.250 ;
        RECT 2510.320 3208.930 2510.580 3209.250 ;
        RECT 19.480 681.885 19.620 3208.930 ;
        RECT 2510.380 3200.000 2510.520 3208.930 ;
        RECT 2510.240 3196.000 2510.520 3200.000 ;
        RECT 19.410 681.515 19.690 681.885 ;
      LAYER via2 ;
        RECT 19.410 681.560 19.690 681.840 ;
      LAYER met3 ;
        RECT -4.800 681.850 2.400 682.300 ;
        RECT 19.385 681.850 19.715 681.865 ;
        RECT -4.800 681.550 19.715 681.850 ;
        RECT -4.800 681.100 2.400 681.550 ;
        RECT 19.385 681.535 19.715 681.550 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2548.950 3196.410 2549.230 3196.525 ;
        RECT 2549.800 3196.410 2550.080 3200.000 ;
        RECT 2548.950 3196.270 2550.080 3196.410 ;
        RECT 2548.950 3196.155 2549.230 3196.270 ;
        RECT 2549.800 3196.000 2550.080 3196.270 ;
        RECT 18.490 3191.395 18.770 3191.765 ;
        RECT 18.560 466.325 18.700 3191.395 ;
        RECT 18.490 465.955 18.770 466.325 ;
      LAYER via2 ;
        RECT 2548.950 3196.200 2549.230 3196.480 ;
        RECT 18.490 3191.440 18.770 3191.720 ;
        RECT 18.490 466.000 18.770 466.280 ;
      LAYER met3 ;
        RECT 2548.925 3196.500 2549.255 3196.505 ;
        RECT 2548.670 3196.490 2549.255 3196.500 ;
        RECT 2548.470 3196.190 2549.255 3196.490 ;
        RECT 2548.670 3196.180 2549.255 3196.190 ;
        RECT 2548.925 3196.175 2549.255 3196.180 ;
        RECT 18.465 3191.730 18.795 3191.745 ;
        RECT 2548.670 3191.730 2549.050 3191.740 ;
        RECT 18.465 3191.430 2549.050 3191.730 ;
        RECT 18.465 3191.415 18.795 3191.430 ;
        RECT 2548.670 3191.420 2549.050 3191.430 ;
        RECT -4.800 466.290 2.400 466.740 ;
        RECT 18.465 466.290 18.795 466.305 ;
        RECT -4.800 465.990 18.795 466.290 ;
        RECT -4.800 465.540 2.400 465.990 ;
        RECT 18.465 465.975 18.795 465.990 ;
      LAYER via3 ;
        RECT 2548.700 3196.180 2549.020 3196.500 ;
        RECT 2548.700 3191.420 2549.020 3191.740 ;
      LAYER met4 ;
        RECT 2548.695 3196.175 2549.025 3196.505 ;
        RECT 2548.710 3191.745 2549.010 3196.175 ;
        RECT 2548.695 3191.415 2549.025 3191.745 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 17.570 3214.515 17.850 3214.885 ;
        RECT 2588.970 3214.515 2589.250 3214.885 ;
        RECT 17.640 250.765 17.780 3214.515 ;
        RECT 2589.040 3200.000 2589.180 3214.515 ;
        RECT 2588.900 3196.000 2589.180 3200.000 ;
        RECT 17.570 250.395 17.850 250.765 ;
      LAYER via2 ;
        RECT 17.570 3214.560 17.850 3214.840 ;
        RECT 2588.970 3214.560 2589.250 3214.840 ;
        RECT 17.570 250.440 17.850 250.720 ;
      LAYER met3 ;
        RECT 17.545 3214.850 17.875 3214.865 ;
        RECT 2588.945 3214.850 2589.275 3214.865 ;
        RECT 17.545 3214.550 2589.275 3214.850 ;
        RECT 17.545 3214.535 17.875 3214.550 ;
        RECT 2588.945 3214.535 2589.275 3214.550 ;
        RECT -4.800 250.730 2.400 251.180 ;
        RECT 17.545 250.730 17.875 250.745 ;
        RECT -4.800 250.430 17.875 250.730 ;
        RECT -4.800 249.980 2.400 250.430 ;
        RECT 17.545 250.415 17.875 250.430 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2627.150 3196.410 2627.430 3196.525 ;
        RECT 2628.460 3196.410 2628.740 3200.000 ;
        RECT 2627.150 3196.270 2628.740 3196.410 ;
        RECT 2627.150 3196.155 2627.430 3196.270 ;
        RECT 2628.460 3196.000 2628.740 3196.270 ;
        RECT 17.110 3190.715 17.390 3191.085 ;
        RECT 17.180 35.885 17.320 3190.715 ;
        RECT 17.110 35.515 17.390 35.885 ;
      LAYER via2 ;
        RECT 2627.150 3196.200 2627.430 3196.480 ;
        RECT 17.110 3190.760 17.390 3191.040 ;
        RECT 17.110 35.560 17.390 35.840 ;
      LAYER met3 ;
        RECT 2627.125 3196.500 2627.455 3196.505 ;
        RECT 2626.870 3196.490 2627.455 3196.500 ;
        RECT 2626.670 3196.190 2627.455 3196.490 ;
        RECT 2626.870 3196.180 2627.455 3196.190 ;
        RECT 2627.125 3196.175 2627.455 3196.180 ;
        RECT 17.085 3191.050 17.415 3191.065 ;
        RECT 2626.870 3191.050 2627.250 3191.060 ;
        RECT 17.085 3190.750 2627.250 3191.050 ;
        RECT 17.085 3190.735 17.415 3190.750 ;
        RECT 2626.870 3190.740 2627.250 3190.750 ;
        RECT -4.800 35.850 2.400 36.300 ;
        RECT 17.085 35.850 17.415 35.865 ;
        RECT -4.800 35.550 17.415 35.850 ;
        RECT -4.800 35.100 2.400 35.550 ;
        RECT 17.085 35.535 17.415 35.550 ;
      LAYER via3 ;
        RECT 2626.900 3196.180 2627.220 3196.500 ;
        RECT 2626.900 3190.740 2627.220 3191.060 ;
      LAYER met4 ;
        RECT 2626.895 3196.175 2627.225 3196.505 ;
        RECT 2626.910 3191.065 2627.210 3196.175 ;
        RECT 2626.895 3190.735 2627.225 3191.065 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1863.070 906.000 1863.390 906.060 ;
        RECT 1910.910 906.000 1911.230 906.060 ;
        RECT 1863.070 905.860 1911.230 906.000 ;
        RECT 1863.070 905.800 1863.390 905.860 ;
        RECT 1910.910 905.800 1911.230 905.860 ;
        RECT 2766.510 904.980 2766.830 905.040 ;
        RECT 2774.790 904.980 2775.110 905.040 ;
        RECT 2766.510 904.840 2775.110 904.980 ;
        RECT 2766.510 904.780 2766.830 904.840 ;
        RECT 2774.790 904.780 2775.110 904.840 ;
        RECT 2379.650 904.640 2379.970 904.700 ;
        RECT 2380.570 904.640 2380.890 904.700 ;
        RECT 2379.650 904.500 2380.890 904.640 ;
        RECT 2379.650 904.440 2379.970 904.500 ;
        RECT 2380.570 904.440 2380.890 904.500 ;
        RECT 2125.270 904.300 2125.590 904.360 ;
        RECT 2172.650 904.300 2172.970 904.360 ;
        RECT 2125.270 904.160 2172.970 904.300 ;
        RECT 2125.270 904.100 2125.590 904.160 ;
        RECT 2172.650 904.100 2172.970 904.160 ;
        RECT 2608.270 904.300 2608.590 904.360 ;
        RECT 2632.190 904.300 2632.510 904.360 ;
        RECT 2608.270 904.160 2632.510 904.300 ;
        RECT 2608.270 904.100 2608.590 904.160 ;
        RECT 2632.190 904.100 2632.510 904.160 ;
      LAYER via ;
        RECT 1863.100 905.800 1863.360 906.060 ;
        RECT 1910.940 905.800 1911.200 906.060 ;
        RECT 2766.540 904.780 2766.800 905.040 ;
        RECT 2774.820 904.780 2775.080 905.040 ;
        RECT 2379.680 904.440 2379.940 904.700 ;
        RECT 2380.600 904.440 2380.860 904.700 ;
        RECT 2125.300 904.100 2125.560 904.360 ;
        RECT 2172.680 904.100 2172.940 904.360 ;
        RECT 2608.300 904.100 2608.560 904.360 ;
        RECT 2632.220 904.100 2632.480 904.360 ;
      LAYER met2 ;
        RECT 1286.640 3196.410 1286.920 3200.000 ;
        RECT 1288.550 3196.410 1288.830 3196.525 ;
        RECT 1286.640 3196.270 1288.830 3196.410 ;
        RECT 1286.640 3196.000 1286.920 3196.270 ;
        RECT 1288.550 3196.155 1288.830 3196.270 ;
        RECT 1717.730 906.595 1718.010 906.965 ;
        RECT 1717.800 906.285 1717.940 906.595 ;
        RECT 1545.230 905.915 1545.510 906.285 ;
        RECT 1717.730 905.915 1718.010 906.285 ;
        RECT 1863.090 905.915 1863.370 906.285 ;
        RECT 1545.300 904.245 1545.440 905.915 ;
        RECT 1863.100 905.770 1863.360 905.915 ;
        RECT 1910.940 905.770 1911.200 906.090 ;
        RECT 2704.430 905.915 2704.710 906.285 ;
        RECT 1911.000 904.925 1911.140 905.770 ;
        RECT 2172.670 905.235 2172.950 905.605 ;
        RECT 1855.730 904.555 1856.010 904.925 ;
        RECT 1910.930 904.555 1911.210 904.925 ;
        RECT 1545.230 903.875 1545.510 904.245 ;
        RECT 1855.800 903.565 1855.940 904.555 ;
        RECT 2172.740 904.390 2172.880 905.235 ;
        RECT 2379.670 904.555 2379.950 904.925 ;
        RECT 2380.590 904.555 2380.870 904.925 ;
        RECT 2572.870 904.555 2573.150 904.925 ;
        RECT 2632.210 904.555 2632.490 904.925 ;
        RECT 2379.680 904.410 2379.940 904.555 ;
        RECT 2380.600 904.410 2380.860 904.555 ;
        RECT 2125.300 904.245 2125.560 904.390 ;
        RECT 2125.290 903.875 2125.570 904.245 ;
        RECT 2172.680 904.070 2172.940 904.390 ;
        RECT 1855.730 903.195 1856.010 903.565 ;
        RECT 2572.940 902.885 2573.080 904.555 ;
        RECT 2632.280 904.390 2632.420 904.555 ;
        RECT 2608.300 904.245 2608.560 904.390 ;
        RECT 2608.290 903.875 2608.570 904.245 ;
        RECT 2632.220 904.070 2632.480 904.390 ;
        RECT 2704.500 904.245 2704.640 905.915 ;
        RECT 2766.540 904.925 2766.800 905.070 ;
        RECT 2774.820 904.925 2775.080 905.070 ;
        RECT 2766.530 904.555 2766.810 904.925 ;
        RECT 2774.810 904.555 2775.090 904.925 ;
        RECT 2704.430 903.875 2704.710 904.245 ;
        RECT 2572.870 902.515 2573.150 902.885 ;
      LAYER via2 ;
        RECT 1288.550 3196.200 1288.830 3196.480 ;
        RECT 1717.730 906.640 1718.010 906.920 ;
        RECT 1545.230 905.960 1545.510 906.240 ;
        RECT 1717.730 905.960 1718.010 906.240 ;
        RECT 1863.090 905.960 1863.370 906.240 ;
        RECT 2704.430 905.960 2704.710 906.240 ;
        RECT 2172.670 905.280 2172.950 905.560 ;
        RECT 1855.730 904.600 1856.010 904.880 ;
        RECT 1910.930 904.600 1911.210 904.880 ;
        RECT 1545.230 903.920 1545.510 904.200 ;
        RECT 2379.670 904.600 2379.950 904.880 ;
        RECT 2380.590 904.600 2380.870 904.880 ;
        RECT 2572.870 904.600 2573.150 904.880 ;
        RECT 2632.210 904.600 2632.490 904.880 ;
        RECT 2125.290 903.920 2125.570 904.200 ;
        RECT 1855.730 903.240 1856.010 903.520 ;
        RECT 2608.290 903.920 2608.570 904.200 ;
        RECT 2766.530 904.600 2766.810 904.880 ;
        RECT 2774.810 904.600 2775.090 904.880 ;
        RECT 2704.430 903.920 2704.710 904.200 ;
        RECT 2572.870 902.560 2573.150 902.840 ;
      LAYER met3 ;
        RECT 1288.525 3196.490 1288.855 3196.505 ;
        RECT 1289.190 3196.490 1289.570 3196.500 ;
        RECT 1288.525 3196.190 1289.570 3196.490 ;
        RECT 1288.525 3196.175 1288.855 3196.190 ;
        RECT 1289.190 3196.180 1289.570 3196.190 ;
        RECT 2917.600 909.650 2924.800 910.100 ;
        RECT 2916.710 909.350 2924.800 909.650 ;
        RECT 1717.705 906.940 1718.035 906.945 ;
        RECT 1717.705 906.930 1718.290 906.940 ;
        RECT 1717.500 906.630 1718.290 906.930 ;
        RECT 1717.705 906.620 1718.290 906.630 ;
        RECT 1717.705 906.615 1718.035 906.620 ;
        RECT 1545.205 906.250 1545.535 906.265 ;
        RECT 1717.705 906.250 1718.035 906.265 ;
        RECT 1863.065 906.250 1863.395 906.265 ;
        RECT 2656.310 906.250 2656.690 906.260 ;
        RECT 2704.405 906.250 2704.735 906.265 ;
        RECT 1473.230 905.950 1545.535 906.250 ;
        RECT 1289.190 904.890 1289.570 904.900 ;
        RECT 1473.230 904.890 1473.530 905.950 ;
        RECT 1545.205 905.935 1545.535 905.950 ;
        RECT 1670.110 905.950 1718.035 906.250 ;
        RECT 1593.710 905.570 1594.090 905.580 ;
        RECT 1670.110 905.570 1670.410 905.950 ;
        RECT 1717.705 905.935 1718.035 905.950 ;
        RECT 1862.390 905.950 1863.395 906.250 ;
        RECT 1289.190 904.590 1473.530 904.890 ;
        RECT 1569.830 905.270 1594.090 905.570 ;
        RECT 1289.190 904.580 1289.570 904.590 ;
        RECT 1545.205 904.210 1545.535 904.225 ;
        RECT 1569.830 904.210 1570.130 905.270 ;
        RECT 1593.710 905.260 1594.090 905.270 ;
        RECT 1659.070 905.270 1670.410 905.570 ;
        RECT 1717.910 905.570 1718.290 905.580 ;
        RECT 1717.910 905.270 1801.970 905.570 ;
        RECT 1659.070 904.890 1659.370 905.270 ;
        RECT 1717.910 905.260 1718.290 905.270 ;
        RECT 1618.590 904.590 1659.370 904.890 ;
        RECT 1801.670 904.890 1801.970 905.270 ;
        RECT 1808.070 904.890 1808.450 904.900 ;
        RECT 1801.670 904.590 1808.450 904.890 ;
        RECT 1545.205 903.910 1570.130 904.210 ;
        RECT 1593.710 904.210 1594.090 904.220 ;
        RECT 1618.590 904.210 1618.890 904.590 ;
        RECT 1808.070 904.580 1808.450 904.590 ;
        RECT 1855.705 904.890 1856.035 904.905 ;
        RECT 1862.390 904.890 1862.690 905.950 ;
        RECT 1863.065 905.935 1863.395 905.950 ;
        RECT 2282.830 905.950 2318.090 906.250 ;
        RECT 2172.645 905.570 2172.975 905.585 ;
        RECT 1946.110 905.270 1994.250 905.570 ;
        RECT 1855.705 904.590 1862.690 904.890 ;
        RECT 1910.905 904.890 1911.235 904.905 ;
        RECT 1946.110 904.890 1946.410 905.270 ;
        RECT 1910.905 904.590 1946.410 904.890 ;
        RECT 1855.705 904.575 1856.035 904.590 ;
        RECT 1910.905 904.575 1911.235 904.590 ;
        RECT 1593.710 903.910 1618.890 904.210 ;
        RECT 1993.950 904.210 1994.250 905.270 ;
        RECT 2172.645 905.270 2187.450 905.570 ;
        RECT 2172.645 905.255 2172.975 905.270 ;
        RECT 2042.710 904.590 2089.930 904.890 ;
        RECT 2042.710 904.210 2043.010 904.590 ;
        RECT 1993.950 903.910 2043.010 904.210 ;
        RECT 2089.630 904.210 2089.930 904.590 ;
        RECT 2125.265 904.210 2125.595 904.225 ;
        RECT 2089.630 903.910 2125.595 904.210 ;
        RECT 2187.150 904.210 2187.450 905.270 ;
        RECT 2282.830 904.890 2283.130 905.950 ;
        RECT 2317.790 905.580 2318.090 905.950 ;
        RECT 2463.150 905.950 2511.290 906.250 ;
        RECT 2317.750 905.260 2318.130 905.580 ;
        RECT 2379.645 904.890 2379.975 904.905 ;
        RECT 2235.910 904.590 2283.130 904.890 ;
        RECT 2332.510 904.590 2379.975 904.890 ;
        RECT 2235.910 904.210 2236.210 904.590 ;
        RECT 2187.150 903.910 2236.210 904.210 ;
        RECT 2317.750 904.210 2318.130 904.220 ;
        RECT 2332.510 904.210 2332.810 904.590 ;
        RECT 2379.645 904.575 2379.975 904.590 ;
        RECT 2380.565 904.890 2380.895 904.905 ;
        RECT 2463.150 904.890 2463.450 905.950 ;
        RECT 2510.990 905.580 2511.290 905.950 ;
        RECT 2656.310 905.950 2704.735 906.250 ;
        RECT 2656.310 905.940 2656.690 905.950 ;
        RECT 2704.405 905.935 2704.735 905.950 ;
        RECT 2510.950 905.260 2511.330 905.580 ;
        RECT 2916.710 905.570 2917.010 909.350 ;
        RECT 2917.600 908.900 2924.800 909.350 ;
        RECT 2863.350 905.270 2917.010 905.570 ;
        RECT 2572.845 904.890 2573.175 904.905 ;
        RECT 2380.565 904.590 2414.690 904.890 ;
        RECT 2380.565 904.575 2380.895 904.590 ;
        RECT 2317.750 903.910 2332.810 904.210 ;
        RECT 2414.390 904.210 2414.690 904.590 ;
        RECT 2429.110 904.590 2463.450 904.890 ;
        RECT 2525.710 904.590 2573.175 904.890 ;
        RECT 2429.110 904.210 2429.410 904.590 ;
        RECT 2414.390 903.910 2429.410 904.210 ;
        RECT 2510.950 904.210 2511.330 904.220 ;
        RECT 2525.710 904.210 2526.010 904.590 ;
        RECT 2572.845 904.575 2573.175 904.590 ;
        RECT 2632.185 904.890 2632.515 904.905 ;
        RECT 2656.310 904.890 2656.690 904.900 ;
        RECT 2766.505 904.890 2766.835 904.905 ;
        RECT 2632.185 904.590 2656.690 904.890 ;
        RECT 2632.185 904.575 2632.515 904.590 ;
        RECT 2656.310 904.580 2656.690 904.590 ;
        RECT 2718.910 904.590 2766.835 904.890 ;
        RECT 2608.265 904.210 2608.595 904.225 ;
        RECT 2510.950 903.910 2526.010 904.210 ;
        RECT 2607.590 903.910 2608.595 904.210 ;
        RECT 1545.205 903.895 1545.535 903.910 ;
        RECT 1593.710 903.900 1594.090 903.910 ;
        RECT 2125.265 903.895 2125.595 903.910 ;
        RECT 2317.750 903.900 2318.130 903.910 ;
        RECT 2510.950 903.900 2511.330 903.910 ;
        RECT 1808.070 903.530 1808.450 903.540 ;
        RECT 1855.705 903.530 1856.035 903.545 ;
        RECT 1808.070 903.230 1856.035 903.530 ;
        RECT 1808.070 903.220 1808.450 903.230 ;
        RECT 1855.705 903.215 1856.035 903.230 ;
        RECT 2572.845 902.850 2573.175 902.865 ;
        RECT 2607.590 902.850 2607.890 903.910 ;
        RECT 2608.265 903.895 2608.595 903.910 ;
        RECT 2704.405 904.210 2704.735 904.225 ;
        RECT 2718.910 904.210 2719.210 904.590 ;
        RECT 2766.505 904.575 2766.835 904.590 ;
        RECT 2774.785 904.890 2775.115 904.905 ;
        RECT 2774.785 904.590 2814.890 904.890 ;
        RECT 2774.785 904.575 2775.115 904.590 ;
        RECT 2704.405 903.910 2719.210 904.210 ;
        RECT 2814.590 904.210 2814.890 904.590 ;
        RECT 2863.350 904.210 2863.650 905.270 ;
        RECT 2814.590 903.910 2863.650 904.210 ;
        RECT 2704.405 903.895 2704.735 903.910 ;
        RECT 2572.845 902.550 2607.890 902.850 ;
        RECT 2572.845 902.535 2573.175 902.550 ;
      LAYER via3 ;
        RECT 1289.220 3196.180 1289.540 3196.500 ;
        RECT 1717.940 906.620 1718.260 906.940 ;
        RECT 1289.220 904.580 1289.540 904.900 ;
        RECT 1593.740 905.260 1594.060 905.580 ;
        RECT 1717.940 905.260 1718.260 905.580 ;
        RECT 1593.740 903.900 1594.060 904.220 ;
        RECT 1808.100 904.580 1808.420 904.900 ;
        RECT 2317.780 905.260 2318.100 905.580 ;
        RECT 2317.780 903.900 2318.100 904.220 ;
        RECT 2656.340 905.940 2656.660 906.260 ;
        RECT 2510.980 905.260 2511.300 905.580 ;
        RECT 2510.980 903.900 2511.300 904.220 ;
        RECT 2656.340 904.580 2656.660 904.900 ;
        RECT 1808.100 903.220 1808.420 903.540 ;
      LAYER met4 ;
        RECT 1289.215 3196.175 1289.545 3196.505 ;
        RECT 1289.230 904.905 1289.530 3196.175 ;
        RECT 1717.935 906.615 1718.265 906.945 ;
        RECT 1717.950 905.585 1718.250 906.615 ;
        RECT 2656.335 905.935 2656.665 906.265 ;
        RECT 1593.735 905.255 1594.065 905.585 ;
        RECT 1717.935 905.255 1718.265 905.585 ;
        RECT 2317.775 905.255 2318.105 905.585 ;
        RECT 2510.975 905.255 2511.305 905.585 ;
        RECT 1289.215 904.575 1289.545 904.905 ;
        RECT 1593.750 904.225 1594.050 905.255 ;
        RECT 1808.095 904.575 1808.425 904.905 ;
        RECT 1593.735 903.895 1594.065 904.225 ;
        RECT 1808.110 903.545 1808.410 904.575 ;
        RECT 2317.790 904.225 2318.090 905.255 ;
        RECT 2510.990 904.225 2511.290 905.255 ;
        RECT 2656.350 904.905 2656.650 905.935 ;
        RECT 2656.335 904.575 2656.665 904.905 ;
        RECT 2317.775 903.895 2318.105 904.225 ;
        RECT 2510.975 903.895 2511.305 904.225 ;
        RECT 1808.095 903.215 1808.425 903.545 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1325.790 3203.720 1326.110 3203.780 ;
        RECT 2901.750 3203.720 2902.070 3203.780 ;
        RECT 1325.790 3203.580 2902.070 3203.720 ;
        RECT 1325.790 3203.520 1326.110 3203.580 ;
        RECT 2901.750 3203.520 2902.070 3203.580 ;
      LAYER via ;
        RECT 1325.820 3203.520 1326.080 3203.780 ;
        RECT 2901.780 3203.520 2902.040 3203.780 ;
      LAYER met2 ;
        RECT 1325.820 3203.490 1326.080 3203.810 ;
        RECT 2901.780 3203.490 2902.040 3203.810 ;
        RECT 1325.880 3200.000 1326.020 3203.490 ;
        RECT 1325.740 3196.000 1326.020 3200.000 ;
        RECT 2901.840 1144.285 2901.980 3203.490 ;
        RECT 2901.770 1143.915 2902.050 1144.285 ;
      LAYER via2 ;
        RECT 2901.770 1143.960 2902.050 1144.240 ;
      LAYER met3 ;
        RECT 2901.745 1144.250 2902.075 1144.265 ;
        RECT 2917.600 1144.250 2924.800 1144.700 ;
        RECT 2901.745 1143.950 2924.800 1144.250 ;
        RECT 2901.745 1143.935 2902.075 1143.950 ;
        RECT 2917.600 1143.500 2924.800 1143.950 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2728.330 1374.860 2728.650 1374.920 ;
        RECT 2752.710 1374.860 2753.030 1374.920 ;
        RECT 2728.330 1374.720 2753.030 1374.860 ;
        RECT 2728.330 1374.660 2728.650 1374.720 ;
        RECT 2752.710 1374.660 2753.030 1374.720 ;
      LAYER via ;
        RECT 2728.360 1374.660 2728.620 1374.920 ;
        RECT 2752.740 1374.660 2753.000 1374.920 ;
      LAYER met2 ;
        RECT 1365.300 3196.410 1365.580 3200.000 ;
        RECT 1365.830 3196.410 1366.110 3196.525 ;
        RECT 1365.300 3196.270 1366.110 3196.410 ;
        RECT 1365.300 3196.000 1365.580 3196.270 ;
        RECT 1365.830 3196.155 1366.110 3196.270 ;
        RECT 2728.360 1374.805 2728.620 1374.950 ;
        RECT 2752.740 1374.805 2753.000 1374.950 ;
        RECT 2728.350 1374.435 2728.630 1374.805 ;
        RECT 2752.730 1374.435 2753.010 1374.805 ;
        RECT 2815.290 1374.435 2815.570 1374.805 ;
        RECT 2815.360 1372.765 2815.500 1374.435 ;
        RECT 2863.130 1374.010 2863.410 1374.125 ;
        RECT 2863.130 1373.870 2863.800 1374.010 ;
        RECT 2863.130 1373.755 2863.410 1373.870 ;
        RECT 2863.660 1373.445 2863.800 1373.870 ;
        RECT 2863.590 1373.075 2863.870 1373.445 ;
        RECT 2815.290 1372.395 2815.570 1372.765 ;
      LAYER via2 ;
        RECT 1365.830 3196.200 1366.110 3196.480 ;
        RECT 2728.350 1374.480 2728.630 1374.760 ;
        RECT 2752.730 1374.480 2753.010 1374.760 ;
        RECT 2815.290 1374.480 2815.570 1374.760 ;
        RECT 2863.130 1373.800 2863.410 1374.080 ;
        RECT 2863.590 1373.120 2863.870 1373.400 ;
        RECT 2815.290 1372.440 2815.570 1372.720 ;
      LAYER met3 ;
        RECT 1365.805 3196.500 1366.135 3196.505 ;
        RECT 1365.550 3196.490 1366.135 3196.500 ;
        RECT 1365.350 3196.190 1366.135 3196.490 ;
        RECT 1365.550 3196.180 1366.135 3196.190 ;
        RECT 1365.805 3196.175 1366.135 3196.180 ;
        RECT 2625.950 3192.410 2626.330 3192.420 ;
        RECT 2645.270 3192.410 2645.650 3192.420 ;
        RECT 2625.950 3192.110 2645.650 3192.410 ;
        RECT 2625.950 3192.100 2626.330 3192.110 ;
        RECT 2645.270 3192.100 2645.650 3192.110 ;
        RECT 1365.550 3190.370 1365.930 3190.380 ;
        RECT 2625.950 3190.370 2626.330 3190.380 ;
        RECT 1365.550 3190.070 2626.330 3190.370 ;
        RECT 1365.550 3190.060 1365.930 3190.070 ;
        RECT 2625.950 3190.060 2626.330 3190.070 ;
        RECT 2917.600 1378.850 2924.800 1379.300 ;
        RECT 2916.710 1378.550 2924.800 1378.850 ;
        RECT 2728.325 1374.770 2728.655 1374.785 ;
        RECT 2670.150 1374.470 2728.655 1374.770 ;
        RECT 2645.270 1373.410 2645.650 1373.420 ;
        RECT 2670.150 1373.410 2670.450 1374.470 ;
        RECT 2728.325 1374.455 2728.655 1374.470 ;
        RECT 2752.705 1374.770 2753.035 1374.785 ;
        RECT 2815.265 1374.770 2815.595 1374.785 ;
        RECT 2752.705 1374.470 2815.595 1374.770 ;
        RECT 2752.705 1374.455 2753.035 1374.470 ;
        RECT 2815.265 1374.455 2815.595 1374.470 ;
        RECT 2863.105 1374.090 2863.435 1374.105 ;
        RECT 2849.550 1373.790 2863.435 1374.090 ;
        RECT 2849.550 1373.410 2849.850 1373.790 ;
        RECT 2863.105 1373.775 2863.435 1373.790 ;
        RECT 2645.270 1373.110 2670.450 1373.410 ;
        RECT 2816.430 1373.110 2849.850 1373.410 ;
        RECT 2863.565 1373.410 2863.895 1373.425 ;
        RECT 2916.710 1373.410 2917.010 1378.550 ;
        RECT 2917.600 1378.100 2924.800 1378.550 ;
        RECT 2863.565 1373.110 2917.010 1373.410 ;
        RECT 2645.270 1373.100 2645.650 1373.110 ;
        RECT 2815.265 1372.730 2815.595 1372.745 ;
        RECT 2816.430 1372.730 2816.730 1373.110 ;
        RECT 2863.565 1373.095 2863.895 1373.110 ;
        RECT 2815.265 1372.430 2816.730 1372.730 ;
        RECT 2815.265 1372.415 2815.595 1372.430 ;
      LAYER via3 ;
        RECT 1365.580 3196.180 1365.900 3196.500 ;
        RECT 2625.980 3192.100 2626.300 3192.420 ;
        RECT 2645.300 3192.100 2645.620 3192.420 ;
        RECT 1365.580 3190.060 1365.900 3190.380 ;
        RECT 2625.980 3190.060 2626.300 3190.380 ;
        RECT 2645.300 1373.100 2645.620 1373.420 ;
      LAYER met4 ;
        RECT 1365.575 3196.175 1365.905 3196.505 ;
        RECT 1365.590 3190.385 1365.890 3196.175 ;
        RECT 2625.975 3192.095 2626.305 3192.425 ;
        RECT 2645.295 3192.095 2645.625 3192.425 ;
        RECT 2625.990 3190.385 2626.290 3192.095 ;
        RECT 1365.575 3190.055 1365.905 3190.385 ;
        RECT 2625.975 3190.055 2626.305 3190.385 ;
        RECT 2645.310 1373.425 2645.610 3192.095 ;
        RECT 2645.295 1373.095 2645.625 1373.425 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2653.350 1614.560 2653.670 1614.620 ;
        RECT 2898.070 1614.560 2898.390 1614.620 ;
        RECT 2653.350 1614.420 2898.390 1614.560 ;
        RECT 2653.350 1614.360 2653.670 1614.420 ;
        RECT 2898.070 1614.360 2898.390 1614.420 ;
      LAYER via ;
        RECT 2653.380 1614.360 2653.640 1614.620 ;
        RECT 2898.100 1614.360 2898.360 1614.620 ;
      LAYER met2 ;
        RECT 1404.860 3196.410 1405.140 3200.000 ;
        RECT 1405.850 3196.410 1406.130 3196.525 ;
        RECT 1404.860 3196.270 1406.130 3196.410 ;
        RECT 1404.860 3196.000 1405.140 3196.270 ;
        RECT 1405.850 3196.155 1406.130 3196.270 ;
        RECT 2653.370 3189.355 2653.650 3189.725 ;
        RECT 2653.440 1614.650 2653.580 3189.355 ;
        RECT 2653.380 1614.330 2653.640 1614.650 ;
        RECT 2898.100 1614.330 2898.360 1614.650 ;
        RECT 2898.160 1613.485 2898.300 1614.330 ;
        RECT 2898.090 1613.115 2898.370 1613.485 ;
      LAYER via2 ;
        RECT 1405.850 3196.200 1406.130 3196.480 ;
        RECT 2653.370 3189.400 2653.650 3189.680 ;
        RECT 2898.090 1613.160 2898.370 1613.440 ;
      LAYER met3 ;
        RECT 1405.825 3196.500 1406.155 3196.505 ;
        RECT 1405.825 3196.490 1406.410 3196.500 ;
        RECT 1405.825 3196.190 1406.610 3196.490 ;
        RECT 1405.825 3196.180 1406.410 3196.190 ;
        RECT 1405.825 3196.175 1406.155 3196.180 ;
        RECT 1406.030 3189.690 1406.410 3189.700 ;
        RECT 2653.345 3189.690 2653.675 3189.705 ;
        RECT 1406.030 3189.390 2653.675 3189.690 ;
        RECT 1406.030 3189.380 1406.410 3189.390 ;
        RECT 2653.345 3189.375 2653.675 3189.390 ;
        RECT 2898.065 1613.450 2898.395 1613.465 ;
        RECT 2917.600 1613.450 2924.800 1613.900 ;
        RECT 2898.065 1613.150 2924.800 1613.450 ;
        RECT 2898.065 1613.135 2898.395 1613.150 ;
        RECT 2917.600 1612.700 2924.800 1613.150 ;
      LAYER via3 ;
        RECT 1406.060 3196.180 1406.380 3196.500 ;
        RECT 1406.060 3189.380 1406.380 3189.700 ;
      LAYER met4 ;
        RECT 1406.055 3196.175 1406.385 3196.505 ;
        RECT 1406.070 3189.705 1406.370 3196.175 ;
        RECT 1406.055 3189.375 1406.385 3189.705 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1444.490 3209.755 1444.770 3210.125 ;
        RECT 1444.560 3200.000 1444.700 3209.755 ;
        RECT 1444.420 3196.000 1444.700 3200.000 ;
      LAYER via2 ;
        RECT 1444.490 3209.800 1444.770 3210.080 ;
      LAYER met3 ;
        RECT 1444.465 3210.090 1444.795 3210.105 ;
        RECT 2639.750 3210.090 2640.130 3210.100 ;
        RECT 1444.465 3209.790 2640.130 3210.090 ;
        RECT 1444.465 3209.775 1444.795 3209.790 ;
        RECT 2639.750 3209.780 2640.130 3209.790 ;
        RECT 2637.910 2573.980 2638.290 2574.300 ;
        RECT 2637.950 2573.620 2638.250 2573.980 ;
        RECT 2637.910 2573.300 2638.290 2573.620 ;
        RECT 2637.910 2561.370 2638.290 2561.380 ;
        RECT 2637.910 2561.070 2639.170 2561.370 ;
        RECT 2637.910 2561.060 2638.290 2561.070 ;
        RECT 2638.870 2560.700 2639.170 2561.070 ;
        RECT 2638.830 2560.380 2639.210 2560.700 ;
        RECT 2638.830 2526.010 2639.210 2526.020 ;
        RECT 2637.030 2525.710 2639.210 2526.010 ;
        RECT 2637.030 2524.660 2637.330 2525.710 ;
        RECT 2638.830 2525.700 2639.210 2525.710 ;
        RECT 2636.990 2524.340 2637.370 2524.660 ;
        RECT 2638.830 2462.460 2639.210 2462.780 ;
        RECT 2638.870 2462.090 2639.170 2462.460 ;
        RECT 2640.670 2462.090 2641.050 2462.100 ;
        RECT 2638.870 2461.790 2641.050 2462.090 ;
        RECT 2640.670 2461.780 2641.050 2461.790 ;
        RECT 2637.910 2415.170 2638.290 2415.180 ;
        RECT 2640.670 2415.170 2641.050 2415.180 ;
        RECT 2637.910 2414.870 2641.050 2415.170 ;
        RECT 2637.910 2414.860 2638.290 2414.870 ;
        RECT 2640.670 2414.860 2641.050 2414.870 ;
        RECT 2637.910 2359.100 2638.290 2359.420 ;
        RECT 2637.950 2358.730 2638.250 2359.100 ;
        RECT 2639.750 2358.730 2640.130 2358.740 ;
        RECT 2637.950 2358.430 2640.130 2358.730 ;
        RECT 2639.750 2358.420 2640.130 2358.430 ;
        RECT 2639.750 2311.810 2640.130 2311.820 ;
        RECT 2640.670 2311.810 2641.050 2311.820 ;
        RECT 2639.750 2311.510 2641.050 2311.810 ;
        RECT 2639.750 2311.500 2640.130 2311.510 ;
        RECT 2640.670 2311.500 2641.050 2311.510 ;
        RECT 2638.830 2270.330 2639.210 2270.340 ;
        RECT 2640.670 2270.330 2641.050 2270.340 ;
        RECT 2638.830 2270.030 2641.050 2270.330 ;
        RECT 2638.830 2270.020 2639.210 2270.030 ;
        RECT 2640.670 2270.020 2641.050 2270.030 ;
        RECT 2638.830 2236.330 2639.210 2236.340 ;
        RECT 2637.950 2236.030 2639.210 2236.330 ;
        RECT 2637.950 2234.980 2638.250 2236.030 ;
        RECT 2638.830 2236.020 2639.210 2236.030 ;
        RECT 2637.910 2234.660 2638.290 2234.980 ;
        RECT 2637.910 2125.490 2638.290 2125.500 ;
        RECT 2635.190 2125.190 2638.290 2125.490 ;
        RECT 2635.190 2124.810 2635.490 2125.190 ;
        RECT 2637.910 2125.180 2638.290 2125.190 ;
        RECT 2637.910 2124.810 2638.290 2124.820 ;
        RECT 2635.190 2124.510 2638.290 2124.810 ;
        RECT 2637.910 2124.500 2638.290 2124.510 ;
        RECT 2917.600 1848.050 2924.800 1848.500 ;
        RECT 2916.710 1847.750 2924.800 1848.050 ;
        RECT 2637.910 1843.970 2638.290 1843.980 ;
        RECT 2637.910 1843.670 2642.850 1843.970 ;
        RECT 2637.910 1843.660 2638.290 1843.670 ;
        RECT 2642.550 1843.290 2642.850 1843.670 ;
        RECT 2691.310 1843.670 2739.450 1843.970 ;
        RECT 2642.550 1842.990 2690.690 1843.290 ;
        RECT 2690.390 1842.610 2690.690 1842.990 ;
        RECT 2691.310 1842.610 2691.610 1843.670 ;
        RECT 2739.150 1843.290 2739.450 1843.670 ;
        RECT 2787.910 1843.670 2836.050 1843.970 ;
        RECT 2739.150 1842.990 2787.290 1843.290 ;
        RECT 2690.390 1842.310 2691.610 1842.610 ;
        RECT 2786.990 1842.610 2787.290 1842.990 ;
        RECT 2787.910 1842.610 2788.210 1843.670 ;
        RECT 2835.750 1843.290 2836.050 1843.670 ;
        RECT 2916.710 1843.290 2917.010 1847.750 ;
        RECT 2917.600 1847.300 2924.800 1847.750 ;
        RECT 2835.750 1842.990 2883.890 1843.290 ;
        RECT 2786.990 1842.310 2788.210 1842.610 ;
        RECT 2883.590 1842.610 2883.890 1842.990 ;
        RECT 2884.510 1842.990 2917.010 1843.290 ;
        RECT 2884.510 1842.610 2884.810 1842.990 ;
        RECT 2883.590 1842.310 2884.810 1842.610 ;
      LAYER via3 ;
        RECT 2639.780 3209.780 2640.100 3210.100 ;
        RECT 2637.940 2573.980 2638.260 2574.300 ;
        RECT 2637.940 2573.300 2638.260 2573.620 ;
        RECT 2637.940 2561.060 2638.260 2561.380 ;
        RECT 2638.860 2560.380 2639.180 2560.700 ;
        RECT 2638.860 2525.700 2639.180 2526.020 ;
        RECT 2637.020 2524.340 2637.340 2524.660 ;
        RECT 2638.860 2462.460 2639.180 2462.780 ;
        RECT 2640.700 2461.780 2641.020 2462.100 ;
        RECT 2637.940 2414.860 2638.260 2415.180 ;
        RECT 2640.700 2414.860 2641.020 2415.180 ;
        RECT 2637.940 2359.100 2638.260 2359.420 ;
        RECT 2639.780 2358.420 2640.100 2358.740 ;
        RECT 2639.780 2311.500 2640.100 2311.820 ;
        RECT 2640.700 2311.500 2641.020 2311.820 ;
        RECT 2638.860 2270.020 2639.180 2270.340 ;
        RECT 2640.700 2270.020 2641.020 2270.340 ;
        RECT 2638.860 2236.020 2639.180 2236.340 ;
        RECT 2637.940 2234.660 2638.260 2234.980 ;
        RECT 2637.940 2125.180 2638.260 2125.500 ;
        RECT 2637.940 2124.500 2638.260 2124.820 ;
        RECT 2637.940 1843.660 2638.260 1843.980 ;
      LAYER met4 ;
        RECT 2639.775 3209.775 2640.105 3210.105 ;
        RECT 2639.790 3058.890 2640.090 3209.775 ;
        RECT 2639.350 3057.710 2640.530 3058.890 ;
        RECT 2639.350 3054.310 2640.530 3055.490 ;
        RECT 2639.790 2769.450 2640.090 3054.310 ;
        RECT 2637.950 2769.150 2640.090 2769.450 ;
        RECT 2637.950 2766.050 2638.250 2769.150 ;
        RECT 2637.950 2765.750 2640.090 2766.050 ;
        RECT 2639.790 2671.290 2640.090 2765.750 ;
        RECT 2639.350 2670.110 2640.530 2671.290 ;
        RECT 2637.510 2666.710 2638.690 2667.890 ;
        RECT 2637.950 2574.305 2638.250 2666.710 ;
        RECT 2637.935 2573.975 2638.265 2574.305 ;
        RECT 2637.935 2573.295 2638.265 2573.625 ;
        RECT 2637.950 2561.385 2638.250 2573.295 ;
        RECT 2637.935 2561.055 2638.265 2561.385 ;
        RECT 2638.855 2560.375 2639.185 2560.705 ;
        RECT 2638.870 2526.025 2639.170 2560.375 ;
        RECT 2638.855 2525.695 2639.185 2526.025 ;
        RECT 2637.015 2524.335 2637.345 2524.665 ;
        RECT 2637.030 2477.050 2637.330 2524.335 ;
        RECT 2637.030 2476.750 2639.170 2477.050 ;
        RECT 2638.870 2462.785 2639.170 2476.750 ;
        RECT 2638.855 2462.455 2639.185 2462.785 ;
        RECT 2640.695 2461.775 2641.025 2462.105 ;
        RECT 2640.710 2415.185 2641.010 2461.775 ;
        RECT 2637.935 2414.855 2638.265 2415.185 ;
        RECT 2640.695 2414.855 2641.025 2415.185 ;
        RECT 2637.950 2359.425 2638.250 2414.855 ;
        RECT 2637.935 2359.095 2638.265 2359.425 ;
        RECT 2639.775 2358.415 2640.105 2358.745 ;
        RECT 2639.790 2311.825 2640.090 2358.415 ;
        RECT 2639.775 2311.495 2640.105 2311.825 ;
        RECT 2640.695 2311.495 2641.025 2311.825 ;
        RECT 2640.710 2270.345 2641.010 2311.495 ;
        RECT 2638.855 2270.015 2639.185 2270.345 ;
        RECT 2640.695 2270.015 2641.025 2270.345 ;
        RECT 2638.870 2236.345 2639.170 2270.015 ;
        RECT 2638.855 2236.015 2639.185 2236.345 ;
        RECT 2637.935 2234.655 2638.265 2234.985 ;
        RECT 2637.950 2125.505 2638.250 2234.655 ;
        RECT 2637.935 2125.175 2638.265 2125.505 ;
        RECT 2637.935 2124.495 2638.265 2124.825 ;
        RECT 2637.950 1947.090 2638.250 2124.495 ;
        RECT 2637.510 1945.910 2638.690 1947.090 ;
        RECT 2637.510 1942.510 2638.690 1943.690 ;
        RECT 2637.950 1843.985 2638.250 1942.510 ;
        RECT 2637.935 1843.655 2638.265 1843.985 ;
      LAYER met5 ;
        RECT 2630.860 3057.500 2640.740 3059.100 ;
        RECT 2630.860 3055.700 2632.460 3057.500 ;
        RECT 2630.860 3054.100 2640.740 3055.700 ;
        RECT 2629.940 2669.900 2640.740 2671.500 ;
        RECT 2629.940 2668.100 2631.540 2669.900 ;
        RECT 2629.940 2666.500 2638.900 2668.100 ;
        RECT 2629.940 1945.700 2638.900 1947.300 ;
        RECT 2629.940 1943.900 2631.540 1945.700 ;
        RECT 2629.940 1942.300 2638.900 1943.900 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1484.030 3214.260 1484.350 3214.320 ;
        RECT 2653.810 3214.260 2654.130 3214.320 ;
        RECT 1484.030 3214.120 2654.130 3214.260 ;
        RECT 1484.030 3214.060 1484.350 3214.120 ;
        RECT 2653.810 3214.060 2654.130 3214.120 ;
        RECT 2653.810 2083.760 2654.130 2083.820 ;
        RECT 2900.830 2083.760 2901.150 2083.820 ;
        RECT 2653.810 2083.620 2901.150 2083.760 ;
        RECT 2653.810 2083.560 2654.130 2083.620 ;
        RECT 2900.830 2083.560 2901.150 2083.620 ;
      LAYER via ;
        RECT 1484.060 3214.060 1484.320 3214.320 ;
        RECT 2653.840 3214.060 2654.100 3214.320 ;
        RECT 2653.840 2083.560 2654.100 2083.820 ;
        RECT 2900.860 2083.560 2901.120 2083.820 ;
      LAYER met2 ;
        RECT 1484.060 3214.030 1484.320 3214.350 ;
        RECT 2653.840 3214.030 2654.100 3214.350 ;
        RECT 1484.120 3200.000 1484.260 3214.030 ;
        RECT 1483.980 3196.000 1484.260 3200.000 ;
        RECT 2653.900 2083.850 2654.040 3214.030 ;
        RECT 2653.840 2083.530 2654.100 2083.850 ;
        RECT 2900.860 2083.530 2901.120 2083.850 ;
        RECT 2900.920 2082.685 2901.060 2083.530 ;
        RECT 2900.850 2082.315 2901.130 2082.685 ;
      LAYER via2 ;
        RECT 2900.850 2082.360 2901.130 2082.640 ;
      LAYER met3 ;
        RECT 2900.825 2082.650 2901.155 2082.665 ;
        RECT 2917.600 2082.650 2924.800 2083.100 ;
        RECT 2900.825 2082.350 2924.800 2082.650 ;
        RECT 2900.825 2082.335 2901.155 2082.350 ;
        RECT 2917.600 2081.900 2924.800 2082.350 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2654.730 2318.360 2655.050 2318.420 ;
        RECT 2898.990 2318.360 2899.310 2318.420 ;
        RECT 2654.730 2318.220 2899.310 2318.360 ;
        RECT 2654.730 2318.160 2655.050 2318.220 ;
        RECT 2898.990 2318.160 2899.310 2318.220 ;
      LAYER via ;
        RECT 2654.760 2318.160 2655.020 2318.420 ;
        RECT 2899.020 2318.160 2899.280 2318.420 ;
      LAYER met2 ;
        RECT 1523.080 3196.410 1523.360 3200.000 ;
        RECT 1524.530 3196.410 1524.810 3196.525 ;
        RECT 1523.080 3196.270 1524.810 3196.410 ;
        RECT 1523.080 3196.000 1523.360 3196.270 ;
        RECT 1524.530 3196.155 1524.810 3196.270 ;
        RECT 2654.750 3191.395 2655.030 3191.765 ;
        RECT 2654.820 2318.450 2654.960 3191.395 ;
        RECT 2654.760 2318.130 2655.020 2318.450 ;
        RECT 2899.020 2318.130 2899.280 2318.450 ;
        RECT 2899.080 2317.285 2899.220 2318.130 ;
        RECT 2899.010 2316.915 2899.290 2317.285 ;
      LAYER via2 ;
        RECT 1524.530 3196.200 1524.810 3196.480 ;
        RECT 2654.750 3191.440 2655.030 3191.720 ;
        RECT 2899.010 2316.960 2899.290 2317.240 ;
      LAYER met3 ;
        RECT 1524.505 3196.490 1524.835 3196.505 ;
        RECT 1537.590 3196.490 1537.970 3196.500 ;
        RECT 1524.505 3196.190 1537.970 3196.490 ;
        RECT 1524.505 3196.175 1524.835 3196.190 ;
        RECT 1537.590 3196.180 1537.970 3196.190 ;
        RECT 2627.790 3191.730 2628.170 3191.740 ;
        RECT 2654.725 3191.730 2655.055 3191.745 ;
        RECT 2627.790 3191.430 2655.055 3191.730 ;
        RECT 2627.790 3191.420 2628.170 3191.430 ;
        RECT 2654.725 3191.415 2655.055 3191.430 ;
        RECT 1537.590 3189.010 1537.970 3189.020 ;
        RECT 2627.790 3189.010 2628.170 3189.020 ;
        RECT 1537.590 3188.710 2628.170 3189.010 ;
        RECT 1537.590 3188.700 1537.970 3188.710 ;
        RECT 2627.790 3188.700 2628.170 3188.710 ;
        RECT 2898.985 2317.250 2899.315 2317.265 ;
        RECT 2917.600 2317.250 2924.800 2317.700 ;
        RECT 2898.985 2316.950 2924.800 2317.250 ;
        RECT 2898.985 2316.935 2899.315 2316.950 ;
        RECT 2917.600 2316.500 2924.800 2316.950 ;
      LAYER via3 ;
        RECT 1537.620 3196.180 1537.940 3196.500 ;
        RECT 2627.820 3191.420 2628.140 3191.740 ;
        RECT 1537.620 3188.700 1537.940 3189.020 ;
        RECT 2627.820 3188.700 2628.140 3189.020 ;
      LAYER met4 ;
        RECT 1537.615 3196.175 1537.945 3196.505 ;
        RECT 1537.630 3189.025 1537.930 3196.175 ;
        RECT 2627.815 3191.415 2628.145 3191.745 ;
        RECT 2627.830 3189.025 2628.130 3191.415 ;
        RECT 1537.615 3188.695 1537.945 3189.025 ;
        RECT 2627.815 3188.695 2628.145 3189.025 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1393.870 146.100 1394.190 146.160 ;
        RECT 1415.490 146.100 1415.810 146.160 ;
        RECT 1393.870 145.960 1415.810 146.100 ;
        RECT 1393.870 145.900 1394.190 145.960 ;
        RECT 1415.490 145.900 1415.810 145.960 ;
        RECT 2331.350 146.100 2331.670 146.160 ;
        RECT 2366.310 146.100 2366.630 146.160 ;
        RECT 2331.350 145.960 2366.630 146.100 ;
        RECT 2331.350 145.900 2331.670 145.960 ;
        RECT 2366.310 145.900 2366.630 145.960 ;
        RECT 2863.110 146.100 2863.430 146.160 ;
        RECT 2883.810 146.100 2884.130 146.160 ;
        RECT 2863.110 145.960 2884.130 146.100 ;
        RECT 2863.110 145.900 2863.430 145.960 ;
        RECT 2883.810 145.900 2884.130 145.960 ;
        RECT 2608.270 145.420 2608.590 145.480 ;
        RECT 2629.430 145.420 2629.750 145.480 ;
        RECT 2608.270 145.280 2629.750 145.420 ;
        RECT 2608.270 145.220 2608.590 145.280 ;
        RECT 2629.430 145.220 2629.750 145.280 ;
      LAYER via ;
        RECT 1393.900 145.900 1394.160 146.160 ;
        RECT 1415.520 145.900 1415.780 146.160 ;
        RECT 2331.380 145.900 2331.640 146.160 ;
        RECT 2366.340 145.900 2366.600 146.160 ;
        RECT 2863.140 145.900 2863.400 146.160 ;
        RECT 2883.840 145.900 2884.100 146.160 ;
        RECT 2608.300 145.220 2608.560 145.480 ;
        RECT 2629.460 145.220 2629.720 145.480 ;
      LAYER met2 ;
        RECT 1181.300 3196.410 1181.580 3200.000 ;
        RECT 1182.750 3196.410 1183.030 3196.525 ;
        RECT 1181.300 3196.270 1183.030 3196.410 ;
        RECT 1181.300 3196.000 1181.580 3196.270 ;
        RECT 1182.750 3196.155 1183.030 3196.270 ;
        RECT 1917.830 147.715 1918.110 148.085 ;
        RECT 2801.030 147.715 2801.310 148.085 ;
        RECT 1586.630 147.035 1586.910 147.405 ;
        RECT 1593.530 147.035 1593.810 147.405 ;
        RECT 1754.990 147.035 1755.270 147.405 ;
        RECT 1466.110 146.355 1466.390 146.725 ;
        RECT 1393.900 146.045 1394.160 146.190 ;
        RECT 1415.520 146.045 1415.780 146.190 ;
        RECT 1370.430 145.930 1370.710 146.045 ;
        RECT 1371.350 145.930 1371.630 146.045 ;
        RECT 1370.430 145.790 1371.630 145.930 ;
        RECT 1370.430 145.675 1370.710 145.790 ;
        RECT 1371.350 145.675 1371.630 145.790 ;
        RECT 1393.890 145.675 1394.170 146.045 ;
        RECT 1415.510 145.675 1415.790 146.045 ;
        RECT 1466.180 144.685 1466.320 146.355 ;
        RECT 1586.700 144.685 1586.840 147.035 ;
        RECT 1593.600 146.725 1593.740 147.035 ;
        RECT 1593.530 146.355 1593.810 146.725 ;
        RECT 1755.060 146.045 1755.200 147.035 ;
        RECT 1869.530 146.355 1869.810 146.725 ;
        RECT 1754.990 145.675 1755.270 146.045 ;
        RECT 1869.600 144.685 1869.740 146.355 ;
        RECT 1917.900 146.045 1918.040 147.715 ;
        RECT 2703.970 147.035 2704.250 147.405 ;
        RECT 2366.330 146.355 2366.610 146.725 ;
        RECT 2366.400 146.190 2366.540 146.355 ;
        RECT 1917.830 145.675 1918.110 146.045 ;
        RECT 1979.470 145.930 1979.750 146.045 ;
        RECT 1980.390 145.930 1980.670 146.045 ;
        RECT 1979.470 145.790 1980.670 145.930 ;
        RECT 2331.380 145.870 2331.640 146.190 ;
        RECT 2366.340 145.870 2366.600 146.190 ;
        RECT 1979.470 145.675 1979.750 145.790 ;
        RECT 1980.390 145.675 1980.670 145.790 ;
        RECT 2331.440 145.365 2331.580 145.870 ;
        RECT 2629.450 145.675 2629.730 146.045 ;
        RECT 2629.520 145.510 2629.660 145.675 ;
        RECT 2608.300 145.365 2608.560 145.510 ;
        RECT 2331.370 144.995 2331.650 145.365 ;
        RECT 2608.290 144.995 2608.570 145.365 ;
        RECT 2629.460 145.190 2629.720 145.510 ;
        RECT 2704.040 145.250 2704.180 147.035 ;
        RECT 2801.100 146.725 2801.240 147.715 ;
        RECT 2801.030 146.355 2801.310 146.725 ;
        RECT 2863.140 146.045 2863.400 146.190 ;
        RECT 2883.840 146.045 2884.100 146.190 ;
        RECT 2863.130 145.675 2863.410 146.045 ;
        RECT 2883.830 145.675 2884.110 146.045 ;
        RECT 2704.430 145.250 2704.710 145.365 ;
        RECT 2704.040 145.110 2704.710 145.250 ;
        RECT 2704.430 144.995 2704.710 145.110 ;
        RECT 1466.110 144.315 1466.390 144.685 ;
        RECT 1586.630 144.315 1586.910 144.685 ;
        RECT 1869.530 144.315 1869.810 144.685 ;
      LAYER via2 ;
        RECT 1182.750 3196.200 1183.030 3196.480 ;
        RECT 1917.830 147.760 1918.110 148.040 ;
        RECT 2801.030 147.760 2801.310 148.040 ;
        RECT 1586.630 147.080 1586.910 147.360 ;
        RECT 1593.530 147.080 1593.810 147.360 ;
        RECT 1754.990 147.080 1755.270 147.360 ;
        RECT 1466.110 146.400 1466.390 146.680 ;
        RECT 1370.430 145.720 1370.710 146.000 ;
        RECT 1371.350 145.720 1371.630 146.000 ;
        RECT 1393.890 145.720 1394.170 146.000 ;
        RECT 1415.510 145.720 1415.790 146.000 ;
        RECT 1593.530 146.400 1593.810 146.680 ;
        RECT 1869.530 146.400 1869.810 146.680 ;
        RECT 1754.990 145.720 1755.270 146.000 ;
        RECT 2703.970 147.080 2704.250 147.360 ;
        RECT 2366.330 146.400 2366.610 146.680 ;
        RECT 1917.830 145.720 1918.110 146.000 ;
        RECT 1979.470 145.720 1979.750 146.000 ;
        RECT 1980.390 145.720 1980.670 146.000 ;
        RECT 2629.450 145.720 2629.730 146.000 ;
        RECT 2331.370 145.040 2331.650 145.320 ;
        RECT 2608.290 145.040 2608.570 145.320 ;
        RECT 2801.030 146.400 2801.310 146.680 ;
        RECT 2863.130 145.720 2863.410 146.000 ;
        RECT 2883.830 145.720 2884.110 146.000 ;
        RECT 2704.430 145.040 2704.710 145.320 ;
        RECT 1466.110 144.360 1466.390 144.640 ;
        RECT 1586.630 144.360 1586.910 144.640 ;
        RECT 1869.530 144.360 1869.810 144.640 ;
      LAYER met3 ;
        RECT 1182.725 3196.490 1183.055 3196.505 ;
        RECT 1186.150 3196.490 1186.530 3196.500 ;
        RECT 1182.725 3196.190 1186.530 3196.490 ;
        RECT 1182.725 3196.175 1183.055 3196.190 ;
        RECT 1186.150 3196.180 1186.530 3196.190 ;
        RECT 1690.310 148.050 1690.690 148.060 ;
        RECT 1869.710 148.050 1870.090 148.060 ;
        RECT 1917.805 148.050 1918.135 148.065 ;
        RECT 1690.310 147.750 1725.610 148.050 ;
        RECT 1690.310 147.740 1690.690 147.750 ;
        RECT 1586.605 147.370 1586.935 147.385 ;
        RECT 1593.505 147.370 1593.835 147.385 ;
        RECT 1231.270 147.070 1280.330 147.370 ;
        RECT 1186.150 146.690 1186.530 146.700 ;
        RECT 1231.270 146.690 1231.570 147.070 ;
        RECT 1186.150 146.390 1231.570 146.690 ;
        RECT 1186.150 146.380 1186.530 146.390 ;
        RECT 1280.030 146.010 1280.330 147.070 ;
        RECT 1586.605 147.070 1593.835 147.370 ;
        RECT 1725.310 147.370 1725.610 147.750 ;
        RECT 1869.710 147.750 1918.135 148.050 ;
        RECT 1869.710 147.740 1870.090 147.750 ;
        RECT 1917.805 147.735 1918.135 147.750 ;
        RECT 2269.910 148.050 2270.290 148.060 ;
        RECT 2752.910 148.050 2753.290 148.060 ;
        RECT 2801.005 148.050 2801.335 148.065 ;
        RECT 2269.910 147.750 2318.090 148.050 ;
        RECT 2269.910 147.740 2270.290 147.750 ;
        RECT 1754.965 147.370 1755.295 147.385 ;
        RECT 2317.790 147.380 2318.090 147.750 ;
        RECT 2752.910 147.750 2801.335 148.050 ;
        RECT 2752.910 147.740 2753.290 147.750 ;
        RECT 2801.005 147.735 2801.335 147.750 ;
        RECT 1725.310 147.070 1755.295 147.370 ;
        RECT 1586.605 147.055 1586.935 147.070 ;
        RECT 1593.505 147.055 1593.835 147.070 ;
        RECT 1754.965 147.055 1755.295 147.070 ;
        RECT 2066.630 147.070 2089.930 147.370 ;
        RECT 1466.085 146.690 1466.415 146.705 ;
        RECT 1593.505 146.700 1593.835 146.705 ;
        RECT 1869.505 146.700 1869.835 146.705 ;
        RECT 1593.505 146.690 1594.090 146.700 ;
        RECT 1690.310 146.690 1690.690 146.700 ;
        RECT 1466.085 146.390 1497.450 146.690 ;
        RECT 1466.085 146.375 1466.415 146.390 ;
        RECT 1370.405 146.010 1370.735 146.025 ;
        RECT 1280.030 145.710 1370.735 146.010 ;
        RECT 1370.405 145.695 1370.735 145.710 ;
        RECT 1371.325 146.010 1371.655 146.025 ;
        RECT 1393.865 146.010 1394.195 146.025 ;
        RECT 1371.325 145.710 1394.195 146.010 ;
        RECT 1371.325 145.695 1371.655 145.710 ;
        RECT 1393.865 145.695 1394.195 145.710 ;
        RECT 1415.485 146.010 1415.815 146.025 ;
        RECT 1441.910 146.010 1442.290 146.020 ;
        RECT 1415.485 145.710 1442.290 146.010 ;
        RECT 1497.150 146.010 1497.450 146.390 ;
        RECT 1593.505 146.390 1594.470 146.690 ;
        RECT 1659.070 146.390 1690.690 146.690 ;
        RECT 1593.505 146.380 1594.090 146.390 ;
        RECT 1593.505 146.375 1593.835 146.380 ;
        RECT 1538.510 146.010 1538.890 146.020 ;
        RECT 1659.070 146.010 1659.370 146.390 ;
        RECT 1690.310 146.380 1690.690 146.390 ;
        RECT 1869.505 146.690 1870.090 146.700 ;
        RECT 1869.505 146.390 1870.470 146.690 ;
        RECT 1869.505 146.380 1870.090 146.390 ;
        RECT 1869.505 146.375 1869.835 146.380 ;
        RECT 1497.150 145.710 1538.890 146.010 ;
        RECT 1415.485 145.695 1415.815 145.710 ;
        RECT 1441.910 145.700 1442.290 145.710 ;
        RECT 1538.510 145.700 1538.890 145.710 ;
        RECT 1618.590 145.710 1659.370 146.010 ;
        RECT 1754.965 146.010 1755.295 146.025 ;
        RECT 1917.805 146.010 1918.135 146.025 ;
        RECT 1979.445 146.010 1979.775 146.025 ;
        RECT 1754.965 145.710 1779.890 146.010 ;
        RECT 1593.710 145.330 1594.090 145.340 ;
        RECT 1618.590 145.330 1618.890 145.710 ;
        RECT 1754.965 145.695 1755.295 145.710 ;
        RECT 1593.710 145.030 1618.890 145.330 ;
        RECT 1593.710 145.020 1594.090 145.030 ;
        RECT 1441.910 144.650 1442.290 144.660 ;
        RECT 1466.085 144.650 1466.415 144.665 ;
        RECT 1441.910 144.350 1466.415 144.650 ;
        RECT 1441.910 144.340 1442.290 144.350 ;
        RECT 1466.085 144.335 1466.415 144.350 ;
        RECT 1538.510 144.650 1538.890 144.660 ;
        RECT 1586.605 144.650 1586.935 144.665 ;
        RECT 1538.510 144.350 1586.935 144.650 ;
        RECT 1779.590 144.650 1779.890 145.710 ;
        RECT 1917.805 145.710 1979.775 146.010 ;
        RECT 1917.805 145.695 1918.135 145.710 ;
        RECT 1979.445 145.695 1979.775 145.710 ;
        RECT 1980.365 146.010 1980.695 146.025 ;
        RECT 2066.630 146.010 2066.930 147.070 ;
        RECT 1980.365 145.710 2066.930 146.010 ;
        RECT 2089.630 146.010 2089.930 147.070 ;
        RECT 2317.750 147.060 2318.130 147.380 ;
        RECT 2510.950 147.370 2511.330 147.380 ;
        RECT 2607.550 147.370 2607.930 147.380 ;
        RECT 2476.030 147.070 2511.330 147.370 ;
        RECT 2366.305 146.690 2366.635 146.705 ;
        RECT 2138.390 146.390 2187.450 146.690 ;
        RECT 2089.630 145.710 2092.690 146.010 ;
        RECT 1980.365 145.695 1980.695 145.710 ;
        RECT 2092.390 145.330 2092.690 145.710 ;
        RECT 2138.390 145.330 2138.690 146.390 ;
        RECT 2092.390 145.030 2138.690 145.330 ;
        RECT 2187.150 145.330 2187.450 146.390 ;
        RECT 2366.305 146.390 2380.650 146.690 ;
        RECT 2366.305 146.375 2366.635 146.390 ;
        RECT 2269.910 146.010 2270.290 146.020 ;
        RECT 2235.910 145.710 2270.290 146.010 ;
        RECT 2235.910 145.330 2236.210 145.710 ;
        RECT 2269.910 145.700 2270.290 145.710 ;
        RECT 2187.150 145.030 2236.210 145.330 ;
        RECT 2317.750 145.330 2318.130 145.340 ;
        RECT 2331.345 145.330 2331.675 145.345 ;
        RECT 2317.750 145.030 2331.675 145.330 ;
        RECT 2380.350 145.330 2380.650 146.390 ;
        RECT 2476.030 146.010 2476.330 147.070 ;
        RECT 2510.950 147.060 2511.330 147.070 ;
        RECT 2572.630 147.070 2607.930 147.370 ;
        RECT 2572.630 146.010 2572.930 147.070 ;
        RECT 2607.550 147.060 2607.930 147.070 ;
        RECT 2656.310 147.370 2656.690 147.380 ;
        RECT 2703.945 147.370 2704.275 147.385 ;
        RECT 2656.310 147.070 2704.275 147.370 ;
        RECT 2656.310 147.060 2656.690 147.070 ;
        RECT 2703.945 147.055 2704.275 147.070 ;
        RECT 2801.005 146.690 2801.335 146.705 ;
        RECT 2917.600 146.690 2924.800 147.140 ;
        RECT 2801.005 146.390 2815.810 146.690 ;
        RECT 2801.005 146.375 2801.335 146.390 ;
        RECT 2429.110 145.710 2476.330 146.010 ;
        RECT 2525.710 145.710 2572.930 146.010 ;
        RECT 2629.425 146.010 2629.755 146.025 ;
        RECT 2656.310 146.010 2656.690 146.020 ;
        RECT 2752.910 146.010 2753.290 146.020 ;
        RECT 2629.425 145.710 2656.690 146.010 ;
        RECT 2429.110 145.330 2429.410 145.710 ;
        RECT 2380.350 145.030 2429.410 145.330 ;
        RECT 2510.950 145.330 2511.330 145.340 ;
        RECT 2525.710 145.330 2526.010 145.710 ;
        RECT 2629.425 145.695 2629.755 145.710 ;
        RECT 2656.310 145.700 2656.690 145.710 ;
        RECT 2718.910 145.710 2753.290 146.010 ;
        RECT 2510.950 145.030 2526.010 145.330 ;
        RECT 2607.550 145.330 2607.930 145.340 ;
        RECT 2608.265 145.330 2608.595 145.345 ;
        RECT 2607.550 145.030 2608.595 145.330 ;
        RECT 2317.750 145.020 2318.130 145.030 ;
        RECT 2331.345 145.015 2331.675 145.030 ;
        RECT 2510.950 145.020 2511.330 145.030 ;
        RECT 2607.550 145.020 2607.930 145.030 ;
        RECT 2608.265 145.015 2608.595 145.030 ;
        RECT 2704.405 145.330 2704.735 145.345 ;
        RECT 2718.910 145.330 2719.210 145.710 ;
        RECT 2752.910 145.700 2753.290 145.710 ;
        RECT 2704.405 145.030 2719.210 145.330 ;
        RECT 2815.510 145.330 2815.810 146.390 ;
        RECT 2916.710 146.390 2924.800 146.690 ;
        RECT 2863.105 146.010 2863.435 146.025 ;
        RECT 2849.550 145.710 2863.435 146.010 ;
        RECT 2849.550 145.330 2849.850 145.710 ;
        RECT 2863.105 145.695 2863.435 145.710 ;
        RECT 2883.805 146.010 2884.135 146.025 ;
        RECT 2916.710 146.010 2917.010 146.390 ;
        RECT 2883.805 145.710 2917.010 146.010 ;
        RECT 2917.600 145.940 2924.800 146.390 ;
        RECT 2883.805 145.695 2884.135 145.710 ;
        RECT 2815.510 145.030 2849.850 145.330 ;
        RECT 2704.405 145.015 2704.735 145.030 ;
        RECT 1820.990 144.650 1822.210 144.820 ;
        RECT 1869.505 144.650 1869.835 144.665 ;
        RECT 1779.590 144.520 1869.835 144.650 ;
        RECT 1779.590 144.350 1821.290 144.520 ;
        RECT 1821.910 144.350 1869.835 144.520 ;
        RECT 1538.510 144.340 1538.890 144.350 ;
        RECT 1586.605 144.335 1586.935 144.350 ;
        RECT 1869.505 144.335 1869.835 144.350 ;
      LAYER via3 ;
        RECT 1186.180 3196.180 1186.500 3196.500 ;
        RECT 1690.340 147.740 1690.660 148.060 ;
        RECT 1186.180 146.380 1186.500 146.700 ;
        RECT 1869.740 147.740 1870.060 148.060 ;
        RECT 2269.940 147.740 2270.260 148.060 ;
        RECT 2752.940 147.740 2753.260 148.060 ;
        RECT 1441.940 145.700 1442.260 146.020 ;
        RECT 1593.740 146.380 1594.060 146.700 ;
        RECT 1538.540 145.700 1538.860 146.020 ;
        RECT 1690.340 146.380 1690.660 146.700 ;
        RECT 1869.740 146.380 1870.060 146.700 ;
        RECT 1593.740 145.020 1594.060 145.340 ;
        RECT 1441.940 144.340 1442.260 144.660 ;
        RECT 1538.540 144.340 1538.860 144.660 ;
        RECT 2317.780 147.060 2318.100 147.380 ;
        RECT 2269.940 145.700 2270.260 146.020 ;
        RECT 2317.780 145.020 2318.100 145.340 ;
        RECT 2510.980 147.060 2511.300 147.380 ;
        RECT 2607.580 147.060 2607.900 147.380 ;
        RECT 2656.340 147.060 2656.660 147.380 ;
        RECT 2510.980 145.020 2511.300 145.340 ;
        RECT 2656.340 145.700 2656.660 146.020 ;
        RECT 2607.580 145.020 2607.900 145.340 ;
        RECT 2752.940 145.700 2753.260 146.020 ;
      LAYER met4 ;
        RECT 1186.175 3196.175 1186.505 3196.505 ;
        RECT 1186.190 146.705 1186.490 3196.175 ;
        RECT 1690.335 147.735 1690.665 148.065 ;
        RECT 1869.735 147.735 1870.065 148.065 ;
        RECT 2269.935 147.735 2270.265 148.065 ;
        RECT 2752.935 147.735 2753.265 148.065 ;
        RECT 1690.350 146.705 1690.650 147.735 ;
        RECT 1869.750 146.705 1870.050 147.735 ;
        RECT 1186.175 146.375 1186.505 146.705 ;
        RECT 1593.735 146.375 1594.065 146.705 ;
        RECT 1690.335 146.375 1690.665 146.705 ;
        RECT 1869.735 146.375 1870.065 146.705 ;
        RECT 1441.935 145.695 1442.265 146.025 ;
        RECT 1538.535 145.695 1538.865 146.025 ;
        RECT 1441.950 144.665 1442.250 145.695 ;
        RECT 1538.550 144.665 1538.850 145.695 ;
        RECT 1593.750 145.345 1594.050 146.375 ;
        RECT 2269.950 146.025 2270.250 147.735 ;
        RECT 2317.775 147.055 2318.105 147.385 ;
        RECT 2510.975 147.055 2511.305 147.385 ;
        RECT 2607.575 147.055 2607.905 147.385 ;
        RECT 2656.335 147.055 2656.665 147.385 ;
        RECT 2269.935 145.695 2270.265 146.025 ;
        RECT 2317.790 145.345 2318.090 147.055 ;
        RECT 2510.990 145.345 2511.290 147.055 ;
        RECT 2607.590 145.345 2607.890 147.055 ;
        RECT 2656.350 146.025 2656.650 147.055 ;
        RECT 2752.950 146.025 2753.250 147.735 ;
        RECT 2656.335 145.695 2656.665 146.025 ;
        RECT 2752.935 145.695 2753.265 146.025 ;
        RECT 1593.735 145.015 1594.065 145.345 ;
        RECT 2317.775 145.015 2318.105 145.345 ;
        RECT 2510.975 145.015 2511.305 145.345 ;
        RECT 2607.575 145.015 2607.905 145.345 ;
        RECT 1441.935 144.335 1442.265 144.665 ;
        RECT 1538.535 144.335 1538.865 144.665 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1576.030 3214.600 1576.350 3214.660 ;
        RECT 2655.190 3214.600 2655.510 3214.660 ;
        RECT 1576.030 3214.460 2655.510 3214.600 ;
        RECT 1576.030 3214.400 1576.350 3214.460 ;
        RECT 2655.190 3214.400 2655.510 3214.460 ;
        RECT 2655.190 2497.540 2655.510 2497.600 ;
        RECT 2900.370 2497.540 2900.690 2497.600 ;
        RECT 2655.190 2497.400 2900.690 2497.540 ;
        RECT 2655.190 2497.340 2655.510 2497.400 ;
        RECT 2900.370 2497.340 2900.690 2497.400 ;
      LAYER via ;
        RECT 1576.060 3214.400 1576.320 3214.660 ;
        RECT 2655.220 3214.400 2655.480 3214.660 ;
        RECT 2655.220 2497.340 2655.480 2497.600 ;
        RECT 2900.400 2497.340 2900.660 2497.600 ;
      LAYER met2 ;
        RECT 1576.060 3214.370 1576.320 3214.690 ;
        RECT 2655.220 3214.370 2655.480 3214.690 ;
        RECT 1576.120 3200.000 1576.260 3214.370 ;
        RECT 1575.980 3196.000 1576.260 3200.000 ;
        RECT 2655.280 2497.630 2655.420 3214.370 ;
        RECT 2655.220 2497.310 2655.480 2497.630 ;
        RECT 2900.400 2497.310 2900.660 2497.630 ;
        RECT 2900.460 2493.405 2900.600 2497.310 ;
        RECT 2900.390 2493.035 2900.670 2493.405 ;
      LAYER via2 ;
        RECT 2900.390 2493.080 2900.670 2493.360 ;
      LAYER met3 ;
        RECT 2900.365 2493.370 2900.695 2493.385 ;
        RECT 2917.600 2493.370 2924.800 2493.820 ;
        RECT 2900.365 2493.070 2924.800 2493.370 ;
        RECT 2900.365 2493.055 2900.695 2493.070 ;
        RECT 2917.600 2492.620 2924.800 2493.070 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1615.590 3214.940 1615.910 3215.000 ;
        RECT 2656.110 3214.940 2656.430 3215.000 ;
        RECT 1615.590 3214.800 2656.430 3214.940 ;
        RECT 1615.590 3214.740 1615.910 3214.800 ;
        RECT 2656.110 3214.740 2656.430 3214.800 ;
        RECT 2656.110 2732.140 2656.430 2732.200 ;
        RECT 2900.370 2732.140 2900.690 2732.200 ;
        RECT 2656.110 2732.000 2900.690 2732.140 ;
        RECT 2656.110 2731.940 2656.430 2732.000 ;
        RECT 2900.370 2731.940 2900.690 2732.000 ;
      LAYER via ;
        RECT 1615.620 3214.740 1615.880 3215.000 ;
        RECT 2656.140 3214.740 2656.400 3215.000 ;
        RECT 2656.140 2731.940 2656.400 2732.200 ;
        RECT 2900.400 2731.940 2900.660 2732.200 ;
      LAYER met2 ;
        RECT 1615.620 3214.710 1615.880 3215.030 ;
        RECT 2656.140 3214.710 2656.400 3215.030 ;
        RECT 1615.680 3200.000 1615.820 3214.710 ;
        RECT 1615.540 3196.000 1615.820 3200.000 ;
        RECT 2656.200 2732.230 2656.340 3214.710 ;
        RECT 2656.140 2731.910 2656.400 2732.230 ;
        RECT 2900.400 2731.910 2900.660 2732.230 ;
        RECT 2900.460 2728.005 2900.600 2731.910 ;
        RECT 2900.390 2727.635 2900.670 2728.005 ;
      LAYER via2 ;
        RECT 2900.390 2727.680 2900.670 2727.960 ;
      LAYER met3 ;
        RECT 2900.365 2727.970 2900.695 2727.985 ;
        RECT 2917.600 2727.970 2924.800 2728.420 ;
        RECT 2900.365 2727.670 2924.800 2727.970 ;
        RECT 2900.365 2727.655 2900.695 2727.670 ;
        RECT 2917.600 2727.220 2924.800 2727.670 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1655.150 3215.280 1655.470 3215.340 ;
        RECT 2651.970 3215.280 2652.290 3215.340 ;
        RECT 1655.150 3215.140 2652.290 3215.280 ;
        RECT 1655.150 3215.080 1655.470 3215.140 ;
        RECT 2651.970 3215.080 2652.290 3215.140 ;
        RECT 2651.970 2966.740 2652.290 2966.800 ;
        RECT 2900.370 2966.740 2900.690 2966.800 ;
        RECT 2651.970 2966.600 2900.690 2966.740 ;
        RECT 2651.970 2966.540 2652.290 2966.600 ;
        RECT 2900.370 2966.540 2900.690 2966.600 ;
      LAYER via ;
        RECT 1655.180 3215.080 1655.440 3215.340 ;
        RECT 2652.000 3215.080 2652.260 3215.340 ;
        RECT 2652.000 2966.540 2652.260 2966.800 ;
        RECT 2900.400 2966.540 2900.660 2966.800 ;
      LAYER met2 ;
        RECT 1655.180 3215.050 1655.440 3215.370 ;
        RECT 2652.000 3215.050 2652.260 3215.370 ;
        RECT 1655.240 3200.000 1655.380 3215.050 ;
        RECT 1655.100 3196.000 1655.380 3200.000 ;
        RECT 2652.060 2966.830 2652.200 3215.050 ;
        RECT 2652.000 2966.510 2652.260 2966.830 ;
        RECT 2900.400 2966.510 2900.660 2966.830 ;
        RECT 2900.460 2962.605 2900.600 2966.510 ;
        RECT 2900.390 2962.235 2900.670 2962.605 ;
      LAYER via2 ;
        RECT 2900.390 2962.280 2900.670 2962.560 ;
      LAYER met3 ;
        RECT 2900.365 2962.570 2900.695 2962.585 ;
        RECT 2917.600 2962.570 2924.800 2963.020 ;
        RECT 2900.365 2962.270 2924.800 2962.570 ;
        RECT 2900.365 2962.255 2900.695 2962.270 ;
        RECT 2917.600 2961.820 2924.800 2962.270 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1696.090 3198.620 1696.410 3198.680 ;
        RECT 2898.990 3198.620 2899.310 3198.680 ;
        RECT 1696.090 3198.480 2899.310 3198.620 ;
        RECT 1696.090 3198.420 1696.410 3198.480 ;
        RECT 2898.990 3198.420 2899.310 3198.480 ;
      LAYER via ;
        RECT 1696.120 3198.420 1696.380 3198.680 ;
        RECT 2899.020 3198.420 2899.280 3198.680 ;
      LAYER met2 ;
        RECT 1694.200 3198.450 1694.480 3200.000 ;
        RECT 1696.120 3198.450 1696.380 3198.710 ;
        RECT 1694.200 3198.390 1696.380 3198.450 ;
        RECT 2899.020 3198.390 2899.280 3198.710 ;
        RECT 1694.200 3198.310 1696.320 3198.390 ;
        RECT 1694.200 3196.000 1694.480 3198.310 ;
        RECT 2899.080 3197.205 2899.220 3198.390 ;
        RECT 2899.010 3196.835 2899.290 3197.205 ;
      LAYER via2 ;
        RECT 2899.010 3196.880 2899.290 3197.160 ;
      LAYER met3 ;
        RECT 2898.985 3197.170 2899.315 3197.185 ;
        RECT 2917.600 3197.170 2924.800 3197.620 ;
        RECT 2898.985 3196.870 2924.800 3197.170 ;
        RECT 2898.985 3196.855 2899.315 3196.870 ;
        RECT 2917.600 3196.420 2924.800 3196.870 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2146.060 3429.680 2149.880 3429.820 ;
        RECT 1738.410 3429.480 1738.730 3429.540 ;
        RECT 2146.060 3429.480 2146.200 3429.680 ;
        RECT 1738.410 3429.340 2146.200 3429.480 ;
        RECT 2149.740 3429.480 2149.880 3429.680 ;
        RECT 2762.920 3429.680 2798.940 3429.820 ;
        RECT 2762.920 3429.480 2763.060 3429.680 ;
        RECT 2149.740 3429.340 2763.060 3429.480 ;
        RECT 2798.800 3429.480 2798.940 3429.680 ;
        RECT 2900.830 3429.480 2901.150 3429.540 ;
        RECT 2798.800 3429.340 2901.150 3429.480 ;
        RECT 1738.410 3429.280 1738.730 3429.340 ;
        RECT 2900.830 3429.280 2901.150 3429.340 ;
      LAYER via ;
        RECT 1738.440 3429.280 1738.700 3429.540 ;
        RECT 2900.860 3429.280 2901.120 3429.540 ;
      LAYER met2 ;
        RECT 2900.850 3431.435 2901.130 3431.805 ;
        RECT 2900.920 3429.570 2901.060 3431.435 ;
        RECT 1738.440 3429.250 1738.700 3429.570 ;
        RECT 2900.860 3429.250 2901.120 3429.570 ;
        RECT 1738.500 3200.490 1738.640 3429.250 ;
        RECT 1735.740 3200.350 1738.640 3200.490 ;
        RECT 1733.760 3199.810 1734.040 3200.000 ;
        RECT 1735.740 3199.810 1735.880 3200.350 ;
        RECT 1733.760 3199.670 1735.880 3199.810 ;
        RECT 1733.760 3196.000 1734.040 3199.670 ;
      LAYER via2 ;
        RECT 2900.850 3431.480 2901.130 3431.760 ;
      LAYER met3 ;
        RECT 2900.825 3431.770 2901.155 3431.785 ;
        RECT 2917.600 3431.770 2924.800 3432.220 ;
        RECT 2900.825 3431.470 2924.800 3431.770 ;
        RECT 2900.825 3431.455 2901.155 3431.470 ;
        RECT 2917.600 3431.020 2924.800 3431.470 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1779.810 3504.620 1780.130 3504.680 ;
        RECT 2717.290 3504.620 2717.610 3504.680 ;
        RECT 1779.810 3504.480 2717.610 3504.620 ;
        RECT 1779.810 3504.420 1780.130 3504.480 ;
        RECT 2717.290 3504.420 2717.610 3504.480 ;
      LAYER via ;
        RECT 1779.840 3504.420 1780.100 3504.680 ;
        RECT 2717.320 3504.420 2717.580 3504.680 ;
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
        RECT 2717.380 3504.710 2717.520 3517.600 ;
        RECT 1779.840 3504.390 1780.100 3504.710 ;
        RECT 2717.320 3504.390 2717.580 3504.710 ;
        RECT 1779.900 3200.490 1780.040 3504.390 ;
        RECT 1776.680 3200.350 1780.040 3200.490 ;
        RECT 1773.320 3199.810 1773.600 3200.000 ;
        RECT 1776.680 3199.810 1776.820 3200.350 ;
        RECT 1773.320 3199.670 1776.820 3199.810 ;
        RECT 1773.320 3196.000 1773.600 3199.670 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1814.310 3500.540 1814.630 3500.600 ;
        RECT 2392.530 3500.540 2392.850 3500.600 ;
        RECT 1814.310 3500.400 2392.850 3500.540 ;
        RECT 1814.310 3500.340 1814.630 3500.400 ;
        RECT 2392.530 3500.340 2392.850 3500.400 ;
      LAYER via ;
        RECT 1814.340 3500.340 1814.600 3500.600 ;
        RECT 2392.560 3500.340 2392.820 3500.600 ;
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
        RECT 2392.620 3500.630 2392.760 3517.600 ;
        RECT 1814.340 3500.310 1814.600 3500.630 ;
        RECT 2392.560 3500.310 2392.820 3500.630 ;
        RECT 1812.880 3199.810 1813.160 3200.000 ;
        RECT 1814.400 3199.810 1814.540 3500.310 ;
        RECT 1812.880 3199.670 1814.540 3199.810 ;
        RECT 1812.880 3196.000 1813.160 3199.670 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1855.710 3499.180 1856.030 3499.240 ;
        RECT 2068.230 3499.180 2068.550 3499.240 ;
        RECT 1855.710 3499.040 2068.550 3499.180 ;
        RECT 1855.710 3498.980 1856.030 3499.040 ;
        RECT 2068.230 3498.980 2068.550 3499.040 ;
      LAYER via ;
        RECT 1855.740 3498.980 1856.000 3499.240 ;
        RECT 2068.260 3498.980 2068.520 3499.240 ;
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
        RECT 2068.320 3499.270 2068.460 3517.600 ;
        RECT 1855.740 3498.950 1856.000 3499.270 ;
        RECT 2068.260 3498.950 2068.520 3499.270 ;
        RECT 1852.440 3199.130 1852.720 3200.000 ;
        RECT 1855.800 3199.130 1855.940 3498.950 ;
        RECT 1852.440 3198.990 1855.940 3199.130 ;
        RECT 1852.440 3196.000 1852.720 3198.990 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1743.930 3498.840 1744.250 3498.900 ;
        RECT 1890.670 3498.840 1890.990 3498.900 ;
        RECT 1743.930 3498.700 1890.990 3498.840 ;
        RECT 1743.930 3498.640 1744.250 3498.700 ;
        RECT 1890.670 3498.640 1890.990 3498.700 ;
      LAYER via ;
        RECT 1743.960 3498.640 1744.220 3498.900 ;
        RECT 1890.700 3498.640 1890.960 3498.900 ;
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
        RECT 1744.020 3498.930 1744.160 3517.600 ;
        RECT 1743.960 3498.610 1744.220 3498.930 ;
        RECT 1890.700 3498.610 1890.960 3498.930 ;
        RECT 1890.760 3199.810 1890.900 3498.610 ;
        RECT 1891.540 3199.810 1891.820 3200.000 ;
        RECT 1890.760 3199.670 1891.820 3199.810 ;
        RECT 1891.540 3196.000 1891.820 3199.670 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1419.170 3499.860 1419.490 3499.920 ;
        RECT 1925.170 3499.860 1925.490 3499.920 ;
        RECT 1419.170 3499.720 1925.490 3499.860 ;
        RECT 1419.170 3499.660 1419.490 3499.720 ;
        RECT 1925.170 3499.660 1925.490 3499.720 ;
      LAYER via ;
        RECT 1419.200 3499.660 1419.460 3499.920 ;
        RECT 1925.200 3499.660 1925.460 3499.920 ;
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
        RECT 1419.260 3499.950 1419.400 3517.600 ;
        RECT 1419.200 3499.630 1419.460 3499.950 ;
        RECT 1925.200 3499.630 1925.460 3499.950 ;
        RECT 1925.260 3200.490 1925.400 3499.630 ;
        RECT 1925.260 3200.350 1928.160 3200.490 ;
        RECT 1928.020 3199.810 1928.160 3200.350 ;
        RECT 1931.100 3199.810 1931.380 3200.000 ;
        RECT 1928.020 3199.670 1931.380 3199.810 ;
        RECT 1931.100 3196.000 1931.380 3199.670 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1993.710 381.380 1994.030 381.440 ;
        RECT 2028.210 381.380 2028.530 381.440 ;
        RECT 1993.710 381.240 2028.530 381.380 ;
        RECT 1993.710 381.180 1994.030 381.240 ;
        RECT 2028.210 381.180 2028.530 381.240 ;
        RECT 1545.210 381.040 1545.530 381.100 ;
        RECT 1586.610 381.040 1586.930 381.100 ;
        RECT 1545.210 380.900 1586.930 381.040 ;
        RECT 1545.210 380.840 1545.530 380.900 ;
        RECT 1586.610 380.840 1586.930 380.900 ;
        RECT 2572.850 380.700 2573.170 380.760 ;
        RECT 2584.350 380.700 2584.670 380.760 ;
        RECT 2572.850 380.560 2584.670 380.700 ;
        RECT 2572.850 380.500 2573.170 380.560 ;
        RECT 2584.350 380.500 2584.670 380.560 ;
        RECT 2379.650 380.360 2379.970 380.420 ;
        RECT 2390.690 380.360 2391.010 380.420 ;
        RECT 2379.650 380.220 2391.010 380.360 ;
        RECT 2379.650 380.160 2379.970 380.220 ;
        RECT 2390.690 380.160 2391.010 380.220 ;
        RECT 1417.330 380.020 1417.650 380.080 ;
        RECT 1452.750 380.020 1453.070 380.080 ;
        RECT 1417.330 379.880 1453.070 380.020 ;
        RECT 1417.330 379.820 1417.650 379.880 ;
        RECT 1452.750 379.820 1453.070 379.880 ;
        RECT 2621.150 380.020 2621.470 380.080 ;
        RECT 2632.190 380.020 2632.510 380.080 ;
        RECT 2621.150 379.880 2632.510 380.020 ;
        RECT 2621.150 379.820 2621.470 379.880 ;
        RECT 2632.190 379.820 2632.510 379.880 ;
      LAYER via ;
        RECT 1993.740 381.180 1994.000 381.440 ;
        RECT 2028.240 381.180 2028.500 381.440 ;
        RECT 1545.240 380.840 1545.500 381.100 ;
        RECT 1586.640 380.840 1586.900 381.100 ;
        RECT 2572.880 380.500 2573.140 380.760 ;
        RECT 2584.380 380.500 2584.640 380.760 ;
        RECT 2379.680 380.160 2379.940 380.420 ;
        RECT 2390.720 380.160 2390.980 380.420 ;
        RECT 1417.360 379.820 1417.620 380.080 ;
        RECT 1452.780 379.820 1453.040 380.080 ;
        RECT 2621.180 379.820 2621.440 380.080 ;
        RECT 2632.220 379.820 2632.480 380.080 ;
      LAYER met2 ;
        RECT 1220.010 3196.410 1220.290 3196.525 ;
        RECT 1220.860 3196.410 1221.140 3200.000 ;
        RECT 1220.010 3196.270 1221.140 3196.410 ;
        RECT 1220.010 3196.155 1220.290 3196.270 ;
        RECT 1220.860 3196.000 1221.140 3196.270 ;
        RECT 1265.550 382.315 1265.830 382.685 ;
        RECT 1265.620 379.965 1265.760 382.315 ;
        RECT 2704.430 381.635 2704.710 382.005 ;
        RECT 1993.740 381.325 1994.000 381.470 ;
        RECT 2028.240 381.325 2028.500 381.470 ;
        RECT 1545.230 380.955 1545.510 381.325 ;
        RECT 1586.630 380.955 1586.910 381.325 ;
        RECT 1593.530 380.955 1593.810 381.325 ;
        RECT 1993.730 380.955 1994.010 381.325 ;
        RECT 2028.230 380.955 2028.510 381.325 ;
        RECT 2090.330 380.955 2090.610 381.325 ;
        RECT 1545.240 380.810 1545.500 380.955 ;
        RECT 1586.640 380.810 1586.900 380.955 ;
        RECT 1593.600 380.645 1593.740 380.955 ;
        RECT 1593.530 380.275 1593.810 380.645 ;
        RECT 2090.400 380.530 2090.540 380.955 ;
        RECT 2572.880 380.645 2573.140 380.790 ;
        RECT 2584.380 380.645 2584.640 380.790 ;
        RECT 2090.790 380.530 2091.070 380.645 ;
        RECT 2090.400 380.390 2091.070 380.530 ;
        RECT 2090.790 380.275 2091.070 380.390 ;
        RECT 2283.530 380.530 2283.810 380.645 ;
        RECT 2284.450 380.530 2284.730 380.645 ;
        RECT 2283.530 380.390 2284.730 380.530 ;
        RECT 2283.530 380.275 2283.810 380.390 ;
        RECT 2284.450 380.275 2284.730 380.390 ;
        RECT 2379.670 380.275 2379.950 380.645 ;
        RECT 2390.710 380.275 2390.990 380.645 ;
        RECT 2572.870 380.275 2573.150 380.645 ;
        RECT 2584.370 380.275 2584.650 380.645 ;
        RECT 2632.210 380.275 2632.490 380.645 ;
        RECT 2379.680 380.130 2379.940 380.275 ;
        RECT 2390.720 380.130 2390.980 380.275 ;
        RECT 2632.280 380.110 2632.420 380.275 ;
        RECT 1417.360 379.965 1417.620 380.110 ;
        RECT 1265.550 379.595 1265.830 379.965 ;
        RECT 1417.350 379.595 1417.630 379.965 ;
        RECT 1452.780 379.790 1453.040 380.110 ;
        RECT 2621.180 379.965 2621.440 380.110 ;
        RECT 1452.840 379.285 1452.980 379.790 ;
        RECT 2621.170 379.595 2621.450 379.965 ;
        RECT 2632.220 379.790 2632.480 380.110 ;
        RECT 2704.500 379.965 2704.640 381.635 ;
        RECT 2801.030 380.955 2801.310 381.325 ;
        RECT 2704.430 379.595 2704.710 379.965 ;
        RECT 2801.100 379.285 2801.240 380.955 ;
        RECT 2863.130 380.275 2863.410 380.645 ;
        RECT 2863.200 379.850 2863.340 380.275 ;
        RECT 2863.590 379.850 2863.870 379.965 ;
        RECT 2863.200 379.710 2863.870 379.850 ;
        RECT 2863.590 379.595 2863.870 379.710 ;
        RECT 1452.770 378.915 1453.050 379.285 ;
        RECT 2801.030 378.915 2801.310 379.285 ;
      LAYER via2 ;
        RECT 1220.010 3196.200 1220.290 3196.480 ;
        RECT 1265.550 382.360 1265.830 382.640 ;
        RECT 2704.430 381.680 2704.710 381.960 ;
        RECT 1545.230 381.000 1545.510 381.280 ;
        RECT 1586.630 381.000 1586.910 381.280 ;
        RECT 1593.530 381.000 1593.810 381.280 ;
        RECT 1993.730 381.000 1994.010 381.280 ;
        RECT 2028.230 381.000 2028.510 381.280 ;
        RECT 2090.330 381.000 2090.610 381.280 ;
        RECT 1593.530 380.320 1593.810 380.600 ;
        RECT 2090.790 380.320 2091.070 380.600 ;
        RECT 2283.530 380.320 2283.810 380.600 ;
        RECT 2284.450 380.320 2284.730 380.600 ;
        RECT 2379.670 380.320 2379.950 380.600 ;
        RECT 2390.710 380.320 2390.990 380.600 ;
        RECT 2572.870 380.320 2573.150 380.600 ;
        RECT 2584.370 380.320 2584.650 380.600 ;
        RECT 2632.210 380.320 2632.490 380.600 ;
        RECT 1265.550 379.640 1265.830 379.920 ;
        RECT 1417.350 379.640 1417.630 379.920 ;
        RECT 2621.170 379.640 2621.450 379.920 ;
        RECT 2801.030 381.000 2801.310 381.280 ;
        RECT 2704.430 379.640 2704.710 379.920 ;
        RECT 2863.130 380.320 2863.410 380.600 ;
        RECT 2863.590 379.640 2863.870 379.920 ;
        RECT 1452.770 378.960 1453.050 379.240 ;
        RECT 2801.030 378.960 2801.310 379.240 ;
      LAYER met3 ;
        RECT 1219.985 3196.500 1220.315 3196.505 ;
        RECT 1219.985 3196.490 1220.570 3196.500 ;
        RECT 1219.985 3196.190 1220.770 3196.490 ;
        RECT 1219.985 3196.180 1220.570 3196.190 ;
        RECT 1219.985 3196.175 1220.315 3196.180 ;
        RECT 1265.525 382.650 1265.855 382.665 ;
        RECT 1265.525 382.350 1290.450 382.650 ;
        RECT 1265.525 382.335 1265.855 382.350 ;
        RECT 1290.150 381.970 1290.450 382.350 ;
        RECT 1786.910 381.970 1787.290 381.980 ;
        RECT 2656.310 381.970 2656.690 381.980 ;
        RECT 2704.405 381.970 2704.735 381.985 ;
        RECT 1290.150 381.670 1318.970 381.970 ;
        RECT 1318.670 380.610 1318.970 381.670 ;
        RECT 1594.670 381.670 1707.210 381.970 ;
        RECT 1545.205 381.290 1545.535 381.305 ;
        RECT 1521.070 380.990 1545.535 381.290 ;
        RECT 1318.670 380.310 1366.810 380.610 ;
        RECT 1220.190 379.930 1220.570 379.940 ;
        RECT 1265.525 379.930 1265.855 379.945 ;
        RECT 1220.190 379.630 1265.855 379.930 ;
        RECT 1366.510 379.930 1366.810 380.310 ;
        RECT 1417.325 379.930 1417.655 379.945 ;
        RECT 1366.510 379.630 1417.655 379.930 ;
        RECT 1220.190 379.620 1220.570 379.630 ;
        RECT 1265.525 379.615 1265.855 379.630 ;
        RECT 1417.325 379.615 1417.655 379.630 ;
        RECT 1452.745 379.250 1453.075 379.265 ;
        RECT 1521.070 379.250 1521.370 380.990 ;
        RECT 1545.205 380.975 1545.535 380.990 ;
        RECT 1586.605 381.290 1586.935 381.305 ;
        RECT 1593.505 381.290 1593.835 381.305 ;
        RECT 1594.670 381.290 1594.970 381.670 ;
        RECT 1586.605 380.990 1594.970 381.290 ;
        RECT 1586.605 380.975 1586.935 380.990 ;
        RECT 1593.505 380.975 1594.050 380.990 ;
        RECT 1593.750 380.625 1594.050 380.975 ;
        RECT 1593.505 380.310 1594.050 380.625 ;
        RECT 1706.910 380.610 1707.210 381.670 ;
        RECT 1786.910 381.670 1852.570 381.970 ;
        RECT 1786.910 381.660 1787.290 381.670 ;
        RECT 1786.910 380.610 1787.290 380.620 ;
        RECT 1706.910 380.310 1715.490 380.610 ;
        RECT 1593.505 380.295 1593.835 380.310 ;
        RECT 1715.190 379.930 1715.490 380.310 ;
        RECT 1752.910 380.310 1787.290 380.610 ;
        RECT 1852.270 380.610 1852.570 381.670 ;
        RECT 2125.510 381.670 2138.690 381.970 ;
        RECT 1993.705 381.290 1994.035 381.305 ;
        RECT 1946.110 380.990 1994.035 381.290 ;
        RECT 1883.510 380.610 1883.890 380.620 ;
        RECT 1852.270 380.310 1883.890 380.610 ;
        RECT 1715.190 379.760 1752.290 379.930 ;
        RECT 1752.910 379.760 1753.210 380.310 ;
        RECT 1786.910 380.300 1787.290 380.310 ;
        RECT 1883.510 380.300 1883.890 380.310 ;
        RECT 1884.430 380.610 1884.810 380.620 ;
        RECT 1946.110 380.610 1946.410 380.990 ;
        RECT 1993.705 380.975 1994.035 380.990 ;
        RECT 2028.205 381.290 2028.535 381.305 ;
        RECT 2090.305 381.290 2090.635 381.305 ;
        RECT 2125.510 381.290 2125.810 381.670 ;
        RECT 2028.205 380.990 2042.090 381.290 ;
        RECT 2028.205 380.975 2028.535 380.990 ;
        RECT 1884.430 380.310 1946.410 380.610 ;
        RECT 1884.430 380.300 1884.810 380.310 ;
        RECT 1715.190 379.630 1753.210 379.760 ;
        RECT 2041.790 379.930 2042.090 380.990 ;
        RECT 2076.750 380.990 2090.635 381.290 ;
        RECT 2076.750 380.610 2077.050 380.990 ;
        RECT 2090.305 380.975 2090.635 380.990 ;
        RECT 2124.590 380.990 2125.810 381.290 ;
        RECT 2138.390 381.290 2138.690 381.670 ;
        RECT 2476.030 381.670 2511.290 381.970 ;
        RECT 2138.390 380.990 2187.450 381.290 ;
        RECT 2042.710 380.310 2077.050 380.610 ;
        RECT 2090.765 380.610 2091.095 380.625 ;
        RECT 2124.590 380.610 2124.890 380.990 ;
        RECT 2090.765 380.310 2124.890 380.610 ;
        RECT 2042.710 379.930 2043.010 380.310 ;
        RECT 2090.765 380.295 2091.095 380.310 ;
        RECT 2041.790 379.630 2043.010 379.930 ;
        RECT 2187.150 379.930 2187.450 380.990 ;
        RECT 2283.505 380.610 2283.835 380.625 ;
        RECT 2235.910 380.310 2283.835 380.610 ;
        RECT 2235.910 379.930 2236.210 380.310 ;
        RECT 2283.505 380.295 2283.835 380.310 ;
        RECT 2284.425 380.610 2284.755 380.625 ;
        RECT 2379.645 380.610 2379.975 380.625 ;
        RECT 2284.425 380.310 2331.890 380.610 ;
        RECT 2284.425 380.295 2284.755 380.310 ;
        RECT 2187.150 379.630 2236.210 379.930 ;
        RECT 2331.590 379.930 2331.890 380.310 ;
        RECT 2332.510 380.310 2379.975 380.610 ;
        RECT 2332.510 379.930 2332.810 380.310 ;
        RECT 2379.645 380.295 2379.975 380.310 ;
        RECT 2390.685 380.610 2391.015 380.625 ;
        RECT 2476.030 380.610 2476.330 381.670 ;
        RECT 2390.685 380.310 2414.690 380.610 ;
        RECT 2390.685 380.295 2391.015 380.310 ;
        RECT 2331.590 379.630 2332.810 379.930 ;
        RECT 2414.390 379.930 2414.690 380.310 ;
        RECT 2429.110 380.310 2476.330 380.610 ;
        RECT 2429.110 379.930 2429.410 380.310 ;
        RECT 2414.390 379.630 2429.410 379.930 ;
        RECT 2510.990 379.930 2511.290 381.670 ;
        RECT 2656.310 381.670 2704.735 381.970 ;
        RECT 2656.310 381.660 2656.690 381.670 ;
        RECT 2704.405 381.655 2704.735 381.670 ;
        RECT 2801.005 381.290 2801.335 381.305 ;
        RECT 2917.600 381.290 2924.800 381.740 ;
        RECT 2801.005 380.990 2815.810 381.290 ;
        RECT 2801.005 380.975 2801.335 380.990 ;
        RECT 2572.845 380.610 2573.175 380.625 ;
        RECT 2525.710 380.310 2573.175 380.610 ;
        RECT 2525.710 379.930 2526.010 380.310 ;
        RECT 2572.845 380.295 2573.175 380.310 ;
        RECT 2584.345 380.610 2584.675 380.625 ;
        RECT 2632.185 380.610 2632.515 380.625 ;
        RECT 2656.310 380.610 2656.690 380.620 ;
        RECT 2752.910 380.610 2753.290 380.620 ;
        RECT 2584.345 380.310 2607.890 380.610 ;
        RECT 2584.345 380.295 2584.675 380.310 ;
        RECT 2510.990 379.630 2526.010 379.930 ;
        RECT 2607.590 379.930 2607.890 380.310 ;
        RECT 2632.185 380.310 2656.690 380.610 ;
        RECT 2632.185 380.295 2632.515 380.310 ;
        RECT 2656.310 380.300 2656.690 380.310 ;
        RECT 2718.910 380.310 2753.290 380.610 ;
        RECT 2621.145 379.930 2621.475 379.945 ;
        RECT 2607.590 379.630 2621.475 379.930 ;
        RECT 1751.990 379.460 1753.210 379.630 ;
        RECT 2621.145 379.615 2621.475 379.630 ;
        RECT 2704.405 379.930 2704.735 379.945 ;
        RECT 2718.910 379.930 2719.210 380.310 ;
        RECT 2752.910 380.300 2753.290 380.310 ;
        RECT 2704.405 379.630 2719.210 379.930 ;
        RECT 2815.510 379.930 2815.810 380.990 ;
        RECT 2916.710 380.990 2924.800 381.290 ;
        RECT 2863.105 380.610 2863.435 380.625 ;
        RECT 2916.710 380.610 2917.010 380.990 ;
        RECT 2849.550 380.310 2863.435 380.610 ;
        RECT 2849.550 379.930 2849.850 380.310 ;
        RECT 2863.105 380.295 2863.435 380.310 ;
        RECT 2884.510 380.310 2917.010 380.610 ;
        RECT 2917.600 380.540 2924.800 380.990 ;
        RECT 2815.510 379.630 2849.850 379.930 ;
        RECT 2863.565 379.930 2863.895 379.945 ;
        RECT 2884.510 379.930 2884.810 380.310 ;
        RECT 2863.565 379.630 2884.810 379.930 ;
        RECT 2704.405 379.615 2704.735 379.630 ;
        RECT 2863.565 379.615 2863.895 379.630 ;
        RECT 1452.745 378.950 1521.370 379.250 ;
        RECT 2752.910 379.250 2753.290 379.260 ;
        RECT 2801.005 379.250 2801.335 379.265 ;
        RECT 2752.910 378.950 2801.335 379.250 ;
        RECT 1452.745 378.935 1453.075 378.950 ;
        RECT 2752.910 378.940 2753.290 378.950 ;
        RECT 2801.005 378.935 2801.335 378.950 ;
      LAYER via3 ;
        RECT 1220.220 3196.180 1220.540 3196.500 ;
        RECT 1220.220 379.620 1220.540 379.940 ;
        RECT 1786.940 381.660 1787.260 381.980 ;
        RECT 1786.940 380.300 1787.260 380.620 ;
        RECT 1883.540 380.300 1883.860 380.620 ;
        RECT 1884.460 380.300 1884.780 380.620 ;
        RECT 2656.340 381.660 2656.660 381.980 ;
        RECT 2656.340 380.300 2656.660 380.620 ;
        RECT 2752.940 380.300 2753.260 380.620 ;
        RECT 2752.940 378.940 2753.260 379.260 ;
      LAYER met4 ;
        RECT 1220.215 3196.175 1220.545 3196.505 ;
        RECT 1220.230 379.945 1220.530 3196.175 ;
        RECT 1786.935 381.655 1787.265 381.985 ;
        RECT 2656.335 381.655 2656.665 381.985 ;
        RECT 1786.950 380.625 1787.250 381.655 ;
        RECT 2656.350 380.625 2656.650 381.655 ;
        RECT 1786.935 380.295 1787.265 380.625 ;
        RECT 1883.535 380.295 1883.865 380.625 ;
        RECT 1884.455 380.295 1884.785 380.625 ;
        RECT 2656.335 380.295 2656.665 380.625 ;
        RECT 2752.935 380.295 2753.265 380.625 ;
        RECT 1220.215 379.615 1220.545 379.945 ;
        RECT 1883.550 379.250 1883.850 380.295 ;
        RECT 1884.470 379.250 1884.770 380.295 ;
        RECT 2752.950 379.265 2753.250 380.295 ;
        RECT 1883.550 378.950 1884.770 379.250 ;
        RECT 2752.935 378.935 2753.265 379.265 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1094.870 3504.960 1095.190 3505.020 ;
        RECT 1966.570 3504.960 1966.890 3505.020 ;
        RECT 1094.870 3504.820 1966.890 3504.960 ;
        RECT 1094.870 3504.760 1095.190 3504.820 ;
        RECT 1966.570 3504.760 1966.890 3504.820 ;
      LAYER via ;
        RECT 1094.900 3504.760 1095.160 3505.020 ;
        RECT 1966.600 3504.760 1966.860 3505.020 ;
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
        RECT 1094.960 3505.050 1095.100 3517.600 ;
        RECT 1094.900 3504.730 1095.160 3505.050 ;
        RECT 1966.600 3504.730 1966.860 3505.050 ;
        RECT 1966.660 3199.810 1966.800 3504.730 ;
        RECT 1970.660 3199.810 1970.940 3200.000 ;
        RECT 1966.660 3199.670 1970.940 3199.810 ;
        RECT 1970.660 3196.000 1970.940 3199.670 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 770.570 3503.600 770.890 3503.660 ;
        RECT 2007.970 3503.600 2008.290 3503.660 ;
        RECT 770.570 3503.460 2008.290 3503.600 ;
        RECT 770.570 3503.400 770.890 3503.460 ;
        RECT 2007.970 3503.400 2008.290 3503.460 ;
      LAYER via ;
        RECT 770.600 3503.400 770.860 3503.660 ;
        RECT 2008.000 3503.400 2008.260 3503.660 ;
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
        RECT 770.660 3503.690 770.800 3517.600 ;
        RECT 770.600 3503.370 770.860 3503.690 ;
        RECT 2008.000 3503.370 2008.260 3503.690 ;
        RECT 2008.060 3199.810 2008.200 3503.370 ;
        RECT 2010.220 3199.810 2010.500 3200.000 ;
        RECT 2008.060 3199.670 2010.500 3199.810 ;
        RECT 2010.220 3196.000 2010.500 3199.670 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 445.810 3502.580 446.130 3502.640 ;
        RECT 2049.370 3502.580 2049.690 3502.640 ;
        RECT 445.810 3502.440 2049.690 3502.580 ;
        RECT 445.810 3502.380 446.130 3502.440 ;
        RECT 2049.370 3502.380 2049.690 3502.440 ;
      LAYER via ;
        RECT 445.840 3502.380 446.100 3502.640 ;
        RECT 2049.400 3502.380 2049.660 3502.640 ;
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
        RECT 445.900 3502.670 446.040 3517.600 ;
        RECT 445.840 3502.350 446.100 3502.670 ;
        RECT 2049.400 3502.350 2049.660 3502.670 ;
        RECT 2049.460 3199.810 2049.600 3502.350 ;
        RECT 2049.780 3199.810 2050.060 3200.000 ;
        RECT 2049.460 3199.670 2050.060 3199.810 ;
        RECT 2049.780 3196.000 2050.060 3199.670 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 121.510 3501.560 121.830 3501.620 ;
        RECT 2083.870 3501.560 2084.190 3501.620 ;
        RECT 121.510 3501.420 2084.190 3501.560 ;
        RECT 121.510 3501.360 121.830 3501.420 ;
        RECT 2083.870 3501.360 2084.190 3501.420 ;
      LAYER via ;
        RECT 121.540 3501.360 121.800 3501.620 ;
        RECT 2083.900 3501.360 2084.160 3501.620 ;
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
        RECT 121.600 3501.650 121.740 3517.600 ;
        RECT 121.540 3501.330 121.800 3501.650 ;
        RECT 2083.900 3501.330 2084.160 3501.650 ;
        RECT 2083.960 3199.130 2084.100 3501.330 ;
        RECT 2088.880 3199.130 2089.160 3200.000 ;
        RECT 2083.960 3198.990 2089.160 3199.130 ;
        RECT 2088.880 3196.000 2089.160 3198.990 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 3339.720 17.410 3339.780 ;
        RECT 2125.270 3339.720 2125.590 3339.780 ;
        RECT 17.090 3339.580 2125.590 3339.720 ;
        RECT 17.090 3339.520 17.410 3339.580 ;
        RECT 2125.270 3339.520 2125.590 3339.580 ;
      LAYER via ;
        RECT 17.120 3339.520 17.380 3339.780 ;
        RECT 2125.300 3339.520 2125.560 3339.780 ;
      LAYER met2 ;
        RECT 17.110 3339.635 17.390 3340.005 ;
        RECT 17.120 3339.490 17.380 3339.635 ;
        RECT 2125.300 3339.490 2125.560 3339.810 ;
        RECT 2125.360 3199.130 2125.500 3339.490 ;
        RECT 2128.440 3199.130 2128.720 3200.000 ;
        RECT 2125.360 3198.990 2128.720 3199.130 ;
        RECT 2128.440 3196.000 2128.720 3198.990 ;
      LAYER via2 ;
        RECT 17.110 3339.680 17.390 3339.960 ;
      LAYER met3 ;
        RECT -4.800 3339.970 2.400 3340.420 ;
        RECT 17.085 3339.970 17.415 3339.985 ;
        RECT -4.800 3339.670 17.415 3339.970 ;
        RECT -4.800 3339.220 2.400 3339.670 ;
        RECT 17.085 3339.655 17.415 3339.670 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 27.210 3213.240 27.530 3213.300 ;
        RECT 2168.050 3213.240 2168.370 3213.300 ;
        RECT 27.210 3213.100 2168.370 3213.240 ;
        RECT 27.210 3213.040 27.530 3213.100 ;
        RECT 2168.050 3213.040 2168.370 3213.100 ;
        RECT 13.870 3052.760 14.190 3052.820 ;
        RECT 27.210 3052.760 27.530 3052.820 ;
        RECT 13.870 3052.620 27.530 3052.760 ;
        RECT 13.870 3052.560 14.190 3052.620 ;
        RECT 27.210 3052.560 27.530 3052.620 ;
      LAYER via ;
        RECT 27.240 3213.040 27.500 3213.300 ;
        RECT 2168.080 3213.040 2168.340 3213.300 ;
        RECT 13.900 3052.560 14.160 3052.820 ;
        RECT 27.240 3052.560 27.500 3052.820 ;
      LAYER met2 ;
        RECT 27.240 3213.010 27.500 3213.330 ;
        RECT 2168.080 3213.010 2168.340 3213.330 ;
        RECT 27.300 3052.850 27.440 3213.010 ;
        RECT 2168.140 3200.000 2168.280 3213.010 ;
        RECT 2168.000 3196.000 2168.280 3200.000 ;
        RECT 13.900 3052.530 14.160 3052.850 ;
        RECT 27.240 3052.530 27.500 3052.850 ;
        RECT 13.960 3052.365 14.100 3052.530 ;
        RECT 13.890 3051.995 14.170 3052.365 ;
      LAYER via2 ;
        RECT 13.890 3052.040 14.170 3052.320 ;
      LAYER met3 ;
        RECT -4.800 3052.330 2.400 3052.780 ;
        RECT 13.865 3052.330 14.195 3052.345 ;
        RECT -4.800 3052.030 14.195 3052.330 ;
        RECT -4.800 3051.580 2.400 3052.030 ;
        RECT 13.865 3052.015 14.195 3052.030 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 26.750 3212.900 27.070 3212.960 ;
        RECT 2207.610 3212.900 2207.930 3212.960 ;
        RECT 26.750 3212.760 2207.930 3212.900 ;
        RECT 26.750 3212.700 27.070 3212.760 ;
        RECT 2207.610 3212.700 2207.930 3212.760 ;
        RECT 13.870 2765.460 14.190 2765.520 ;
        RECT 26.750 2765.460 27.070 2765.520 ;
        RECT 13.870 2765.320 27.070 2765.460 ;
        RECT 13.870 2765.260 14.190 2765.320 ;
        RECT 26.750 2765.260 27.070 2765.320 ;
      LAYER via ;
        RECT 26.780 3212.700 27.040 3212.960 ;
        RECT 2207.640 3212.700 2207.900 3212.960 ;
        RECT 13.900 2765.260 14.160 2765.520 ;
        RECT 26.780 2765.260 27.040 2765.520 ;
      LAYER met2 ;
        RECT 26.780 3212.670 27.040 3212.990 ;
        RECT 2207.640 3212.670 2207.900 3212.990 ;
        RECT 26.840 2765.550 26.980 3212.670 ;
        RECT 2207.700 3200.000 2207.840 3212.670 ;
        RECT 2207.560 3196.000 2207.840 3200.000 ;
        RECT 13.900 2765.405 14.160 2765.550 ;
        RECT 13.890 2765.035 14.170 2765.405 ;
        RECT 26.780 2765.230 27.040 2765.550 ;
      LAYER via2 ;
        RECT 13.890 2765.080 14.170 2765.360 ;
      LAYER met3 ;
        RECT -4.800 2765.370 2.400 2765.820 ;
        RECT 13.865 2765.370 14.195 2765.385 ;
        RECT -4.800 2765.070 14.195 2765.370 ;
        RECT -4.800 2764.620 2.400 2765.070 ;
        RECT 13.865 2765.055 14.195 2765.070 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 25.830 3211.880 26.150 3211.940 ;
        RECT 2247.170 3211.880 2247.490 3211.940 ;
        RECT 25.830 3211.740 2247.490 3211.880 ;
        RECT 25.830 3211.680 26.150 3211.740 ;
        RECT 2247.170 3211.680 2247.490 3211.740 ;
        RECT 13.870 2482.240 14.190 2482.300 ;
        RECT 25.830 2482.240 26.150 2482.300 ;
        RECT 13.870 2482.100 26.150 2482.240 ;
        RECT 13.870 2482.040 14.190 2482.100 ;
        RECT 25.830 2482.040 26.150 2482.100 ;
      LAYER via ;
        RECT 25.860 3211.680 26.120 3211.940 ;
        RECT 2247.200 3211.680 2247.460 3211.940 ;
        RECT 13.900 2482.040 14.160 2482.300 ;
        RECT 25.860 2482.040 26.120 2482.300 ;
      LAYER met2 ;
        RECT 25.860 3211.650 26.120 3211.970 ;
        RECT 2247.200 3211.650 2247.460 3211.970 ;
        RECT 25.920 2482.330 26.060 3211.650 ;
        RECT 2247.260 3200.000 2247.400 3211.650 ;
        RECT 2247.120 3196.000 2247.400 3200.000 ;
        RECT 13.900 2482.010 14.160 2482.330 ;
        RECT 25.860 2482.010 26.120 2482.330 ;
        RECT 13.960 2477.765 14.100 2482.010 ;
        RECT 13.890 2477.395 14.170 2477.765 ;
      LAYER via2 ;
        RECT 13.890 2477.440 14.170 2477.720 ;
      LAYER met3 ;
        RECT -4.800 2477.730 2.400 2478.180 ;
        RECT 13.865 2477.730 14.195 2477.745 ;
        RECT -4.800 2477.430 14.195 2477.730 ;
        RECT -4.800 2476.980 2.400 2477.430 ;
        RECT 13.865 2477.415 14.195 2477.430 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 13.870 2190.180 14.190 2190.240 ;
        RECT 26.290 2190.180 26.610 2190.240 ;
        RECT 13.870 2190.040 26.610 2190.180 ;
        RECT 13.870 2189.980 14.190 2190.040 ;
        RECT 26.290 2189.980 26.610 2190.040 ;
      LAYER via ;
        RECT 13.900 2189.980 14.160 2190.240 ;
        RECT 26.320 2189.980 26.580 2190.240 ;
      LAYER met2 ;
        RECT 2285.830 3196.410 2286.110 3196.525 ;
        RECT 2286.680 3196.410 2286.960 3200.000 ;
        RECT 2285.830 3196.270 2286.960 3196.410 ;
        RECT 2285.830 3196.155 2286.110 3196.270 ;
        RECT 2286.680 3196.000 2286.960 3196.270 ;
        RECT 26.310 3193.435 26.590 3193.805 ;
        RECT 26.380 2190.270 26.520 3193.435 ;
        RECT 13.900 2190.125 14.160 2190.270 ;
        RECT 13.890 2189.755 14.170 2190.125 ;
        RECT 26.320 2189.950 26.580 2190.270 ;
      LAYER via2 ;
        RECT 2285.830 3196.200 2286.110 3196.480 ;
        RECT 26.310 3193.480 26.590 3193.760 ;
        RECT 13.890 2189.800 14.170 2190.080 ;
      LAYER met3 ;
        RECT 2088.670 3197.850 2089.050 3197.860 ;
        RECT 2113.510 3197.850 2113.890 3197.860 ;
        RECT 2088.670 3197.550 2113.890 3197.850 ;
        RECT 2088.670 3197.540 2089.050 3197.550 ;
        RECT 2113.510 3197.540 2113.890 3197.550 ;
        RECT 1810.830 3196.490 1811.210 3196.500 ;
        RECT 1825.550 3196.490 1825.930 3196.500 ;
        RECT 2285.805 3196.490 2286.135 3196.505 ;
        RECT 1810.830 3196.190 1825.930 3196.490 ;
        RECT 1810.830 3196.180 1811.210 3196.190 ;
        RECT 1825.550 3196.180 1825.930 3196.190 ;
        RECT 2285.590 3196.175 2286.135 3196.490 ;
        RECT 2186.190 3195.130 2186.570 3195.140 ;
        RECT 2282.790 3195.130 2283.170 3195.140 ;
        RECT 2285.590 3195.130 2285.890 3196.175 ;
        RECT 2186.190 3194.830 2188.370 3195.130 ;
        RECT 2186.190 3194.820 2186.570 3194.830 ;
        RECT 26.285 3193.770 26.615 3193.785 ;
        RECT 1776.790 3193.770 1777.170 3193.780 ;
        RECT 1810.830 3193.770 1811.210 3193.780 ;
        RECT 26.285 3193.470 1678.690 3193.770 ;
        RECT 26.285 3193.455 26.615 3193.470 ;
        RECT 1678.390 3192.410 1678.690 3193.470 ;
        RECT 1776.790 3193.470 1811.210 3193.770 ;
        RECT 1776.790 3193.460 1777.170 3193.470 ;
        RECT 1810.830 3193.460 1811.210 3193.470 ;
        RECT 1873.390 3193.770 1873.770 3193.780 ;
        RECT 1921.230 3193.770 1921.610 3193.780 ;
        RECT 1873.390 3193.470 1921.610 3193.770 ;
        RECT 1873.390 3193.460 1873.770 3193.470 ;
        RECT 1921.230 3193.460 1921.610 3193.470 ;
        RECT 2113.510 3193.770 2113.890 3193.780 ;
        RECT 2186.190 3193.770 2186.570 3193.780 ;
        RECT 2113.510 3193.470 2186.570 3193.770 ;
        RECT 2188.070 3193.770 2188.370 3194.830 ;
        RECT 2282.790 3194.830 2285.890 3195.130 ;
        RECT 2282.790 3194.820 2283.170 3194.830 ;
        RECT 2282.790 3193.770 2283.170 3193.780 ;
        RECT 2188.070 3193.470 2283.170 3193.770 ;
        RECT 2113.510 3193.460 2113.890 3193.470 ;
        RECT 2186.190 3193.460 2186.570 3193.470 ;
        RECT 2282.790 3193.460 2283.170 3193.470 ;
        RECT 1776.790 3192.410 1777.170 3192.420 ;
        RECT 1678.390 3192.110 1777.170 3192.410 ;
        RECT 1776.790 3192.100 1777.170 3192.110 ;
        RECT 1825.550 3192.410 1825.930 3192.420 ;
        RECT 1873.390 3192.410 1873.770 3192.420 ;
        RECT 1825.550 3192.110 1873.770 3192.410 ;
        RECT 1825.550 3192.100 1825.930 3192.110 ;
        RECT 1873.390 3192.100 1873.770 3192.110 ;
        RECT 1921.230 3192.410 1921.610 3192.420 ;
        RECT 2088.670 3192.410 2089.050 3192.420 ;
        RECT 1921.230 3192.110 2089.050 3192.410 ;
        RECT 1921.230 3192.100 1921.610 3192.110 ;
        RECT 2088.670 3192.100 2089.050 3192.110 ;
        RECT -4.800 2190.090 2.400 2190.540 ;
        RECT 13.865 2190.090 14.195 2190.105 ;
        RECT -4.800 2189.790 14.195 2190.090 ;
        RECT -4.800 2189.340 2.400 2189.790 ;
        RECT 13.865 2189.775 14.195 2189.790 ;
      LAYER via3 ;
        RECT 2088.700 3197.540 2089.020 3197.860 ;
        RECT 2113.540 3197.540 2113.860 3197.860 ;
        RECT 1810.860 3196.180 1811.180 3196.500 ;
        RECT 1825.580 3196.180 1825.900 3196.500 ;
        RECT 2186.220 3194.820 2186.540 3195.140 ;
        RECT 1776.820 3193.460 1777.140 3193.780 ;
        RECT 1810.860 3193.460 1811.180 3193.780 ;
        RECT 1873.420 3193.460 1873.740 3193.780 ;
        RECT 1921.260 3193.460 1921.580 3193.780 ;
        RECT 2113.540 3193.460 2113.860 3193.780 ;
        RECT 2186.220 3193.460 2186.540 3193.780 ;
        RECT 2282.820 3194.820 2283.140 3195.140 ;
        RECT 2282.820 3193.460 2283.140 3193.780 ;
        RECT 1776.820 3192.100 1777.140 3192.420 ;
        RECT 1825.580 3192.100 1825.900 3192.420 ;
        RECT 1873.420 3192.100 1873.740 3192.420 ;
        RECT 1921.260 3192.100 1921.580 3192.420 ;
        RECT 2088.700 3192.100 2089.020 3192.420 ;
      LAYER met4 ;
        RECT 2088.695 3197.535 2089.025 3197.865 ;
        RECT 2113.535 3197.535 2113.865 3197.865 ;
        RECT 1810.855 3196.175 1811.185 3196.505 ;
        RECT 1825.575 3196.175 1825.905 3196.505 ;
        RECT 1810.870 3193.785 1811.170 3196.175 ;
        RECT 1776.815 3193.455 1777.145 3193.785 ;
        RECT 1810.855 3193.455 1811.185 3193.785 ;
        RECT 1776.830 3192.425 1777.130 3193.455 ;
        RECT 1825.590 3192.425 1825.890 3196.175 ;
        RECT 1873.415 3193.455 1873.745 3193.785 ;
        RECT 1921.255 3193.455 1921.585 3193.785 ;
        RECT 1873.430 3192.425 1873.730 3193.455 ;
        RECT 1921.270 3192.425 1921.570 3193.455 ;
        RECT 2088.710 3192.425 2089.010 3197.535 ;
        RECT 2113.550 3193.785 2113.850 3197.535 ;
        RECT 2186.215 3194.815 2186.545 3195.145 ;
        RECT 2282.815 3194.815 2283.145 3195.145 ;
        RECT 2186.230 3193.785 2186.530 3194.815 ;
        RECT 2282.830 3193.785 2283.130 3194.815 ;
        RECT 2113.535 3193.455 2113.865 3193.785 ;
        RECT 2186.215 3193.455 2186.545 3193.785 ;
        RECT 2282.815 3193.455 2283.145 3193.785 ;
        RECT 1776.815 3192.095 1777.145 3192.425 ;
        RECT 1825.575 3192.095 1825.905 3192.425 ;
        RECT 1873.415 3192.095 1873.745 3192.425 ;
        RECT 1921.255 3192.095 1921.585 3192.425 ;
        RECT 2088.695 3192.095 2089.025 3192.425 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 31.810 3210.860 32.130 3210.920 ;
        RECT 2325.830 3210.860 2326.150 3210.920 ;
        RECT 31.810 3210.720 2326.150 3210.860 ;
        RECT 31.810 3210.660 32.130 3210.720 ;
        RECT 2325.830 3210.660 2326.150 3210.720 ;
        RECT 16.170 1903.220 16.490 1903.280 ;
        RECT 31.810 1903.220 32.130 1903.280 ;
        RECT 16.170 1903.080 32.130 1903.220 ;
        RECT 16.170 1903.020 16.490 1903.080 ;
        RECT 31.810 1903.020 32.130 1903.080 ;
      LAYER via ;
        RECT 31.840 3210.660 32.100 3210.920 ;
        RECT 2325.860 3210.660 2326.120 3210.920 ;
        RECT 16.200 1903.020 16.460 1903.280 ;
        RECT 31.840 1903.020 32.100 1903.280 ;
      LAYER met2 ;
        RECT 31.840 3210.630 32.100 3210.950 ;
        RECT 2325.860 3210.630 2326.120 3210.950 ;
        RECT 31.900 1903.310 32.040 3210.630 ;
        RECT 2325.920 3200.000 2326.060 3210.630 ;
        RECT 2325.780 3196.000 2326.060 3200.000 ;
        RECT 16.200 1903.165 16.460 1903.310 ;
        RECT 16.190 1902.795 16.470 1903.165 ;
        RECT 31.840 1902.990 32.100 1903.310 ;
      LAYER via2 ;
        RECT 16.190 1902.840 16.470 1903.120 ;
      LAYER met3 ;
        RECT -4.800 1903.130 2.400 1903.580 ;
        RECT 16.165 1903.130 16.495 1903.145 ;
        RECT -4.800 1902.830 16.495 1903.130 ;
        RECT -4.800 1902.380 2.400 1902.830 ;
        RECT 16.165 1902.815 16.495 1902.830 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1729.670 616.320 1729.990 616.380 ;
        RECT 1772.910 616.320 1773.230 616.380 ;
        RECT 1729.670 616.180 1773.230 616.320 ;
        RECT 1729.670 616.120 1729.990 616.180 ;
        RECT 1772.910 616.120 1773.230 616.180 ;
        RECT 2270.170 615.300 2270.490 615.360 ;
        RECT 2290.870 615.300 2291.190 615.360 ;
        RECT 2270.170 615.160 2291.190 615.300 ;
        RECT 2270.170 615.100 2270.490 615.160 ;
        RECT 2290.870 615.100 2291.190 615.160 ;
        RECT 2572.850 615.300 2573.170 615.360 ;
        RECT 2584.350 615.300 2584.670 615.360 ;
        RECT 2572.850 615.160 2584.670 615.300 ;
        RECT 2572.850 615.100 2573.170 615.160 ;
        RECT 2584.350 615.100 2584.670 615.160 ;
        RECT 2379.650 614.960 2379.970 615.020 ;
        RECT 2390.690 614.960 2391.010 615.020 ;
        RECT 2379.650 614.820 2391.010 614.960 ;
        RECT 2379.650 614.760 2379.970 614.820 ;
        RECT 2390.690 614.760 2391.010 614.820 ;
        RECT 2125.270 614.620 2125.590 614.680 ;
        RECT 2172.650 614.620 2172.970 614.680 ;
        RECT 2125.270 614.480 2172.970 614.620 ;
        RECT 2125.270 614.420 2125.590 614.480 ;
        RECT 2172.650 614.420 2172.970 614.480 ;
        RECT 2621.150 614.620 2621.470 614.680 ;
        RECT 2632.190 614.620 2632.510 614.680 ;
        RECT 2621.150 614.480 2632.510 614.620 ;
        RECT 2621.150 614.420 2621.470 614.480 ;
        RECT 2632.190 614.420 2632.510 614.480 ;
      LAYER via ;
        RECT 1729.700 616.120 1729.960 616.380 ;
        RECT 1772.940 616.120 1773.200 616.380 ;
        RECT 2270.200 615.100 2270.460 615.360 ;
        RECT 2290.900 615.100 2291.160 615.360 ;
        RECT 2572.880 615.100 2573.140 615.360 ;
        RECT 2584.380 615.100 2584.640 615.360 ;
        RECT 2379.680 614.760 2379.940 615.020 ;
        RECT 2390.720 614.760 2390.980 615.020 ;
        RECT 2125.300 614.420 2125.560 614.680 ;
        RECT 2172.680 614.420 2172.940 614.680 ;
        RECT 2621.180 614.420 2621.440 614.680 ;
        RECT 2632.220 614.420 2632.480 614.680 ;
      LAYER met2 ;
        RECT 1259.960 3196.410 1260.240 3200.000 ;
        RECT 1261.410 3196.410 1261.690 3196.525 ;
        RECT 1259.960 3196.270 1261.690 3196.410 ;
        RECT 1259.960 3196.000 1260.240 3196.270 ;
        RECT 1261.410 3196.155 1261.690 3196.270 ;
        RECT 1724.630 616.235 1724.910 616.605 ;
        RECT 1729.690 616.235 1729.970 616.605 ;
        RECT 1724.700 614.565 1724.840 616.235 ;
        RECT 1729.700 616.090 1729.960 616.235 ;
        RECT 1772.940 616.090 1773.200 616.410 ;
        RECT 2704.430 616.235 2704.710 616.605 ;
        RECT 1773.000 615.925 1773.140 616.090 ;
        RECT 1772.930 615.555 1773.210 615.925 ;
        RECT 2172.670 615.555 2172.950 615.925 ;
        RECT 2172.740 614.710 2172.880 615.555 ;
        RECT 2270.200 615.245 2270.460 615.390 ;
        RECT 2290.900 615.245 2291.160 615.390 ;
        RECT 2572.880 615.245 2573.140 615.390 ;
        RECT 2584.380 615.245 2584.640 615.390 ;
        RECT 2270.190 614.875 2270.470 615.245 ;
        RECT 2290.890 614.875 2291.170 615.245 ;
        RECT 2379.670 614.875 2379.950 615.245 ;
        RECT 2390.710 614.875 2390.990 615.245 ;
        RECT 2572.870 614.875 2573.150 615.245 ;
        RECT 2584.370 614.875 2584.650 615.245 ;
        RECT 2632.210 614.875 2632.490 615.245 ;
        RECT 2379.680 614.730 2379.940 614.875 ;
        RECT 2390.720 614.730 2390.980 614.875 ;
        RECT 2632.280 614.710 2632.420 614.875 ;
        RECT 2125.300 614.565 2125.560 614.710 ;
        RECT 1724.630 614.195 1724.910 614.565 ;
        RECT 2125.290 614.195 2125.570 614.565 ;
        RECT 2172.680 614.390 2172.940 614.710 ;
        RECT 2621.180 614.565 2621.440 614.710 ;
        RECT 2621.170 614.195 2621.450 614.565 ;
        RECT 2632.220 614.390 2632.480 614.710 ;
        RECT 2704.500 614.565 2704.640 616.235 ;
        RECT 2801.030 615.555 2801.310 615.925 ;
        RECT 2704.430 614.195 2704.710 614.565 ;
        RECT 2801.100 613.885 2801.240 615.555 ;
        RECT 2863.130 614.875 2863.410 615.245 ;
        RECT 2863.200 614.450 2863.340 614.875 ;
        RECT 2863.590 614.450 2863.870 614.565 ;
        RECT 2863.200 614.310 2863.870 614.450 ;
        RECT 2863.590 614.195 2863.870 614.310 ;
        RECT 2801.030 613.515 2801.310 613.885 ;
      LAYER via2 ;
        RECT 1261.410 3196.200 1261.690 3196.480 ;
        RECT 1724.630 616.280 1724.910 616.560 ;
        RECT 1729.690 616.280 1729.970 616.560 ;
        RECT 2704.430 616.280 2704.710 616.560 ;
        RECT 1772.930 615.600 1773.210 615.880 ;
        RECT 2172.670 615.600 2172.950 615.880 ;
        RECT 2270.190 614.920 2270.470 615.200 ;
        RECT 2290.890 614.920 2291.170 615.200 ;
        RECT 2379.670 614.920 2379.950 615.200 ;
        RECT 2390.710 614.920 2390.990 615.200 ;
        RECT 2572.870 614.920 2573.150 615.200 ;
        RECT 2584.370 614.920 2584.650 615.200 ;
        RECT 2632.210 614.920 2632.490 615.200 ;
        RECT 1724.630 614.240 1724.910 614.520 ;
        RECT 2125.290 614.240 2125.570 614.520 ;
        RECT 2621.170 614.240 2621.450 614.520 ;
        RECT 2801.030 615.600 2801.310 615.880 ;
        RECT 2704.430 614.240 2704.710 614.520 ;
        RECT 2863.130 614.920 2863.410 615.200 ;
        RECT 2863.590 614.240 2863.870 614.520 ;
        RECT 2801.030 613.560 2801.310 613.840 ;
      LAYER met3 ;
        RECT 1261.385 3196.500 1261.715 3196.505 ;
        RECT 1261.385 3196.490 1261.970 3196.500 ;
        RECT 1261.385 3196.190 1262.170 3196.490 ;
        RECT 1261.385 3196.180 1261.970 3196.190 ;
        RECT 1261.385 3196.175 1261.715 3196.180 ;
        RECT 1828.310 617.250 1828.690 617.260 ;
        RECT 1828.310 616.950 1876.490 617.250 ;
        RECT 1828.310 616.940 1828.690 616.950 ;
        RECT 1538.510 616.570 1538.890 616.580 ;
        RECT 1724.605 616.570 1724.935 616.585 ;
        RECT 1729.665 616.570 1729.995 616.585 ;
        RECT 1538.510 616.270 1611.530 616.570 ;
        RECT 1538.510 616.260 1538.890 616.270 ;
        RECT 1261.590 615.890 1261.970 615.900 ;
        RECT 1611.230 615.890 1611.530 616.270 ;
        RECT 1724.605 616.270 1729.995 616.570 ;
        RECT 1876.190 616.570 1876.490 616.950 ;
        RECT 2656.310 616.570 2656.690 616.580 ;
        RECT 2704.405 616.570 2704.735 616.585 ;
        RECT 1876.190 616.270 1898.570 616.570 ;
        RECT 1724.605 616.255 1724.935 616.270 ;
        RECT 1729.665 616.255 1729.995 616.270 ;
        RECT 1676.510 615.890 1676.890 615.900 ;
        RECT 1261.590 615.590 1393.490 615.890 ;
        RECT 1261.590 615.580 1261.970 615.590 ;
        RECT 1393.190 615.210 1393.490 615.590 ;
        RECT 1462.190 615.590 1510.330 615.890 ;
        RECT 1611.230 615.590 1676.890 615.890 ;
        RECT 1462.190 615.210 1462.490 615.590 ;
        RECT 1393.190 614.910 1462.490 615.210 ;
        RECT 1510.030 615.210 1510.330 615.590 ;
        RECT 1676.510 615.580 1676.890 615.590 ;
        RECT 1772.905 615.890 1773.235 615.905 ;
        RECT 1772.905 615.590 1804.730 615.890 ;
        RECT 1772.905 615.575 1773.235 615.590 ;
        RECT 1538.510 615.210 1538.890 615.220 ;
        RECT 1510.030 614.910 1538.890 615.210 ;
        RECT 1804.430 615.210 1804.730 615.590 ;
        RECT 1828.310 615.210 1828.690 615.220 ;
        RECT 1804.430 614.910 1828.690 615.210 ;
        RECT 1898.270 615.210 1898.570 616.270 ;
        RECT 2476.030 616.270 2511.290 616.570 ;
        RECT 2172.645 615.890 2172.975 615.905 ;
        RECT 1970.030 615.590 1994.250 615.890 ;
        RECT 1970.030 615.210 1970.330 615.590 ;
        RECT 1898.270 614.910 1970.330 615.210 ;
        RECT 1538.510 614.900 1538.890 614.910 ;
        RECT 1828.310 614.900 1828.690 614.910 ;
        RECT 1676.510 614.530 1676.890 614.540 ;
        RECT 1724.605 614.530 1724.935 614.545 ;
        RECT 1676.510 614.230 1724.935 614.530 ;
        RECT 1993.950 614.530 1994.250 615.590 ;
        RECT 2172.645 615.590 2187.450 615.890 ;
        RECT 2172.645 615.575 2172.975 615.590 ;
        RECT 2042.710 614.910 2090.850 615.210 ;
        RECT 2042.710 614.530 2043.010 614.910 ;
        RECT 1993.950 614.230 2043.010 614.530 ;
        RECT 2090.550 614.530 2090.850 614.910 ;
        RECT 2125.265 614.530 2125.595 614.545 ;
        RECT 2090.550 614.230 2125.595 614.530 ;
        RECT 2187.150 614.530 2187.450 615.590 ;
        RECT 2270.165 615.210 2270.495 615.225 ;
        RECT 2235.910 614.910 2270.495 615.210 ;
        RECT 2235.910 614.530 2236.210 614.910 ;
        RECT 2270.165 614.895 2270.495 614.910 ;
        RECT 2290.865 615.210 2291.195 615.225 ;
        RECT 2379.645 615.210 2379.975 615.225 ;
        RECT 2290.865 614.910 2318.090 615.210 ;
        RECT 2290.865 614.895 2291.195 614.910 ;
        RECT 2187.150 614.230 2236.210 614.530 ;
        RECT 2317.790 614.530 2318.090 614.910 ;
        RECT 2332.510 614.910 2379.975 615.210 ;
        RECT 2332.510 614.530 2332.810 614.910 ;
        RECT 2379.645 614.895 2379.975 614.910 ;
        RECT 2390.685 615.210 2391.015 615.225 ;
        RECT 2476.030 615.210 2476.330 616.270 ;
        RECT 2390.685 614.910 2414.690 615.210 ;
        RECT 2390.685 614.895 2391.015 614.910 ;
        RECT 2317.790 614.230 2332.810 614.530 ;
        RECT 2414.390 614.530 2414.690 614.910 ;
        RECT 2429.110 614.910 2476.330 615.210 ;
        RECT 2429.110 614.530 2429.410 614.910 ;
        RECT 2414.390 614.230 2429.410 614.530 ;
        RECT 2510.990 614.530 2511.290 616.270 ;
        RECT 2656.310 616.270 2704.735 616.570 ;
        RECT 2656.310 616.260 2656.690 616.270 ;
        RECT 2704.405 616.255 2704.735 616.270 ;
        RECT 2801.005 615.890 2801.335 615.905 ;
        RECT 2917.600 615.890 2924.800 616.340 ;
        RECT 2801.005 615.590 2815.810 615.890 ;
        RECT 2801.005 615.575 2801.335 615.590 ;
        RECT 2572.845 615.210 2573.175 615.225 ;
        RECT 2525.710 614.910 2573.175 615.210 ;
        RECT 2525.710 614.530 2526.010 614.910 ;
        RECT 2572.845 614.895 2573.175 614.910 ;
        RECT 2584.345 615.210 2584.675 615.225 ;
        RECT 2632.185 615.210 2632.515 615.225 ;
        RECT 2656.310 615.210 2656.690 615.220 ;
        RECT 2752.910 615.210 2753.290 615.220 ;
        RECT 2584.345 614.910 2607.890 615.210 ;
        RECT 2584.345 614.895 2584.675 614.910 ;
        RECT 2510.990 614.230 2526.010 614.530 ;
        RECT 2607.590 614.530 2607.890 614.910 ;
        RECT 2632.185 614.910 2656.690 615.210 ;
        RECT 2632.185 614.895 2632.515 614.910 ;
        RECT 2656.310 614.900 2656.690 614.910 ;
        RECT 2718.910 614.910 2753.290 615.210 ;
        RECT 2621.145 614.530 2621.475 614.545 ;
        RECT 2607.590 614.230 2621.475 614.530 ;
        RECT 1676.510 614.220 1676.890 614.230 ;
        RECT 1724.605 614.215 1724.935 614.230 ;
        RECT 2125.265 614.215 2125.595 614.230 ;
        RECT 2621.145 614.215 2621.475 614.230 ;
        RECT 2704.405 614.530 2704.735 614.545 ;
        RECT 2718.910 614.530 2719.210 614.910 ;
        RECT 2752.910 614.900 2753.290 614.910 ;
        RECT 2704.405 614.230 2719.210 614.530 ;
        RECT 2815.510 614.530 2815.810 615.590 ;
        RECT 2916.710 615.590 2924.800 615.890 ;
        RECT 2863.105 615.210 2863.435 615.225 ;
        RECT 2916.710 615.210 2917.010 615.590 ;
        RECT 2849.550 614.910 2863.435 615.210 ;
        RECT 2849.550 614.530 2849.850 614.910 ;
        RECT 2863.105 614.895 2863.435 614.910 ;
        RECT 2884.510 614.910 2917.010 615.210 ;
        RECT 2917.600 615.140 2924.800 615.590 ;
        RECT 2815.510 614.230 2849.850 614.530 ;
        RECT 2863.565 614.530 2863.895 614.545 ;
        RECT 2884.510 614.530 2884.810 614.910 ;
        RECT 2863.565 614.230 2884.810 614.530 ;
        RECT 2704.405 614.215 2704.735 614.230 ;
        RECT 2863.565 614.215 2863.895 614.230 ;
        RECT 2752.910 613.850 2753.290 613.860 ;
        RECT 2801.005 613.850 2801.335 613.865 ;
        RECT 2752.910 613.550 2801.335 613.850 ;
        RECT 2752.910 613.540 2753.290 613.550 ;
        RECT 2801.005 613.535 2801.335 613.550 ;
      LAYER via3 ;
        RECT 1261.620 3196.180 1261.940 3196.500 ;
        RECT 1828.340 616.940 1828.660 617.260 ;
        RECT 1538.540 616.260 1538.860 616.580 ;
        RECT 1261.620 615.580 1261.940 615.900 ;
        RECT 1676.540 615.580 1676.860 615.900 ;
        RECT 1538.540 614.900 1538.860 615.220 ;
        RECT 1828.340 614.900 1828.660 615.220 ;
        RECT 1676.540 614.220 1676.860 614.540 ;
        RECT 2656.340 616.260 2656.660 616.580 ;
        RECT 2656.340 614.900 2656.660 615.220 ;
        RECT 2752.940 614.900 2753.260 615.220 ;
        RECT 2752.940 613.540 2753.260 613.860 ;
      LAYER met4 ;
        RECT 1261.615 3196.175 1261.945 3196.505 ;
        RECT 1261.630 615.905 1261.930 3196.175 ;
        RECT 1828.335 616.935 1828.665 617.265 ;
        RECT 1538.535 616.255 1538.865 616.585 ;
        RECT 1261.615 615.575 1261.945 615.905 ;
        RECT 1538.550 615.225 1538.850 616.255 ;
        RECT 1676.535 615.575 1676.865 615.905 ;
        RECT 1538.535 614.895 1538.865 615.225 ;
        RECT 1676.550 614.545 1676.850 615.575 ;
        RECT 1828.350 615.225 1828.650 616.935 ;
        RECT 2656.335 616.255 2656.665 616.585 ;
        RECT 2656.350 615.225 2656.650 616.255 ;
        RECT 1828.335 614.895 1828.665 615.225 ;
        RECT 2656.335 614.895 2656.665 615.225 ;
        RECT 2752.935 614.895 2753.265 615.225 ;
        RECT 1676.535 614.215 1676.865 614.545 ;
        RECT 2752.950 613.865 2753.250 614.895 ;
        RECT 2752.935 613.535 2753.265 613.865 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2365.410 3213.155 2365.690 3213.525 ;
        RECT 2365.480 3200.000 2365.620 3213.155 ;
        RECT 2365.340 3196.000 2365.620 3200.000 ;
        RECT 15.730 1621.275 16.010 1621.645 ;
        RECT 15.800 1615.525 15.940 1621.275 ;
        RECT 15.730 1615.155 16.010 1615.525 ;
      LAYER via2 ;
        RECT 2365.410 3213.200 2365.690 3213.480 ;
        RECT 15.730 1621.320 16.010 1621.600 ;
        RECT 15.730 1615.200 16.010 1615.480 ;
      LAYER met3 ;
        RECT 1294.710 3213.490 1295.090 3213.500 ;
        RECT 2365.385 3213.490 2365.715 3213.505 ;
        RECT 1294.710 3213.190 2365.715 3213.490 ;
        RECT 1294.710 3213.180 1295.090 3213.190 ;
        RECT 2365.385 3213.175 2365.715 3213.190 ;
        RECT 15.705 1621.610 16.035 1621.625 ;
        RECT 1294.710 1621.610 1295.090 1621.620 ;
        RECT 15.705 1621.310 1295.090 1621.610 ;
        RECT 15.705 1621.295 16.035 1621.310 ;
        RECT 1294.710 1621.300 1295.090 1621.310 ;
        RECT -4.800 1615.490 2.400 1615.940 ;
        RECT 15.705 1615.490 16.035 1615.505 ;
        RECT -4.800 1615.190 16.035 1615.490 ;
        RECT -4.800 1614.740 2.400 1615.190 ;
        RECT 15.705 1615.175 16.035 1615.190 ;
      LAYER via3 ;
        RECT 1294.740 3213.180 1295.060 3213.500 ;
        RECT 1294.740 1621.300 1295.060 1621.620 ;
      LAYER met4 ;
        RECT 1294.735 3213.175 1295.065 3213.505 ;
        RECT 1294.750 1621.625 1295.050 3213.175 ;
        RECT 1294.735 1621.295 1295.065 1621.625 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 31.350 3210.180 31.670 3210.240 ;
        RECT 2404.950 3210.180 2405.270 3210.240 ;
        RECT 31.350 3210.040 2405.270 3210.180 ;
        RECT 31.350 3209.980 31.670 3210.040 ;
        RECT 2404.950 3209.980 2405.270 3210.040 ;
        RECT 15.710 1400.700 16.030 1400.760 ;
        RECT 31.350 1400.700 31.670 1400.760 ;
        RECT 15.710 1400.560 31.670 1400.700 ;
        RECT 15.710 1400.500 16.030 1400.560 ;
        RECT 31.350 1400.500 31.670 1400.560 ;
      LAYER via ;
        RECT 31.380 3209.980 31.640 3210.240 ;
        RECT 2404.980 3209.980 2405.240 3210.240 ;
        RECT 15.740 1400.500 16.000 1400.760 ;
        RECT 31.380 1400.500 31.640 1400.760 ;
      LAYER met2 ;
        RECT 31.380 3209.950 31.640 3210.270 ;
        RECT 2404.980 3209.950 2405.240 3210.270 ;
        RECT 31.440 1400.790 31.580 3209.950 ;
        RECT 2405.040 3200.000 2405.180 3209.950 ;
        RECT 2404.900 3196.000 2405.180 3200.000 ;
        RECT 15.740 1400.645 16.000 1400.790 ;
        RECT 15.730 1400.275 16.010 1400.645 ;
        RECT 31.380 1400.470 31.640 1400.790 ;
      LAYER via2 ;
        RECT 15.730 1400.320 16.010 1400.600 ;
      LAYER met3 ;
        RECT -4.800 1400.610 2.400 1401.060 ;
        RECT 15.705 1400.610 16.035 1400.625 ;
        RECT -4.800 1400.310 16.035 1400.610 ;
        RECT -4.800 1399.860 2.400 1400.310 ;
        RECT 15.705 1400.295 16.035 1400.310 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 13.870 1185.820 14.190 1185.880 ;
        RECT 24.450 1185.820 24.770 1185.880 ;
        RECT 13.870 1185.680 24.770 1185.820 ;
        RECT 13.870 1185.620 14.190 1185.680 ;
        RECT 24.450 1185.620 24.770 1185.680 ;
      LAYER via ;
        RECT 13.900 1185.620 14.160 1185.880 ;
        RECT 24.480 1185.620 24.740 1185.880 ;
      LAYER met2 ;
        RECT 2443.150 3196.410 2443.430 3196.525 ;
        RECT 2444.460 3196.410 2444.740 3200.000 ;
        RECT 2443.150 3196.270 2444.740 3196.410 ;
        RECT 2443.150 3196.155 2443.430 3196.270 ;
        RECT 2444.460 3196.000 2444.740 3196.270 ;
        RECT 24.470 3192.075 24.750 3192.445 ;
        RECT 34.590 3192.075 34.870 3192.445 ;
        RECT 86.110 3192.075 86.390 3192.445 ;
        RECT 131.190 3192.330 131.470 3192.445 ;
        RECT 131.190 3192.190 131.860 3192.330 ;
        RECT 131.190 3192.075 131.470 3192.190 ;
        RECT 24.540 1185.910 24.680 3192.075 ;
        RECT 34.660 3190.405 34.800 3192.075 ;
        RECT 86.180 3190.405 86.320 3192.075 ;
        RECT 131.720 3190.405 131.860 3192.190 ;
        RECT 182.710 3192.075 182.990 3192.445 ;
        RECT 227.790 3192.330 228.070 3192.445 ;
        RECT 227.790 3192.190 228.460 3192.330 ;
        RECT 227.790 3192.075 228.070 3192.190 ;
        RECT 182.780 3190.405 182.920 3192.075 ;
        RECT 228.320 3190.405 228.460 3192.190 ;
        RECT 279.310 3192.075 279.590 3192.445 ;
        RECT 324.390 3192.330 324.670 3192.445 ;
        RECT 324.390 3192.190 325.060 3192.330 ;
        RECT 324.390 3192.075 324.670 3192.190 ;
        RECT 279.380 3190.405 279.520 3192.075 ;
        RECT 324.920 3190.405 325.060 3192.190 ;
        RECT 375.910 3192.075 376.190 3192.445 ;
        RECT 420.990 3192.330 421.270 3192.445 ;
        RECT 420.990 3192.190 421.660 3192.330 ;
        RECT 420.990 3192.075 421.270 3192.190 ;
        RECT 375.980 3190.405 376.120 3192.075 ;
        RECT 421.520 3190.405 421.660 3192.190 ;
        RECT 472.510 3192.075 472.790 3192.445 ;
        RECT 517.590 3192.330 517.870 3192.445 ;
        RECT 517.590 3192.190 518.260 3192.330 ;
        RECT 517.590 3192.075 517.870 3192.190 ;
        RECT 472.580 3190.405 472.720 3192.075 ;
        RECT 518.120 3190.405 518.260 3192.190 ;
        RECT 569.110 3192.075 569.390 3192.445 ;
        RECT 614.190 3192.330 614.470 3192.445 ;
        RECT 614.190 3192.190 614.860 3192.330 ;
        RECT 614.190 3192.075 614.470 3192.190 ;
        RECT 569.180 3190.405 569.320 3192.075 ;
        RECT 614.720 3190.405 614.860 3192.190 ;
        RECT 665.710 3192.075 665.990 3192.445 ;
        RECT 710.790 3192.330 711.070 3192.445 ;
        RECT 710.790 3192.190 711.460 3192.330 ;
        RECT 710.790 3192.075 711.070 3192.190 ;
        RECT 665.780 3190.405 665.920 3192.075 ;
        RECT 711.320 3190.405 711.460 3192.190 ;
        RECT 762.310 3192.075 762.590 3192.445 ;
        RECT 807.390 3192.330 807.670 3192.445 ;
        RECT 807.390 3192.190 808.060 3192.330 ;
        RECT 807.390 3192.075 807.670 3192.190 ;
        RECT 762.380 3190.405 762.520 3192.075 ;
        RECT 807.920 3190.405 808.060 3192.190 ;
        RECT 858.910 3192.075 859.190 3192.445 ;
        RECT 903.990 3192.330 904.270 3192.445 ;
        RECT 903.990 3192.190 904.660 3192.330 ;
        RECT 903.990 3192.075 904.270 3192.190 ;
        RECT 858.980 3190.405 859.120 3192.075 ;
        RECT 904.520 3190.405 904.660 3192.190 ;
        RECT 955.510 3192.075 955.790 3192.445 ;
        RECT 1000.590 3192.330 1000.870 3192.445 ;
        RECT 1000.590 3192.190 1001.260 3192.330 ;
        RECT 1000.590 3192.075 1000.870 3192.190 ;
        RECT 955.580 3190.405 955.720 3192.075 ;
        RECT 1001.120 3190.405 1001.260 3192.190 ;
        RECT 1052.110 3192.075 1052.390 3192.445 ;
        RECT 1100.410 3192.075 1100.690 3192.445 ;
        RECT 1052.180 3190.405 1052.320 3192.075 ;
        RECT 34.590 3190.035 34.870 3190.405 ;
        RECT 86.110 3190.035 86.390 3190.405 ;
        RECT 131.650 3190.035 131.930 3190.405 ;
        RECT 182.710 3190.035 182.990 3190.405 ;
        RECT 228.250 3190.035 228.530 3190.405 ;
        RECT 279.310 3190.035 279.590 3190.405 ;
        RECT 324.850 3190.035 325.130 3190.405 ;
        RECT 375.910 3190.035 376.190 3190.405 ;
        RECT 421.450 3190.035 421.730 3190.405 ;
        RECT 472.510 3190.035 472.790 3190.405 ;
        RECT 518.050 3190.035 518.330 3190.405 ;
        RECT 569.110 3190.035 569.390 3190.405 ;
        RECT 614.650 3190.035 614.930 3190.405 ;
        RECT 665.710 3190.035 665.990 3190.405 ;
        RECT 711.250 3190.035 711.530 3190.405 ;
        RECT 762.310 3190.035 762.590 3190.405 ;
        RECT 807.850 3190.035 808.130 3190.405 ;
        RECT 858.910 3190.035 859.190 3190.405 ;
        RECT 904.450 3190.035 904.730 3190.405 ;
        RECT 955.510 3190.035 955.790 3190.405 ;
        RECT 1001.050 3190.035 1001.330 3190.405 ;
        RECT 1052.110 3190.035 1052.390 3190.405 ;
        RECT 1100.480 3189.725 1100.620 3192.075 ;
        RECT 1100.410 3189.355 1100.690 3189.725 ;
        RECT 13.900 1185.590 14.160 1185.910 ;
        RECT 24.480 1185.590 24.740 1185.910 ;
        RECT 13.960 1185.085 14.100 1185.590 ;
        RECT 13.890 1184.715 14.170 1185.085 ;
      LAYER via2 ;
        RECT 2443.150 3196.200 2443.430 3196.480 ;
        RECT 24.470 3192.120 24.750 3192.400 ;
        RECT 34.590 3192.120 34.870 3192.400 ;
        RECT 86.110 3192.120 86.390 3192.400 ;
        RECT 131.190 3192.120 131.470 3192.400 ;
        RECT 182.710 3192.120 182.990 3192.400 ;
        RECT 227.790 3192.120 228.070 3192.400 ;
        RECT 279.310 3192.120 279.590 3192.400 ;
        RECT 324.390 3192.120 324.670 3192.400 ;
        RECT 375.910 3192.120 376.190 3192.400 ;
        RECT 420.990 3192.120 421.270 3192.400 ;
        RECT 472.510 3192.120 472.790 3192.400 ;
        RECT 517.590 3192.120 517.870 3192.400 ;
        RECT 569.110 3192.120 569.390 3192.400 ;
        RECT 614.190 3192.120 614.470 3192.400 ;
        RECT 665.710 3192.120 665.990 3192.400 ;
        RECT 710.790 3192.120 711.070 3192.400 ;
        RECT 762.310 3192.120 762.590 3192.400 ;
        RECT 807.390 3192.120 807.670 3192.400 ;
        RECT 858.910 3192.120 859.190 3192.400 ;
        RECT 903.990 3192.120 904.270 3192.400 ;
        RECT 955.510 3192.120 955.790 3192.400 ;
        RECT 1000.590 3192.120 1000.870 3192.400 ;
        RECT 1052.110 3192.120 1052.390 3192.400 ;
        RECT 1100.410 3192.120 1100.690 3192.400 ;
        RECT 34.590 3190.080 34.870 3190.360 ;
        RECT 86.110 3190.080 86.390 3190.360 ;
        RECT 131.650 3190.080 131.930 3190.360 ;
        RECT 182.710 3190.080 182.990 3190.360 ;
        RECT 228.250 3190.080 228.530 3190.360 ;
        RECT 279.310 3190.080 279.590 3190.360 ;
        RECT 324.850 3190.080 325.130 3190.360 ;
        RECT 375.910 3190.080 376.190 3190.360 ;
        RECT 421.450 3190.080 421.730 3190.360 ;
        RECT 472.510 3190.080 472.790 3190.360 ;
        RECT 518.050 3190.080 518.330 3190.360 ;
        RECT 569.110 3190.080 569.390 3190.360 ;
        RECT 614.650 3190.080 614.930 3190.360 ;
        RECT 665.710 3190.080 665.990 3190.360 ;
        RECT 711.250 3190.080 711.530 3190.360 ;
        RECT 762.310 3190.080 762.590 3190.360 ;
        RECT 807.850 3190.080 808.130 3190.360 ;
        RECT 858.910 3190.080 859.190 3190.360 ;
        RECT 904.450 3190.080 904.730 3190.360 ;
        RECT 955.510 3190.080 955.790 3190.360 ;
        RECT 1001.050 3190.080 1001.330 3190.360 ;
        RECT 1052.110 3190.080 1052.390 3190.360 ;
        RECT 1100.410 3189.400 1100.690 3189.680 ;
        RECT 13.890 1184.760 14.170 1185.040 ;
      LAYER met3 ;
        RECT 2443.125 3196.500 2443.455 3196.505 ;
        RECT 2042.670 3196.490 2043.050 3196.500 ;
        RECT 2442.870 3196.490 2443.455 3196.500 ;
        RECT 2015.110 3196.190 2043.050 3196.490 ;
        RECT 2442.670 3196.190 2443.455 3196.490 ;
        RECT 1579.910 3195.810 1580.290 3195.820 ;
        RECT 1627.750 3195.810 1628.130 3195.820 ;
        RECT 1579.910 3195.510 1628.130 3195.810 ;
        RECT 1579.910 3195.500 1580.290 3195.510 ;
        RECT 1627.750 3195.500 1628.130 3195.510 ;
        RECT 1712.390 3195.810 1712.770 3195.820 ;
        RECT 1777.710 3195.810 1778.090 3195.820 ;
        RECT 1712.390 3195.510 1778.090 3195.810 ;
        RECT 1712.390 3195.500 1712.770 3195.510 ;
        RECT 1777.710 3195.500 1778.090 3195.510 ;
        RECT 1820.950 3195.810 1821.330 3195.820 ;
        RECT 1874.310 3195.810 1874.690 3195.820 ;
        RECT 1820.950 3195.510 1827.730 3195.810 ;
        RECT 1820.950 3195.500 1821.330 3195.510 ;
        RECT 1387.630 3195.130 1388.010 3195.140 ;
        RECT 1676.510 3195.130 1676.890 3195.140 ;
        RECT 1827.430 3195.130 1827.730 3195.510 ;
        RECT 1850.430 3195.510 1874.690 3195.810 ;
        RECT 1850.430 3195.130 1850.730 3195.510 ;
        RECT 1874.310 3195.500 1874.690 3195.510 ;
        RECT 1920.310 3195.810 1920.690 3195.820 ;
        RECT 1992.990 3195.810 1993.370 3195.820 ;
        RECT 1920.310 3195.510 1993.370 3195.810 ;
        RECT 1920.310 3195.500 1920.690 3195.510 ;
        RECT 1992.990 3195.500 1993.370 3195.510 ;
        RECT 1994.830 3195.810 1995.210 3195.820 ;
        RECT 2015.110 3195.810 2015.410 3196.190 ;
        RECT 2042.670 3196.180 2043.050 3196.190 ;
        RECT 2442.870 3196.180 2443.455 3196.190 ;
        RECT 2443.125 3196.175 2443.455 3196.180 ;
        RECT 1994.830 3195.510 2015.410 3195.810 ;
        RECT 1994.830 3195.500 1995.210 3195.510 ;
        RECT 1387.630 3194.830 1433.970 3195.130 ;
        RECT 1387.630 3194.820 1388.010 3194.830 ;
        RECT 1433.670 3194.460 1433.970 3194.830 ;
        RECT 1676.510 3194.830 1681.450 3195.130 ;
        RECT 1827.430 3194.830 1850.730 3195.130 ;
        RECT 2042.670 3195.130 2043.050 3195.140 ;
        RECT 2042.670 3194.830 2045.770 3195.130 ;
        RECT 1676.510 3194.820 1676.890 3194.830 ;
        RECT 1433.630 3194.140 1434.010 3194.460 ;
        RECT 1681.150 3194.450 1681.450 3194.830 ;
        RECT 2042.670 3194.820 2043.050 3194.830 ;
        RECT 1712.390 3194.450 1712.770 3194.460 ;
        RECT 1681.150 3194.150 1712.770 3194.450 ;
        RECT 2045.470 3194.450 2045.770 3194.830 ;
        RECT 2089.590 3194.450 2089.970 3194.460 ;
        RECT 2045.470 3194.150 2089.970 3194.450 ;
        RECT 1712.390 3194.140 1712.770 3194.150 ;
        RECT 2089.590 3194.140 2089.970 3194.150 ;
        RECT 24.445 3192.410 24.775 3192.425 ;
        RECT 34.565 3192.410 34.895 3192.425 ;
        RECT 24.445 3192.110 34.895 3192.410 ;
        RECT 24.445 3192.095 24.775 3192.110 ;
        RECT 34.565 3192.095 34.895 3192.110 ;
        RECT 86.085 3192.410 86.415 3192.425 ;
        RECT 131.165 3192.410 131.495 3192.425 ;
        RECT 86.085 3192.110 131.495 3192.410 ;
        RECT 86.085 3192.095 86.415 3192.110 ;
        RECT 131.165 3192.095 131.495 3192.110 ;
        RECT 182.685 3192.410 183.015 3192.425 ;
        RECT 227.765 3192.410 228.095 3192.425 ;
        RECT 182.685 3192.110 228.095 3192.410 ;
        RECT 182.685 3192.095 183.015 3192.110 ;
        RECT 227.765 3192.095 228.095 3192.110 ;
        RECT 279.285 3192.410 279.615 3192.425 ;
        RECT 324.365 3192.410 324.695 3192.425 ;
        RECT 279.285 3192.110 324.695 3192.410 ;
        RECT 279.285 3192.095 279.615 3192.110 ;
        RECT 324.365 3192.095 324.695 3192.110 ;
        RECT 375.885 3192.410 376.215 3192.425 ;
        RECT 420.965 3192.410 421.295 3192.425 ;
        RECT 375.885 3192.110 421.295 3192.410 ;
        RECT 375.885 3192.095 376.215 3192.110 ;
        RECT 420.965 3192.095 421.295 3192.110 ;
        RECT 472.485 3192.410 472.815 3192.425 ;
        RECT 517.565 3192.410 517.895 3192.425 ;
        RECT 472.485 3192.110 517.895 3192.410 ;
        RECT 472.485 3192.095 472.815 3192.110 ;
        RECT 517.565 3192.095 517.895 3192.110 ;
        RECT 569.085 3192.410 569.415 3192.425 ;
        RECT 614.165 3192.410 614.495 3192.425 ;
        RECT 569.085 3192.110 614.495 3192.410 ;
        RECT 569.085 3192.095 569.415 3192.110 ;
        RECT 614.165 3192.095 614.495 3192.110 ;
        RECT 665.685 3192.410 666.015 3192.425 ;
        RECT 710.765 3192.410 711.095 3192.425 ;
        RECT 665.685 3192.110 711.095 3192.410 ;
        RECT 665.685 3192.095 666.015 3192.110 ;
        RECT 710.765 3192.095 711.095 3192.110 ;
        RECT 762.285 3192.410 762.615 3192.425 ;
        RECT 807.365 3192.410 807.695 3192.425 ;
        RECT 762.285 3192.110 807.695 3192.410 ;
        RECT 762.285 3192.095 762.615 3192.110 ;
        RECT 807.365 3192.095 807.695 3192.110 ;
        RECT 858.885 3192.410 859.215 3192.425 ;
        RECT 903.965 3192.410 904.295 3192.425 ;
        RECT 858.885 3192.110 904.295 3192.410 ;
        RECT 858.885 3192.095 859.215 3192.110 ;
        RECT 903.965 3192.095 904.295 3192.110 ;
        RECT 955.485 3192.410 955.815 3192.425 ;
        RECT 1000.565 3192.410 1000.895 3192.425 ;
        RECT 955.485 3192.110 1000.895 3192.410 ;
        RECT 955.485 3192.095 955.815 3192.110 ;
        RECT 1000.565 3192.095 1000.895 3192.110 ;
        RECT 1052.085 3192.410 1052.415 3192.425 ;
        RECT 1100.385 3192.410 1100.715 3192.425 ;
        RECT 1052.085 3192.110 1100.715 3192.410 ;
        RECT 1052.085 3192.095 1052.415 3192.110 ;
        RECT 1100.385 3192.095 1100.715 3192.110 ;
        RECT 1171.430 3192.410 1171.810 3192.420 ;
        RECT 1197.190 3192.410 1197.570 3192.420 ;
        RECT 1171.430 3192.110 1197.570 3192.410 ;
        RECT 1171.430 3192.100 1171.810 3192.110 ;
        RECT 1197.190 3192.100 1197.570 3192.110 ;
        RECT 1221.110 3192.410 1221.490 3192.420 ;
        RECT 1290.110 3192.410 1290.490 3192.420 ;
        RECT 1221.110 3192.110 1290.490 3192.410 ;
        RECT 1221.110 3192.100 1221.490 3192.110 ;
        RECT 1290.110 3192.100 1290.490 3192.110 ;
        RECT 1337.950 3192.410 1338.330 3192.420 ;
        RECT 1387.630 3192.410 1388.010 3192.420 ;
        RECT 1337.950 3192.110 1388.010 3192.410 ;
        RECT 1337.950 3192.100 1338.330 3192.110 ;
        RECT 1387.630 3192.100 1388.010 3192.110 ;
        RECT 1433.630 3192.410 1434.010 3192.420 ;
        RECT 1483.310 3192.410 1483.690 3192.420 ;
        RECT 1433.630 3192.110 1483.690 3192.410 ;
        RECT 1433.630 3192.100 1434.010 3192.110 ;
        RECT 1483.310 3192.100 1483.690 3192.110 ;
        RECT 1532.990 3192.410 1533.370 3192.420 ;
        RECT 1579.910 3192.410 1580.290 3192.420 ;
        RECT 1532.990 3192.110 1580.290 3192.410 ;
        RECT 1532.990 3192.100 1533.370 3192.110 ;
        RECT 1579.910 3192.100 1580.290 3192.110 ;
        RECT 1627.750 3192.410 1628.130 3192.420 ;
        RECT 1676.510 3192.410 1676.890 3192.420 ;
        RECT 1627.750 3192.110 1676.890 3192.410 ;
        RECT 1627.750 3192.100 1628.130 3192.110 ;
        RECT 1676.510 3192.100 1676.890 3192.110 ;
        RECT 1777.710 3192.410 1778.090 3192.420 ;
        RECT 1820.950 3192.410 1821.330 3192.420 ;
        RECT 1777.710 3192.110 1821.330 3192.410 ;
        RECT 1777.710 3192.100 1778.090 3192.110 ;
        RECT 1820.950 3192.100 1821.330 3192.110 ;
        RECT 1874.310 3192.410 1874.690 3192.420 ;
        RECT 1920.310 3192.410 1920.690 3192.420 ;
        RECT 1874.310 3192.110 1920.690 3192.410 ;
        RECT 1874.310 3192.100 1874.690 3192.110 ;
        RECT 1920.310 3192.100 1920.690 3192.110 ;
        RECT 2089.590 3192.410 2089.970 3192.420 ;
        RECT 2442.870 3192.410 2443.250 3192.420 ;
        RECT 2089.590 3192.110 2443.250 3192.410 ;
        RECT 2089.590 3192.100 2089.970 3192.110 ;
        RECT 2442.870 3192.100 2443.250 3192.110 ;
        RECT 34.565 3190.370 34.895 3190.385 ;
        RECT 86.085 3190.370 86.415 3190.385 ;
        RECT 34.565 3190.070 86.415 3190.370 ;
        RECT 34.565 3190.055 34.895 3190.070 ;
        RECT 86.085 3190.055 86.415 3190.070 ;
        RECT 131.625 3190.370 131.955 3190.385 ;
        RECT 182.685 3190.370 183.015 3190.385 ;
        RECT 131.625 3190.070 183.015 3190.370 ;
        RECT 131.625 3190.055 131.955 3190.070 ;
        RECT 182.685 3190.055 183.015 3190.070 ;
        RECT 228.225 3190.370 228.555 3190.385 ;
        RECT 279.285 3190.370 279.615 3190.385 ;
        RECT 228.225 3190.070 279.615 3190.370 ;
        RECT 228.225 3190.055 228.555 3190.070 ;
        RECT 279.285 3190.055 279.615 3190.070 ;
        RECT 324.825 3190.370 325.155 3190.385 ;
        RECT 375.885 3190.370 376.215 3190.385 ;
        RECT 324.825 3190.070 376.215 3190.370 ;
        RECT 324.825 3190.055 325.155 3190.070 ;
        RECT 375.885 3190.055 376.215 3190.070 ;
        RECT 421.425 3190.370 421.755 3190.385 ;
        RECT 472.485 3190.370 472.815 3190.385 ;
        RECT 421.425 3190.070 472.815 3190.370 ;
        RECT 421.425 3190.055 421.755 3190.070 ;
        RECT 472.485 3190.055 472.815 3190.070 ;
        RECT 518.025 3190.370 518.355 3190.385 ;
        RECT 569.085 3190.370 569.415 3190.385 ;
        RECT 518.025 3190.070 569.415 3190.370 ;
        RECT 518.025 3190.055 518.355 3190.070 ;
        RECT 569.085 3190.055 569.415 3190.070 ;
        RECT 614.625 3190.370 614.955 3190.385 ;
        RECT 665.685 3190.370 666.015 3190.385 ;
        RECT 614.625 3190.070 666.015 3190.370 ;
        RECT 614.625 3190.055 614.955 3190.070 ;
        RECT 665.685 3190.055 666.015 3190.070 ;
        RECT 711.225 3190.370 711.555 3190.385 ;
        RECT 762.285 3190.370 762.615 3190.385 ;
        RECT 711.225 3190.070 762.615 3190.370 ;
        RECT 711.225 3190.055 711.555 3190.070 ;
        RECT 762.285 3190.055 762.615 3190.070 ;
        RECT 807.825 3190.370 808.155 3190.385 ;
        RECT 858.885 3190.370 859.215 3190.385 ;
        RECT 807.825 3190.070 859.215 3190.370 ;
        RECT 807.825 3190.055 808.155 3190.070 ;
        RECT 858.885 3190.055 859.215 3190.070 ;
        RECT 904.425 3190.370 904.755 3190.385 ;
        RECT 955.485 3190.370 955.815 3190.385 ;
        RECT 904.425 3190.070 955.815 3190.370 ;
        RECT 904.425 3190.055 904.755 3190.070 ;
        RECT 955.485 3190.055 955.815 3190.070 ;
        RECT 1001.025 3190.370 1001.355 3190.385 ;
        RECT 1052.085 3190.370 1052.415 3190.385 ;
        RECT 1001.025 3190.070 1052.415 3190.370 ;
        RECT 1001.025 3190.055 1001.355 3190.070 ;
        RECT 1052.085 3190.055 1052.415 3190.070 ;
        RECT 1290.110 3190.370 1290.490 3190.380 ;
        RECT 1337.950 3190.370 1338.330 3190.380 ;
        RECT 1290.110 3190.070 1338.330 3190.370 ;
        RECT 1290.110 3190.060 1290.490 3190.070 ;
        RECT 1337.950 3190.060 1338.330 3190.070 ;
        RECT 1100.385 3189.690 1100.715 3189.705 ;
        RECT 1171.430 3189.690 1171.810 3189.700 ;
        RECT 1100.385 3189.390 1171.810 3189.690 ;
        RECT 1100.385 3189.375 1100.715 3189.390 ;
        RECT 1171.430 3189.380 1171.810 3189.390 ;
        RECT 1197.190 3189.690 1197.570 3189.700 ;
        RECT 1221.110 3189.690 1221.490 3189.700 ;
        RECT 1197.190 3189.390 1221.490 3189.690 ;
        RECT 1197.190 3189.380 1197.570 3189.390 ;
        RECT 1221.110 3189.380 1221.490 3189.390 ;
        RECT 1483.310 3189.010 1483.690 3189.020 ;
        RECT 1532.990 3189.010 1533.370 3189.020 ;
        RECT 1483.310 3188.710 1533.370 3189.010 ;
        RECT 1483.310 3188.700 1483.690 3188.710 ;
        RECT 1532.990 3188.700 1533.370 3188.710 ;
        RECT -4.800 1185.050 2.400 1185.500 ;
        RECT 13.865 1185.050 14.195 1185.065 ;
        RECT -4.800 1184.750 14.195 1185.050 ;
        RECT -4.800 1184.300 2.400 1184.750 ;
        RECT 13.865 1184.735 14.195 1184.750 ;
      LAYER via3 ;
        RECT 1579.940 3195.500 1580.260 3195.820 ;
        RECT 1627.780 3195.500 1628.100 3195.820 ;
        RECT 1712.420 3195.500 1712.740 3195.820 ;
        RECT 1777.740 3195.500 1778.060 3195.820 ;
        RECT 1820.980 3195.500 1821.300 3195.820 ;
        RECT 1387.660 3194.820 1387.980 3195.140 ;
        RECT 1676.540 3194.820 1676.860 3195.140 ;
        RECT 1874.340 3195.500 1874.660 3195.820 ;
        RECT 1920.340 3195.500 1920.660 3195.820 ;
        RECT 1993.020 3195.500 1993.340 3195.820 ;
        RECT 1994.860 3195.500 1995.180 3195.820 ;
        RECT 2042.700 3196.180 2043.020 3196.500 ;
        RECT 2442.900 3196.180 2443.220 3196.500 ;
        RECT 1433.660 3194.140 1433.980 3194.460 ;
        RECT 2042.700 3194.820 2043.020 3195.140 ;
        RECT 1712.420 3194.140 1712.740 3194.460 ;
        RECT 2089.620 3194.140 2089.940 3194.460 ;
        RECT 1171.460 3192.100 1171.780 3192.420 ;
        RECT 1197.220 3192.100 1197.540 3192.420 ;
        RECT 1221.140 3192.100 1221.460 3192.420 ;
        RECT 1290.140 3192.100 1290.460 3192.420 ;
        RECT 1337.980 3192.100 1338.300 3192.420 ;
        RECT 1387.660 3192.100 1387.980 3192.420 ;
        RECT 1433.660 3192.100 1433.980 3192.420 ;
        RECT 1483.340 3192.100 1483.660 3192.420 ;
        RECT 1533.020 3192.100 1533.340 3192.420 ;
        RECT 1579.940 3192.100 1580.260 3192.420 ;
        RECT 1627.780 3192.100 1628.100 3192.420 ;
        RECT 1676.540 3192.100 1676.860 3192.420 ;
        RECT 1777.740 3192.100 1778.060 3192.420 ;
        RECT 1820.980 3192.100 1821.300 3192.420 ;
        RECT 1874.340 3192.100 1874.660 3192.420 ;
        RECT 1920.340 3192.100 1920.660 3192.420 ;
        RECT 2089.620 3192.100 2089.940 3192.420 ;
        RECT 2442.900 3192.100 2443.220 3192.420 ;
        RECT 1290.140 3190.060 1290.460 3190.380 ;
        RECT 1337.980 3190.060 1338.300 3190.380 ;
        RECT 1171.460 3189.380 1171.780 3189.700 ;
        RECT 1197.220 3189.380 1197.540 3189.700 ;
        RECT 1221.140 3189.380 1221.460 3189.700 ;
        RECT 1483.340 3188.700 1483.660 3189.020 ;
        RECT 1533.020 3188.700 1533.340 3189.020 ;
      LAYER met4 ;
        RECT 2042.695 3196.175 2043.025 3196.505 ;
        RECT 2442.895 3196.175 2443.225 3196.505 ;
        RECT 1579.935 3195.495 1580.265 3195.825 ;
        RECT 1627.775 3195.495 1628.105 3195.825 ;
        RECT 1712.415 3195.495 1712.745 3195.825 ;
        RECT 1777.735 3195.495 1778.065 3195.825 ;
        RECT 1820.975 3195.495 1821.305 3195.825 ;
        RECT 1874.335 3195.495 1874.665 3195.825 ;
        RECT 1920.335 3195.495 1920.665 3195.825 ;
        RECT 1993.015 3195.495 1993.345 3195.825 ;
        RECT 1994.855 3195.495 1995.185 3195.825 ;
        RECT 1387.655 3194.815 1387.985 3195.145 ;
        RECT 1387.670 3192.425 1387.970 3194.815 ;
        RECT 1433.655 3194.135 1433.985 3194.465 ;
        RECT 1433.670 3192.425 1433.970 3194.135 ;
        RECT 1579.950 3192.425 1580.250 3195.495 ;
        RECT 1627.790 3192.425 1628.090 3195.495 ;
        RECT 1676.535 3194.815 1676.865 3195.145 ;
        RECT 1676.550 3192.425 1676.850 3194.815 ;
        RECT 1712.430 3194.465 1712.730 3195.495 ;
        RECT 1712.415 3194.135 1712.745 3194.465 ;
        RECT 1777.750 3192.425 1778.050 3195.495 ;
        RECT 1820.990 3192.425 1821.290 3195.495 ;
        RECT 1874.350 3192.425 1874.650 3195.495 ;
        RECT 1920.350 3192.425 1920.650 3195.495 ;
        RECT 1993.030 3194.450 1993.330 3195.495 ;
        RECT 1994.870 3194.450 1995.170 3195.495 ;
        RECT 2042.710 3195.145 2043.010 3196.175 ;
        RECT 2042.695 3194.815 2043.025 3195.145 ;
        RECT 1993.030 3194.150 1995.170 3194.450 ;
        RECT 2089.615 3194.135 2089.945 3194.465 ;
        RECT 2089.630 3192.425 2089.930 3194.135 ;
        RECT 2442.910 3192.425 2443.210 3196.175 ;
        RECT 1171.455 3192.095 1171.785 3192.425 ;
        RECT 1197.215 3192.095 1197.545 3192.425 ;
        RECT 1221.135 3192.095 1221.465 3192.425 ;
        RECT 1290.135 3192.095 1290.465 3192.425 ;
        RECT 1337.975 3192.095 1338.305 3192.425 ;
        RECT 1387.655 3192.095 1387.985 3192.425 ;
        RECT 1433.655 3192.095 1433.985 3192.425 ;
        RECT 1483.335 3192.095 1483.665 3192.425 ;
        RECT 1533.015 3192.095 1533.345 3192.425 ;
        RECT 1579.935 3192.095 1580.265 3192.425 ;
        RECT 1627.775 3192.095 1628.105 3192.425 ;
        RECT 1676.535 3192.095 1676.865 3192.425 ;
        RECT 1777.735 3192.095 1778.065 3192.425 ;
        RECT 1820.975 3192.095 1821.305 3192.425 ;
        RECT 1874.335 3192.095 1874.665 3192.425 ;
        RECT 1920.335 3192.095 1920.665 3192.425 ;
        RECT 2089.615 3192.095 2089.945 3192.425 ;
        RECT 2442.895 3192.095 2443.225 3192.425 ;
        RECT 1171.470 3189.705 1171.770 3192.095 ;
        RECT 1197.230 3189.705 1197.530 3192.095 ;
        RECT 1221.150 3189.705 1221.450 3192.095 ;
        RECT 1290.150 3190.385 1290.450 3192.095 ;
        RECT 1337.990 3190.385 1338.290 3192.095 ;
        RECT 1290.135 3190.055 1290.465 3190.385 ;
        RECT 1337.975 3190.055 1338.305 3190.385 ;
        RECT 1171.455 3189.375 1171.785 3189.705 ;
        RECT 1197.215 3189.375 1197.545 3189.705 ;
        RECT 1221.135 3189.375 1221.465 3189.705 ;
        RECT 1483.350 3189.025 1483.650 3192.095 ;
        RECT 1533.030 3189.025 1533.330 3192.095 ;
        RECT 1483.335 3188.695 1483.665 3189.025 ;
        RECT 1533.015 3188.695 1533.345 3189.025 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 19.850 3209.500 20.170 3209.560 ;
        RECT 2484.070 3209.500 2484.390 3209.560 ;
        RECT 19.850 3209.360 2484.390 3209.500 ;
        RECT 19.850 3209.300 20.170 3209.360 ;
        RECT 2484.070 3209.300 2484.390 3209.360 ;
      LAYER via ;
        RECT 19.880 3209.300 20.140 3209.560 ;
        RECT 2484.100 3209.300 2484.360 3209.560 ;
      LAYER met2 ;
        RECT 19.880 3209.270 20.140 3209.590 ;
        RECT 2484.100 3209.270 2484.360 3209.590 ;
        RECT 19.940 969.525 20.080 3209.270 ;
        RECT 2484.160 3200.000 2484.300 3209.270 ;
        RECT 2484.020 3196.000 2484.300 3200.000 ;
        RECT 19.870 969.155 20.150 969.525 ;
      LAYER via2 ;
        RECT 19.870 969.200 20.150 969.480 ;
      LAYER met3 ;
        RECT -4.800 969.490 2.400 969.940 ;
        RECT 19.845 969.490 20.175 969.505 ;
        RECT -4.800 969.190 20.175 969.490 ;
        RECT -4.800 968.740 2.400 969.190 ;
        RECT 19.845 969.175 20.175 969.190 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2523.190 3209.075 2523.470 3209.445 ;
        RECT 2523.260 3200.000 2523.400 3209.075 ;
        RECT 2523.120 3196.000 2523.400 3200.000 ;
        RECT 16.650 758.355 16.930 758.725 ;
        RECT 16.720 753.965 16.860 758.355 ;
        RECT 16.650 753.595 16.930 753.965 ;
      LAYER via2 ;
        RECT 2523.190 3209.120 2523.470 3209.400 ;
        RECT 16.650 758.400 16.930 758.680 ;
        RECT 16.650 753.640 16.930 753.920 ;
      LAYER met3 ;
        RECT 1292.870 3209.410 1293.250 3209.420 ;
        RECT 2523.165 3209.410 2523.495 3209.425 ;
        RECT 1292.870 3209.110 2523.495 3209.410 ;
        RECT 1292.870 3209.100 1293.250 3209.110 ;
        RECT 2523.165 3209.095 2523.495 3209.110 ;
        RECT 16.625 758.690 16.955 758.705 ;
        RECT 1292.870 758.690 1293.250 758.700 ;
        RECT 16.625 758.390 1293.250 758.690 ;
        RECT 16.625 758.375 16.955 758.390 ;
        RECT 1292.870 758.380 1293.250 758.390 ;
        RECT -4.800 753.930 2.400 754.380 ;
        RECT 16.625 753.930 16.955 753.945 ;
        RECT -4.800 753.630 16.955 753.930 ;
        RECT -4.800 753.180 2.400 753.630 ;
        RECT 16.625 753.615 16.955 753.630 ;
      LAYER via3 ;
        RECT 1292.900 3209.100 1293.220 3209.420 ;
        RECT 1292.900 758.380 1293.220 758.700 ;
      LAYER met4 ;
        RECT 1292.895 3209.095 1293.225 3209.425 ;
        RECT 1292.910 758.705 1293.210 3209.095 ;
        RECT 1292.895 758.375 1293.225 758.705 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.930 3208.820 19.250 3208.880 ;
        RECT 2562.730 3208.820 2563.050 3208.880 ;
        RECT 18.930 3208.680 2563.050 3208.820 ;
        RECT 18.930 3208.620 19.250 3208.680 ;
        RECT 2562.730 3208.620 2563.050 3208.680 ;
      LAYER via ;
        RECT 18.960 3208.620 19.220 3208.880 ;
        RECT 2562.760 3208.620 2563.020 3208.880 ;
      LAYER met2 ;
        RECT 18.960 3208.590 19.220 3208.910 ;
        RECT 2562.760 3208.590 2563.020 3208.910 ;
        RECT 19.020 538.405 19.160 3208.590 ;
        RECT 2562.820 3200.000 2562.960 3208.590 ;
        RECT 2562.680 3196.000 2562.960 3200.000 ;
        RECT 18.950 538.035 19.230 538.405 ;
      LAYER via2 ;
        RECT 18.950 538.080 19.230 538.360 ;
      LAYER met3 ;
        RECT -4.800 538.370 2.400 538.820 ;
        RECT 18.925 538.370 19.255 538.385 ;
        RECT -4.800 538.070 19.255 538.370 ;
        RECT -4.800 537.620 2.400 538.070 ;
        RECT 18.925 538.055 19.255 538.070 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2601.445 3194.725 2601.615 3199.655 ;
      LAYER mcon ;
        RECT 2601.445 3199.485 2601.615 3199.655 ;
      LAYER met1 ;
        RECT 2601.370 3199.640 2601.690 3199.700 ;
        RECT 2601.175 3199.500 2601.690 3199.640 ;
        RECT 2601.370 3199.440 2601.690 3199.500 ;
        RECT 18.010 3194.880 18.330 3194.940 ;
        RECT 2601.385 3194.880 2601.675 3194.925 ;
        RECT 18.010 3194.740 2601.675 3194.880 ;
        RECT 18.010 3194.680 18.330 3194.740 ;
        RECT 2601.385 3194.695 2601.675 3194.740 ;
      LAYER via ;
        RECT 2601.400 3199.440 2601.660 3199.700 ;
        RECT 18.040 3194.680 18.300 3194.940 ;
      LAYER met2 ;
        RECT 2602.240 3199.810 2602.520 3200.000 ;
        RECT 2601.460 3199.730 2602.520 3199.810 ;
        RECT 2601.400 3199.670 2602.520 3199.730 ;
        RECT 2601.400 3199.410 2601.660 3199.670 ;
        RECT 2602.240 3196.000 2602.520 3199.670 ;
        RECT 18.040 3194.650 18.300 3194.970 ;
        RECT 18.100 322.845 18.240 3194.650 ;
        RECT 18.030 322.475 18.310 322.845 ;
      LAYER via2 ;
        RECT 18.030 322.520 18.310 322.800 ;
      LAYER met3 ;
        RECT -4.800 322.810 2.400 323.260 ;
        RECT 18.005 322.810 18.335 322.825 ;
        RECT -4.800 322.510 18.335 322.810 ;
        RECT -4.800 322.060 2.400 322.510 ;
        RECT 18.005 322.495 18.335 322.510 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2640.490 3196.410 2640.770 3196.525 ;
        RECT 2641.800 3196.410 2642.080 3200.000 ;
        RECT 2640.490 3196.270 2642.080 3196.410 ;
        RECT 2640.490 3196.155 2640.770 3196.270 ;
        RECT 2641.800 3196.000 2642.080 3196.270 ;
      LAYER via2 ;
        RECT 2640.490 3196.200 2640.770 3196.480 ;
      LAYER met3 ;
        RECT 2636.070 3196.490 2636.450 3196.500 ;
        RECT 2640.465 3196.490 2640.795 3196.505 ;
        RECT 2636.070 3196.190 2640.795 3196.490 ;
        RECT 2636.070 3196.180 2636.450 3196.190 ;
        RECT 2640.465 3196.175 2640.795 3196.190 ;
        RECT 2636.070 2852.410 2636.450 2852.420 ;
        RECT 2635.190 2852.110 2636.450 2852.410 ;
        RECT 2635.190 2850.370 2635.490 2852.110 ;
        RECT 2636.070 2852.100 2636.450 2852.110 ;
        RECT 2636.070 2850.370 2636.450 2850.380 ;
        RECT 2635.190 2850.070 2636.450 2850.370 ;
        RECT 2636.070 2850.060 2636.450 2850.070 ;
        RECT 2636.070 2141.810 2636.450 2141.820 ;
        RECT 2638.830 2141.810 2639.210 2141.820 ;
        RECT 2636.070 2141.510 2639.210 2141.810 ;
        RECT 2636.070 2141.500 2636.450 2141.510 ;
        RECT 2638.830 2141.500 2639.210 2141.510 ;
        RECT 2636.070 2108.490 2636.450 2108.500 ;
        RECT 2638.830 2108.490 2639.210 2108.500 ;
        RECT 2636.070 2108.190 2639.210 2108.490 ;
        RECT 2636.070 2108.180 2636.450 2108.190 ;
        RECT 2638.830 2108.180 2639.210 2108.190 ;
        RECT 2636.070 109.970 2636.450 109.980 ;
        RECT 3.070 109.670 2636.450 109.970 ;
        RECT -4.800 107.250 2.400 107.700 ;
        RECT 3.070 107.250 3.370 109.670 ;
        RECT 2636.070 109.660 2636.450 109.670 ;
        RECT -4.800 106.950 3.370 107.250 ;
        RECT -4.800 106.500 2.400 106.950 ;
      LAYER via3 ;
        RECT 2636.100 3196.180 2636.420 3196.500 ;
        RECT 2636.100 2852.100 2636.420 2852.420 ;
        RECT 2636.100 2850.060 2636.420 2850.380 ;
        RECT 2636.100 2141.500 2636.420 2141.820 ;
        RECT 2638.860 2141.500 2639.180 2141.820 ;
        RECT 2636.100 2108.180 2636.420 2108.500 ;
        RECT 2638.860 2108.180 2639.180 2108.500 ;
        RECT 2636.100 109.660 2636.420 109.980 ;
      LAYER met4 ;
        RECT 2636.095 3196.175 2636.425 3196.505 ;
        RECT 2636.110 2852.425 2636.410 3196.175 ;
        RECT 2636.095 2852.095 2636.425 2852.425 ;
        RECT 2636.095 2850.055 2636.425 2850.385 ;
        RECT 2636.110 2141.825 2636.410 2850.055 ;
        RECT 2636.095 2141.495 2636.425 2141.825 ;
        RECT 2638.855 2141.495 2639.185 2141.825 ;
        RECT 2638.870 2108.505 2639.170 2141.495 ;
        RECT 2636.095 2108.175 2636.425 2108.505 ;
        RECT 2638.855 2108.175 2639.185 2108.505 ;
        RECT 2636.110 109.985 2636.410 2108.175 ;
        RECT 2636.095 109.655 2636.425 109.985 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1441.710 850.580 1442.030 850.640 ;
        RECT 1483.110 850.580 1483.430 850.640 ;
        RECT 1441.710 850.440 1483.430 850.580 ;
        RECT 1441.710 850.380 1442.030 850.440 ;
        RECT 1483.110 850.380 1483.430 850.440 ;
        RECT 1641.810 850.240 1642.130 850.300 ;
        RECT 1683.210 850.240 1683.530 850.300 ;
        RECT 1641.810 850.100 1683.530 850.240 ;
        RECT 1641.810 850.040 1642.130 850.100 ;
        RECT 1683.210 850.040 1683.530 850.100 ;
        RECT 1828.570 849.900 1828.890 849.960 ;
        RECT 1841.450 849.900 1841.770 849.960 ;
        RECT 1828.570 849.760 1841.770 849.900 ;
        RECT 1828.570 849.700 1828.890 849.760 ;
        RECT 1841.450 849.700 1841.770 849.760 ;
        RECT 2270.170 849.900 2270.490 849.960 ;
        RECT 2290.870 849.900 2291.190 849.960 ;
        RECT 2270.170 849.760 2291.190 849.900 ;
        RECT 2270.170 849.700 2270.490 849.760 ;
        RECT 2290.870 849.700 2291.190 849.760 ;
        RECT 2572.850 849.900 2573.170 849.960 ;
        RECT 2584.350 849.900 2584.670 849.960 ;
        RECT 2572.850 849.760 2584.670 849.900 ;
        RECT 2572.850 849.700 2573.170 849.760 ;
        RECT 2584.350 849.700 2584.670 849.760 ;
        RECT 2379.650 849.560 2379.970 849.620 ;
        RECT 2380.570 849.560 2380.890 849.620 ;
        RECT 2379.650 849.420 2380.890 849.560 ;
        RECT 2379.650 849.360 2379.970 849.420 ;
        RECT 2380.570 849.360 2380.890 849.420 ;
        RECT 1545.210 849.220 1545.530 849.280 ;
        RECT 1586.610 849.220 1586.930 849.280 ;
        RECT 1545.210 849.080 1586.930 849.220 ;
        RECT 1545.210 849.020 1545.530 849.080 ;
        RECT 1586.610 849.020 1586.930 849.080 ;
        RECT 2125.270 849.220 2125.590 849.280 ;
        RECT 2172.650 849.220 2172.970 849.280 ;
        RECT 2125.270 849.080 2172.970 849.220 ;
        RECT 2125.270 849.020 2125.590 849.080 ;
        RECT 2172.650 849.020 2172.970 849.080 ;
        RECT 2621.150 849.220 2621.470 849.280 ;
        RECT 2632.190 849.220 2632.510 849.280 ;
        RECT 2621.150 849.080 2632.510 849.220 ;
        RECT 2621.150 849.020 2621.470 849.080 ;
        RECT 2632.190 849.020 2632.510 849.080 ;
        RECT 1496.910 848.540 1497.230 848.600 ;
        RECT 1514.850 848.540 1515.170 848.600 ;
        RECT 1496.910 848.400 1515.170 848.540 ;
        RECT 1496.910 848.340 1497.230 848.400 ;
        RECT 1514.850 848.340 1515.170 848.400 ;
      LAYER via ;
        RECT 1441.740 850.380 1442.000 850.640 ;
        RECT 1483.140 850.380 1483.400 850.640 ;
        RECT 1641.840 850.040 1642.100 850.300 ;
        RECT 1683.240 850.040 1683.500 850.300 ;
        RECT 1828.600 849.700 1828.860 849.960 ;
        RECT 1841.480 849.700 1841.740 849.960 ;
        RECT 2270.200 849.700 2270.460 849.960 ;
        RECT 2290.900 849.700 2291.160 849.960 ;
        RECT 2572.880 849.700 2573.140 849.960 ;
        RECT 2584.380 849.700 2584.640 849.960 ;
        RECT 2379.680 849.360 2379.940 849.620 ;
        RECT 2380.600 849.360 2380.860 849.620 ;
        RECT 1545.240 849.020 1545.500 849.280 ;
        RECT 1586.640 849.020 1586.900 849.280 ;
        RECT 2125.300 849.020 2125.560 849.280 ;
        RECT 2172.680 849.020 2172.940 849.280 ;
        RECT 2621.180 849.020 2621.440 849.280 ;
        RECT 2632.220 849.020 2632.480 849.280 ;
        RECT 1496.940 848.340 1497.200 848.600 ;
        RECT 1514.880 848.340 1515.140 848.600 ;
      LAYER met2 ;
        RECT 1299.520 3196.410 1299.800 3200.000 ;
        RECT 1301.430 3196.410 1301.710 3196.525 ;
        RECT 1299.520 3196.270 1301.710 3196.410 ;
        RECT 1299.520 3196.000 1299.800 3196.270 ;
        RECT 1301.430 3196.155 1301.710 3196.270 ;
        RECT 1344.670 856.275 1344.950 856.645 ;
        RECT 1344.740 850.525 1344.880 856.275 ;
        RECT 2704.430 850.835 2704.710 851.205 ;
        RECT 1441.740 850.525 1442.000 850.670 ;
        RECT 1483.140 850.525 1483.400 850.670 ;
        RECT 1344.670 850.155 1344.950 850.525 ;
        RECT 1441.730 850.155 1442.010 850.525 ;
        RECT 1483.130 850.155 1483.410 850.525 ;
        RECT 1490.030 850.155 1490.310 850.525 ;
        RECT 1586.630 850.155 1586.910 850.525 ;
        RECT 1641.830 850.155 1642.110 850.525 ;
        RECT 1683.230 850.155 1683.510 850.525 ;
        RECT 1896.670 850.410 1896.950 850.525 ;
        RECT 1897.590 850.410 1897.870 850.525 ;
        RECT 1896.670 850.270 1897.870 850.410 ;
        RECT 1896.670 850.155 1896.950 850.270 ;
        RECT 1897.590 850.155 1897.870 850.270 ;
        RECT 2172.670 850.155 2172.950 850.525 ;
        RECT 1490.100 849.165 1490.240 850.155 ;
        RECT 1586.700 849.310 1586.840 850.155 ;
        RECT 1641.840 850.010 1642.100 850.155 ;
        RECT 1683.240 850.010 1683.500 850.155 ;
        RECT 1828.600 849.845 1828.860 849.990 ;
        RECT 1841.480 849.845 1841.740 849.990 ;
        RECT 1828.590 849.475 1828.870 849.845 ;
        RECT 1841.470 849.475 1841.750 849.845 ;
        RECT 2090.330 849.475 2090.610 849.845 ;
        RECT 1545.240 849.165 1545.500 849.310 ;
        RECT 1490.030 848.795 1490.310 849.165 ;
        RECT 1545.230 848.795 1545.510 849.165 ;
        RECT 1586.640 848.990 1586.900 849.310 ;
        RECT 1496.940 848.485 1497.200 848.630 ;
        RECT 1514.880 848.485 1515.140 848.630 ;
        RECT 1496.930 848.115 1497.210 848.485 ;
        RECT 1514.870 848.115 1515.150 848.485 ;
        RECT 2090.400 847.805 2090.540 849.475 ;
        RECT 2172.740 849.310 2172.880 850.155 ;
        RECT 2270.200 849.845 2270.460 849.990 ;
        RECT 2290.900 849.845 2291.160 849.990 ;
        RECT 2572.880 849.845 2573.140 849.990 ;
        RECT 2584.380 849.845 2584.640 849.990 ;
        RECT 2270.190 849.475 2270.470 849.845 ;
        RECT 2290.890 849.475 2291.170 849.845 ;
        RECT 2379.670 849.475 2379.950 849.845 ;
        RECT 2380.590 849.475 2380.870 849.845 ;
        RECT 2572.870 849.475 2573.150 849.845 ;
        RECT 2584.370 849.475 2584.650 849.845 ;
        RECT 2632.210 849.475 2632.490 849.845 ;
        RECT 2379.680 849.330 2379.940 849.475 ;
        RECT 2380.600 849.330 2380.860 849.475 ;
        RECT 2632.280 849.310 2632.420 849.475 ;
        RECT 2125.300 849.165 2125.560 849.310 ;
        RECT 2125.290 848.795 2125.570 849.165 ;
        RECT 2172.680 848.990 2172.940 849.310 ;
        RECT 2621.180 849.165 2621.440 849.310 ;
        RECT 2621.170 848.795 2621.450 849.165 ;
        RECT 2632.220 848.990 2632.480 849.310 ;
        RECT 2704.500 849.165 2704.640 850.835 ;
        RECT 2801.030 850.155 2801.310 850.525 ;
        RECT 2704.430 848.795 2704.710 849.165 ;
        RECT 2801.100 848.485 2801.240 850.155 ;
        RECT 2863.130 849.475 2863.410 849.845 ;
        RECT 2863.200 849.050 2863.340 849.475 ;
        RECT 2863.590 849.050 2863.870 849.165 ;
        RECT 2863.200 848.910 2863.870 849.050 ;
        RECT 2863.590 848.795 2863.870 848.910 ;
        RECT 2801.030 848.115 2801.310 848.485 ;
        RECT 2090.330 847.435 2090.610 847.805 ;
      LAYER via2 ;
        RECT 1301.430 3196.200 1301.710 3196.480 ;
        RECT 1344.670 856.320 1344.950 856.600 ;
        RECT 2704.430 850.880 2704.710 851.160 ;
        RECT 1344.670 850.200 1344.950 850.480 ;
        RECT 1441.730 850.200 1442.010 850.480 ;
        RECT 1483.130 850.200 1483.410 850.480 ;
        RECT 1490.030 850.200 1490.310 850.480 ;
        RECT 1586.630 850.200 1586.910 850.480 ;
        RECT 1641.830 850.200 1642.110 850.480 ;
        RECT 1683.230 850.200 1683.510 850.480 ;
        RECT 1896.670 850.200 1896.950 850.480 ;
        RECT 1897.590 850.200 1897.870 850.480 ;
        RECT 2172.670 850.200 2172.950 850.480 ;
        RECT 1828.590 849.520 1828.870 849.800 ;
        RECT 1841.470 849.520 1841.750 849.800 ;
        RECT 2090.330 849.520 2090.610 849.800 ;
        RECT 1490.030 848.840 1490.310 849.120 ;
        RECT 1545.230 848.840 1545.510 849.120 ;
        RECT 1496.930 848.160 1497.210 848.440 ;
        RECT 1514.870 848.160 1515.150 848.440 ;
        RECT 2270.190 849.520 2270.470 849.800 ;
        RECT 2290.890 849.520 2291.170 849.800 ;
        RECT 2379.670 849.520 2379.950 849.800 ;
        RECT 2380.590 849.520 2380.870 849.800 ;
        RECT 2572.870 849.520 2573.150 849.800 ;
        RECT 2584.370 849.520 2584.650 849.800 ;
        RECT 2632.210 849.520 2632.490 849.800 ;
        RECT 2125.290 848.840 2125.570 849.120 ;
        RECT 2621.170 848.840 2621.450 849.120 ;
        RECT 2801.030 850.200 2801.310 850.480 ;
        RECT 2704.430 848.840 2704.710 849.120 ;
        RECT 2863.130 849.520 2863.410 849.800 ;
        RECT 2863.590 848.840 2863.870 849.120 ;
        RECT 2801.030 848.160 2801.310 848.440 ;
        RECT 2090.330 847.480 2090.610 847.760 ;
      LAYER met3 ;
        RECT 1301.405 3196.490 1301.735 3196.505 ;
        RECT 1306.670 3196.490 1307.050 3196.500 ;
        RECT 1301.405 3196.190 1307.050 3196.490 ;
        RECT 1301.405 3196.175 1301.735 3196.190 ;
        RECT 1306.670 3196.180 1307.050 3196.190 ;
        RECT 1306.670 856.610 1307.050 856.620 ;
        RECT 1344.645 856.610 1344.975 856.625 ;
        RECT 1306.670 856.310 1344.975 856.610 ;
        RECT 1306.670 856.300 1307.050 856.310 ;
        RECT 1344.645 856.295 1344.975 856.310 ;
        RECT 2656.310 851.170 2656.690 851.180 ;
        RECT 2704.405 851.170 2704.735 851.185 ;
        RECT 1751.990 850.870 1753.210 851.170 ;
        RECT 1344.645 850.490 1344.975 850.505 ;
        RECT 1441.705 850.490 1442.035 850.505 ;
        RECT 1344.645 850.190 1442.035 850.490 ;
        RECT 1344.645 850.175 1344.975 850.190 ;
        RECT 1441.705 850.175 1442.035 850.190 ;
        RECT 1483.105 850.490 1483.435 850.505 ;
        RECT 1490.005 850.490 1490.335 850.505 ;
        RECT 1483.105 850.190 1490.335 850.490 ;
        RECT 1483.105 850.175 1483.435 850.190 ;
        RECT 1490.005 850.175 1490.335 850.190 ;
        RECT 1586.605 850.490 1586.935 850.505 ;
        RECT 1641.805 850.490 1642.135 850.505 ;
        RECT 1586.605 850.190 1642.135 850.490 ;
        RECT 1586.605 850.175 1586.935 850.190 ;
        RECT 1641.805 850.175 1642.135 850.190 ;
        RECT 1683.205 850.490 1683.535 850.505 ;
        RECT 1683.205 850.190 1714.570 850.490 ;
        RECT 1683.205 850.175 1683.535 850.190 ;
        RECT 1714.270 849.810 1714.570 850.190 ;
        RECT 1751.990 849.810 1752.290 850.870 ;
        RECT 1752.910 850.490 1753.210 850.870 ;
        RECT 2476.030 850.870 2511.290 851.170 ;
        RECT 1896.645 850.490 1896.975 850.505 ;
        RECT 1752.910 850.190 1787.250 850.490 ;
        RECT 1714.270 849.510 1752.290 849.810 ;
        RECT 1786.950 849.810 1787.250 850.190 ;
        RECT 1876.190 850.190 1896.975 850.490 ;
        RECT 1828.565 849.810 1828.895 849.825 ;
        RECT 1786.950 849.510 1828.895 849.810 ;
        RECT 1828.565 849.495 1828.895 849.510 ;
        RECT 1841.445 849.810 1841.775 849.825 ;
        RECT 1876.190 849.810 1876.490 850.190 ;
        RECT 1896.645 850.175 1896.975 850.190 ;
        RECT 1897.565 850.490 1897.895 850.505 ;
        RECT 2172.645 850.490 2172.975 850.505 ;
        RECT 1897.565 850.190 1907.770 850.490 ;
        RECT 1897.565 850.175 1897.895 850.190 ;
        RECT 1841.445 849.510 1876.490 849.810 ;
        RECT 1907.470 849.810 1907.770 850.190 ;
        RECT 1932.310 850.190 1994.250 850.490 ;
        RECT 1932.310 849.810 1932.610 850.190 ;
        RECT 1907.470 849.510 1932.610 849.810 ;
        RECT 1841.445 849.495 1841.775 849.510 ;
        RECT 1490.005 849.130 1490.335 849.145 ;
        RECT 1545.205 849.130 1545.535 849.145 ;
        RECT 1490.005 848.830 1491.010 849.130 ;
        RECT 1490.005 848.815 1490.335 848.830 ;
        RECT 1490.710 848.450 1491.010 848.830 ;
        RECT 1538.550 848.830 1545.535 849.130 ;
        RECT 1993.950 849.130 1994.250 850.190 ;
        RECT 2172.645 850.190 2187.450 850.490 ;
        RECT 2172.645 850.175 2172.975 850.190 ;
        RECT 2090.305 849.810 2090.635 849.825 ;
        RECT 2042.710 849.510 2090.635 849.810 ;
        RECT 2042.710 849.130 2043.010 849.510 ;
        RECT 2090.305 849.495 2090.635 849.510 ;
        RECT 2125.265 849.130 2125.595 849.145 ;
        RECT 1993.950 848.830 2043.010 849.130 ;
        RECT 2124.590 848.830 2125.595 849.130 ;
        RECT 2187.150 849.130 2187.450 850.190 ;
        RECT 2270.165 849.810 2270.495 849.825 ;
        RECT 2235.910 849.510 2270.495 849.810 ;
        RECT 2235.910 849.130 2236.210 849.510 ;
        RECT 2270.165 849.495 2270.495 849.510 ;
        RECT 2290.865 849.810 2291.195 849.825 ;
        RECT 2379.645 849.810 2379.975 849.825 ;
        RECT 2290.865 849.510 2318.090 849.810 ;
        RECT 2290.865 849.495 2291.195 849.510 ;
        RECT 2187.150 848.830 2236.210 849.130 ;
        RECT 2317.790 849.130 2318.090 849.510 ;
        RECT 2332.510 849.510 2379.975 849.810 ;
        RECT 2332.510 849.130 2332.810 849.510 ;
        RECT 2379.645 849.495 2379.975 849.510 ;
        RECT 2380.565 849.810 2380.895 849.825 ;
        RECT 2476.030 849.810 2476.330 850.870 ;
        RECT 2380.565 849.510 2414.690 849.810 ;
        RECT 2380.565 849.495 2380.895 849.510 ;
        RECT 2317.790 848.830 2332.810 849.130 ;
        RECT 2414.390 849.130 2414.690 849.510 ;
        RECT 2429.110 849.510 2476.330 849.810 ;
        RECT 2429.110 849.130 2429.410 849.510 ;
        RECT 2414.390 848.830 2429.410 849.130 ;
        RECT 2510.990 849.130 2511.290 850.870 ;
        RECT 2656.310 850.870 2704.735 851.170 ;
        RECT 2656.310 850.860 2656.690 850.870 ;
        RECT 2704.405 850.855 2704.735 850.870 ;
        RECT 2801.005 850.490 2801.335 850.505 ;
        RECT 2917.600 850.490 2924.800 850.940 ;
        RECT 2801.005 850.190 2815.810 850.490 ;
        RECT 2801.005 850.175 2801.335 850.190 ;
        RECT 2572.845 849.810 2573.175 849.825 ;
        RECT 2525.710 849.510 2573.175 849.810 ;
        RECT 2525.710 849.130 2526.010 849.510 ;
        RECT 2572.845 849.495 2573.175 849.510 ;
        RECT 2584.345 849.810 2584.675 849.825 ;
        RECT 2632.185 849.810 2632.515 849.825 ;
        RECT 2656.310 849.810 2656.690 849.820 ;
        RECT 2752.910 849.810 2753.290 849.820 ;
        RECT 2584.345 849.510 2607.890 849.810 ;
        RECT 2584.345 849.495 2584.675 849.510 ;
        RECT 2510.990 848.830 2526.010 849.130 ;
        RECT 2607.590 849.130 2607.890 849.510 ;
        RECT 2632.185 849.510 2656.690 849.810 ;
        RECT 2632.185 849.495 2632.515 849.510 ;
        RECT 2656.310 849.500 2656.690 849.510 ;
        RECT 2718.910 849.510 2753.290 849.810 ;
        RECT 2621.145 849.130 2621.475 849.145 ;
        RECT 2607.590 848.830 2621.475 849.130 ;
        RECT 1496.905 848.450 1497.235 848.465 ;
        RECT 1490.710 848.150 1497.235 848.450 ;
        RECT 1496.905 848.135 1497.235 848.150 ;
        RECT 1514.845 848.450 1515.175 848.465 ;
        RECT 1538.550 848.450 1538.850 848.830 ;
        RECT 1545.205 848.815 1545.535 848.830 ;
        RECT 1514.845 848.150 1538.850 848.450 ;
        RECT 1514.845 848.135 1515.175 848.150 ;
        RECT 2090.305 847.770 2090.635 847.785 ;
        RECT 2124.590 847.770 2124.890 848.830 ;
        RECT 2125.265 848.815 2125.595 848.830 ;
        RECT 2621.145 848.815 2621.475 848.830 ;
        RECT 2704.405 849.130 2704.735 849.145 ;
        RECT 2718.910 849.130 2719.210 849.510 ;
        RECT 2752.910 849.500 2753.290 849.510 ;
        RECT 2704.405 848.830 2719.210 849.130 ;
        RECT 2815.510 849.130 2815.810 850.190 ;
        RECT 2916.710 850.190 2924.800 850.490 ;
        RECT 2863.105 849.810 2863.435 849.825 ;
        RECT 2916.710 849.810 2917.010 850.190 ;
        RECT 2849.550 849.510 2863.435 849.810 ;
        RECT 2849.550 849.130 2849.850 849.510 ;
        RECT 2863.105 849.495 2863.435 849.510 ;
        RECT 2884.510 849.510 2917.010 849.810 ;
        RECT 2917.600 849.740 2924.800 850.190 ;
        RECT 2815.510 848.830 2849.850 849.130 ;
        RECT 2863.565 849.130 2863.895 849.145 ;
        RECT 2884.510 849.130 2884.810 849.510 ;
        RECT 2863.565 848.830 2884.810 849.130 ;
        RECT 2704.405 848.815 2704.735 848.830 ;
        RECT 2863.565 848.815 2863.895 848.830 ;
        RECT 2752.910 848.450 2753.290 848.460 ;
        RECT 2801.005 848.450 2801.335 848.465 ;
        RECT 2752.910 848.150 2801.335 848.450 ;
        RECT 2752.910 848.140 2753.290 848.150 ;
        RECT 2801.005 848.135 2801.335 848.150 ;
        RECT 2090.305 847.470 2124.890 847.770 ;
        RECT 2090.305 847.455 2090.635 847.470 ;
      LAYER via3 ;
        RECT 1306.700 3196.180 1307.020 3196.500 ;
        RECT 1306.700 856.300 1307.020 856.620 ;
        RECT 2656.340 850.860 2656.660 851.180 ;
        RECT 2656.340 849.500 2656.660 849.820 ;
        RECT 2752.940 849.500 2753.260 849.820 ;
        RECT 2752.940 848.140 2753.260 848.460 ;
      LAYER met4 ;
        RECT 1306.695 3196.175 1307.025 3196.505 ;
        RECT 1306.710 856.625 1307.010 3196.175 ;
        RECT 1306.695 856.295 1307.025 856.625 ;
        RECT 2656.335 850.855 2656.665 851.185 ;
        RECT 2656.350 849.825 2656.650 850.855 ;
        RECT 2656.335 849.495 2656.665 849.825 ;
        RECT 2752.935 849.495 2753.265 849.825 ;
        RECT 2752.950 848.465 2753.250 849.495 ;
        RECT 2752.935 848.135 2753.265 848.465 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1340.970 3196.580 1341.290 3196.640 ;
        RECT 2901.290 3196.580 2901.610 3196.640 ;
        RECT 1340.970 3196.440 2901.610 3196.580 ;
        RECT 1340.970 3196.380 1341.290 3196.440 ;
        RECT 2901.290 3196.380 2901.610 3196.440 ;
      LAYER via ;
        RECT 1341.000 3196.380 1341.260 3196.640 ;
        RECT 2901.320 3196.380 2901.580 3196.640 ;
      LAYER met2 ;
        RECT 1339.080 3196.410 1339.360 3200.000 ;
        RECT 1341.000 3196.410 1341.260 3196.670 ;
        RECT 1339.080 3196.350 1341.260 3196.410 ;
        RECT 2901.320 3196.350 2901.580 3196.670 ;
        RECT 1339.080 3196.270 1341.200 3196.350 ;
        RECT 1339.080 3196.000 1339.360 3196.270 ;
        RECT 2901.380 1085.125 2901.520 3196.350 ;
        RECT 2901.310 1084.755 2901.590 1085.125 ;
      LAYER via2 ;
        RECT 2901.310 1084.800 2901.590 1085.080 ;
      LAYER met3 ;
        RECT 2901.285 1085.090 2901.615 1085.105 ;
        RECT 2917.600 1085.090 2924.800 1085.540 ;
        RECT 2901.285 1084.790 2924.800 1085.090 ;
        RECT 2901.285 1084.775 2901.615 1084.790 ;
        RECT 2917.600 1084.340 2924.800 1084.790 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1379.610 3196.920 1379.930 3196.980 ;
        RECT 2902.670 3196.920 2902.990 3196.980 ;
        RECT 1379.610 3196.780 2902.990 3196.920 ;
        RECT 1379.610 3196.720 1379.930 3196.780 ;
        RECT 2902.670 3196.720 2902.990 3196.780 ;
      LAYER via ;
        RECT 1379.640 3196.720 1379.900 3196.980 ;
        RECT 2902.700 3196.720 2902.960 3196.980 ;
      LAYER met2 ;
        RECT 1378.640 3197.090 1378.920 3200.000 ;
        RECT 1378.640 3197.010 1379.840 3197.090 ;
        RECT 1378.640 3196.950 1379.900 3197.010 ;
        RECT 1378.640 3196.000 1378.920 3196.950 ;
        RECT 1379.640 3196.690 1379.900 3196.950 ;
        RECT 2902.700 3196.690 2902.960 3197.010 ;
        RECT 2902.760 1319.725 2902.900 3196.690 ;
        RECT 2902.690 1319.355 2902.970 1319.725 ;
      LAYER via2 ;
        RECT 2902.690 1319.400 2902.970 1319.680 ;
      LAYER met3 ;
        RECT 2902.665 1319.690 2902.995 1319.705 ;
        RECT 2917.600 1319.690 2924.800 1320.140 ;
        RECT 2902.665 1319.390 2924.800 1319.690 ;
        RECT 2902.665 1319.375 2902.995 1319.390 ;
        RECT 2917.600 1318.940 2924.800 1319.390 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1420.090 3197.260 1420.410 3197.320 ;
        RECT 2903.130 3197.260 2903.450 3197.320 ;
        RECT 1420.090 3197.120 2903.450 3197.260 ;
        RECT 1420.090 3197.060 1420.410 3197.120 ;
        RECT 2903.130 3197.060 2903.450 3197.120 ;
      LAYER via ;
        RECT 1420.120 3197.060 1420.380 3197.320 ;
        RECT 2903.160 3197.060 2903.420 3197.320 ;
      LAYER met2 ;
        RECT 1418.200 3197.090 1418.480 3200.000 ;
        RECT 1420.120 3197.090 1420.380 3197.350 ;
        RECT 1418.200 3197.030 1420.380 3197.090 ;
        RECT 2903.160 3197.030 2903.420 3197.350 ;
        RECT 1418.200 3196.950 1420.320 3197.030 ;
        RECT 1418.200 3196.000 1418.480 3196.950 ;
        RECT 2903.220 1554.325 2903.360 3197.030 ;
        RECT 2903.150 1553.955 2903.430 1554.325 ;
      LAYER via2 ;
        RECT 2903.150 1554.000 2903.430 1554.280 ;
      LAYER met3 ;
        RECT 2903.125 1554.290 2903.455 1554.305 ;
        RECT 2917.600 1554.290 2924.800 1554.740 ;
        RECT 2903.125 1553.990 2924.800 1554.290 ;
        RECT 2903.125 1553.975 2903.455 1553.990 ;
        RECT 2917.600 1553.540 2924.800 1553.990 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1458.730 3197.600 1459.050 3197.660 ;
        RECT 2903.590 3197.600 2903.910 3197.660 ;
        RECT 1458.730 3197.460 2903.910 3197.600 ;
        RECT 1458.730 3197.400 1459.050 3197.460 ;
        RECT 2903.590 3197.400 2903.910 3197.460 ;
      LAYER via ;
        RECT 1458.760 3197.400 1459.020 3197.660 ;
        RECT 2903.620 3197.400 2903.880 3197.660 ;
      LAYER met2 ;
        RECT 1457.300 3197.770 1457.580 3200.000 ;
        RECT 1457.300 3197.690 1458.960 3197.770 ;
        RECT 1457.300 3197.630 1459.020 3197.690 ;
        RECT 1457.300 3196.000 1457.580 3197.630 ;
        RECT 1458.760 3197.370 1459.020 3197.630 ;
        RECT 2903.620 3197.370 2903.880 3197.690 ;
        RECT 2903.680 1789.605 2903.820 3197.370 ;
        RECT 2903.610 1789.235 2903.890 1789.605 ;
      LAYER via2 ;
        RECT 2903.610 1789.280 2903.890 1789.560 ;
      LAYER met3 ;
        RECT 2903.585 1789.570 2903.915 1789.585 ;
        RECT 2917.600 1789.570 2924.800 1790.020 ;
        RECT 2903.585 1789.270 2924.800 1789.570 ;
        RECT 2903.585 1789.255 2903.915 1789.270 ;
        RECT 2917.600 1788.820 2924.800 1789.270 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1497.370 3197.940 1497.690 3198.000 ;
        RECT 2904.050 3197.940 2904.370 3198.000 ;
        RECT 1497.370 3197.800 2904.370 3197.940 ;
        RECT 1497.370 3197.740 1497.690 3197.800 ;
        RECT 2904.050 3197.740 2904.370 3197.800 ;
      LAYER via ;
        RECT 1497.400 3197.740 1497.660 3198.000 ;
        RECT 2904.080 3197.740 2904.340 3198.000 ;
      LAYER met2 ;
        RECT 1496.860 3197.770 1497.140 3200.000 ;
        RECT 1497.400 3197.770 1497.660 3198.030 ;
        RECT 1496.860 3197.710 1497.660 3197.770 ;
        RECT 2904.080 3197.710 2904.340 3198.030 ;
        RECT 1496.860 3197.630 1497.600 3197.710 ;
        RECT 1496.860 3196.000 1497.140 3197.630 ;
        RECT 2904.140 2024.205 2904.280 3197.710 ;
        RECT 2904.070 2023.835 2904.350 2024.205 ;
      LAYER via2 ;
        RECT 2904.070 2023.880 2904.350 2024.160 ;
      LAYER met3 ;
        RECT 2904.045 2024.170 2904.375 2024.185 ;
        RECT 2917.600 2024.170 2924.800 2024.620 ;
        RECT 2904.045 2023.870 2924.800 2024.170 ;
        RECT 2904.045 2023.855 2904.375 2023.870 ;
        RECT 2917.600 2023.420 2924.800 2023.870 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1537.850 3198.280 1538.170 3198.340 ;
        RECT 2904.510 3198.280 2904.830 3198.340 ;
        RECT 1537.850 3198.140 2904.830 3198.280 ;
        RECT 1537.850 3198.080 1538.170 3198.140 ;
        RECT 2904.510 3198.080 2904.830 3198.140 ;
      LAYER via ;
        RECT 1537.880 3198.080 1538.140 3198.340 ;
        RECT 2904.540 3198.080 2904.800 3198.340 ;
      LAYER met2 ;
        RECT 1536.420 3198.450 1536.700 3200.000 ;
        RECT 1536.420 3198.370 1538.080 3198.450 ;
        RECT 1536.420 3198.310 1538.140 3198.370 ;
        RECT 1536.420 3196.000 1536.700 3198.310 ;
        RECT 1537.880 3198.050 1538.140 3198.310 ;
        RECT 2904.540 3198.050 2904.800 3198.370 ;
        RECT 2904.600 2258.805 2904.740 3198.050 ;
        RECT 2904.530 2258.435 2904.810 2258.805 ;
      LAYER via2 ;
        RECT 2904.530 2258.480 2904.810 2258.760 ;
      LAYER met3 ;
        RECT 2904.505 2258.770 2904.835 2258.785 ;
        RECT 2917.600 2258.770 2924.800 2259.220 ;
        RECT 2904.505 2258.470 2924.800 2258.770 ;
        RECT 2904.505 2258.455 2904.835 2258.470 ;
        RECT 2917.600 2258.020 2924.800 2258.470 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1470.305 1628.345 1470.475 1676.455 ;
        RECT 1470.765 1256.045 1470.935 1304.155 ;
        RECT 1470.765 421.005 1470.935 468.435 ;
        RECT 1469.845 59.245 1470.015 62.475 ;
      LAYER mcon ;
        RECT 1470.305 1676.285 1470.475 1676.455 ;
        RECT 1470.765 1303.985 1470.935 1304.155 ;
        RECT 1470.765 468.265 1470.935 468.435 ;
        RECT 1469.845 62.305 1470.015 62.475 ;
      LAYER met1 ;
        RECT 1470.245 1676.440 1470.535 1676.485 ;
        RECT 1472.530 1676.440 1472.850 1676.500 ;
        RECT 1470.245 1676.300 1472.850 1676.440 ;
        RECT 1470.245 1676.255 1470.535 1676.300 ;
        RECT 1472.530 1676.240 1472.850 1676.300 ;
        RECT 1470.230 1628.500 1470.550 1628.560 ;
        RECT 1470.035 1628.360 1470.550 1628.500 ;
        RECT 1470.230 1628.300 1470.550 1628.360 ;
        RECT 1470.690 1580.220 1471.010 1580.280 ;
        RECT 1471.610 1580.220 1471.930 1580.280 ;
        RECT 1470.690 1580.080 1471.930 1580.220 ;
        RECT 1470.690 1580.020 1471.010 1580.080 ;
        RECT 1471.610 1580.020 1471.930 1580.080 ;
        RECT 1470.690 1559.620 1471.010 1559.880 ;
        RECT 1470.780 1559.200 1470.920 1559.620 ;
        RECT 1470.690 1558.940 1471.010 1559.200 ;
        RECT 1470.690 1365.820 1471.010 1366.080 ;
        RECT 1470.780 1365.400 1470.920 1365.820 ;
        RECT 1470.690 1365.140 1471.010 1365.400 ;
        RECT 1470.690 1304.140 1471.010 1304.200 ;
        RECT 1470.495 1304.000 1471.010 1304.140 ;
        RECT 1470.690 1303.940 1471.010 1304.000 ;
        RECT 1470.690 1256.200 1471.010 1256.260 ;
        RECT 1470.495 1256.060 1471.010 1256.200 ;
        RECT 1470.690 1256.000 1471.010 1256.060 ;
        RECT 1469.770 1159.300 1470.090 1159.360 ;
        RECT 1470.690 1159.300 1471.010 1159.360 ;
        RECT 1469.770 1159.160 1471.010 1159.300 ;
        RECT 1469.770 1159.100 1470.090 1159.160 ;
        RECT 1470.690 1159.100 1471.010 1159.160 ;
        RECT 1470.690 1000.520 1471.010 1000.580 ;
        RECT 1471.150 1000.520 1471.470 1000.580 ;
        RECT 1470.690 1000.380 1471.470 1000.520 ;
        RECT 1470.690 1000.320 1471.010 1000.380 ;
        RECT 1471.150 1000.320 1471.470 1000.380 ;
        RECT 1471.150 869.960 1471.470 870.020 ;
        RECT 1470.780 869.820 1471.470 869.960 ;
        RECT 1470.780 869.340 1470.920 869.820 ;
        RECT 1471.150 869.760 1471.470 869.820 ;
        RECT 1470.690 869.080 1471.010 869.340 ;
        RECT 1470.230 724.440 1470.550 724.500 ;
        RECT 1471.150 724.440 1471.470 724.500 ;
        RECT 1470.230 724.300 1471.470 724.440 ;
        RECT 1470.230 724.240 1470.550 724.300 ;
        RECT 1471.150 724.240 1471.470 724.300 ;
        RECT 1470.230 572.940 1470.550 573.200 ;
        RECT 1470.320 572.800 1470.460 572.940 ;
        RECT 1470.690 572.800 1471.010 572.860 ;
        RECT 1470.320 572.660 1471.010 572.800 ;
        RECT 1470.690 572.600 1471.010 572.660 ;
        RECT 1470.690 548.460 1471.010 548.720 ;
        RECT 1470.780 548.040 1470.920 548.460 ;
        RECT 1470.690 547.780 1471.010 548.040 ;
        RECT 1470.690 468.900 1471.010 469.160 ;
        RECT 1470.780 468.465 1470.920 468.900 ;
        RECT 1470.705 468.235 1470.995 468.465 ;
        RECT 1470.690 421.160 1471.010 421.220 ;
        RECT 1470.495 421.020 1471.010 421.160 ;
        RECT 1470.690 420.960 1471.010 421.020 ;
        RECT 1470.230 362.340 1470.550 362.400 ;
        RECT 1471.150 362.340 1471.470 362.400 ;
        RECT 1470.230 362.200 1471.470 362.340 ;
        RECT 1470.230 362.140 1470.550 362.200 ;
        RECT 1471.150 362.140 1471.470 362.200 ;
        RECT 1469.770 331.060 1470.090 331.120 ;
        RECT 1471.150 331.060 1471.470 331.120 ;
        RECT 1469.770 330.920 1471.470 331.060 ;
        RECT 1469.770 330.860 1470.090 330.920 ;
        RECT 1471.150 330.860 1471.470 330.920 ;
        RECT 1469.770 144.740 1470.090 144.800 ;
        RECT 1470.690 144.740 1471.010 144.800 ;
        RECT 1469.770 144.600 1471.010 144.740 ;
        RECT 1469.770 144.540 1470.090 144.600 ;
        RECT 1470.690 144.540 1471.010 144.600 ;
        RECT 1469.770 62.460 1470.090 62.520 ;
        RECT 1469.575 62.320 1470.090 62.460 ;
        RECT 1469.770 62.260 1470.090 62.320 ;
        RECT 634.410 59.400 634.730 59.460 ;
        RECT 1469.785 59.400 1470.075 59.445 ;
        RECT 634.410 59.260 1470.075 59.400 ;
        RECT 634.410 59.200 634.730 59.260 ;
        RECT 1469.785 59.215 1470.075 59.260 ;
      LAYER via ;
        RECT 1472.560 1676.240 1472.820 1676.500 ;
        RECT 1470.260 1628.300 1470.520 1628.560 ;
        RECT 1470.720 1580.020 1470.980 1580.280 ;
        RECT 1471.640 1580.020 1471.900 1580.280 ;
        RECT 1470.720 1559.620 1470.980 1559.880 ;
        RECT 1470.720 1558.940 1470.980 1559.200 ;
        RECT 1470.720 1365.820 1470.980 1366.080 ;
        RECT 1470.720 1365.140 1470.980 1365.400 ;
        RECT 1470.720 1303.940 1470.980 1304.200 ;
        RECT 1470.720 1256.000 1470.980 1256.260 ;
        RECT 1469.800 1159.100 1470.060 1159.360 ;
        RECT 1470.720 1159.100 1470.980 1159.360 ;
        RECT 1470.720 1000.320 1470.980 1000.580 ;
        RECT 1471.180 1000.320 1471.440 1000.580 ;
        RECT 1471.180 869.760 1471.440 870.020 ;
        RECT 1470.720 869.080 1470.980 869.340 ;
        RECT 1470.260 724.240 1470.520 724.500 ;
        RECT 1471.180 724.240 1471.440 724.500 ;
        RECT 1470.260 572.940 1470.520 573.200 ;
        RECT 1470.720 572.600 1470.980 572.860 ;
        RECT 1470.720 548.460 1470.980 548.720 ;
        RECT 1470.720 547.780 1470.980 548.040 ;
        RECT 1470.720 468.900 1470.980 469.160 ;
        RECT 1470.720 420.960 1470.980 421.220 ;
        RECT 1470.260 362.140 1470.520 362.400 ;
        RECT 1471.180 362.140 1471.440 362.400 ;
        RECT 1469.800 330.860 1470.060 331.120 ;
        RECT 1471.180 330.860 1471.440 331.120 ;
        RECT 1469.800 144.540 1470.060 144.800 ;
        RECT 1470.720 144.540 1470.980 144.800 ;
        RECT 1469.800 62.260 1470.060 62.520 ;
        RECT 634.440 59.200 634.700 59.460 ;
      LAYER met2 ;
        RECT 1474.320 1701.090 1474.600 1704.000 ;
        RECT 1472.620 1700.950 1474.600 1701.090 ;
        RECT 1472.620 1676.530 1472.760 1700.950 ;
        RECT 1474.320 1700.000 1474.600 1700.950 ;
        RECT 1472.560 1676.210 1472.820 1676.530 ;
        RECT 1470.260 1628.330 1470.520 1628.590 ;
        RECT 1470.710 1628.330 1470.990 1628.445 ;
        RECT 1470.260 1628.270 1470.990 1628.330 ;
        RECT 1470.320 1628.190 1470.990 1628.270 ;
        RECT 1470.710 1628.075 1470.990 1628.190 ;
        RECT 1471.630 1628.075 1471.910 1628.445 ;
        RECT 1471.700 1580.310 1471.840 1628.075 ;
        RECT 1470.720 1579.990 1470.980 1580.310 ;
        RECT 1471.640 1579.990 1471.900 1580.310 ;
        RECT 1470.780 1559.910 1470.920 1579.990 ;
        RECT 1470.720 1559.590 1470.980 1559.910 ;
        RECT 1470.720 1558.910 1470.980 1559.230 ;
        RECT 1470.780 1366.110 1470.920 1558.910 ;
        RECT 1470.720 1365.790 1470.980 1366.110 ;
        RECT 1470.720 1365.110 1470.980 1365.430 ;
        RECT 1470.780 1304.230 1470.920 1365.110 ;
        RECT 1470.720 1303.910 1470.980 1304.230 ;
        RECT 1470.720 1255.970 1470.980 1256.290 ;
        RECT 1470.780 1207.525 1470.920 1255.970 ;
        RECT 1469.790 1207.155 1470.070 1207.525 ;
        RECT 1470.710 1207.155 1470.990 1207.525 ;
        RECT 1469.860 1159.390 1470.000 1207.155 ;
        RECT 1469.800 1159.070 1470.060 1159.390 ;
        RECT 1470.720 1159.070 1470.980 1159.390 ;
        RECT 1470.780 1110.965 1470.920 1159.070 ;
        RECT 1469.790 1110.595 1470.070 1110.965 ;
        RECT 1470.710 1110.595 1470.990 1110.965 ;
        RECT 1469.860 1091.810 1470.000 1110.595 ;
        RECT 1469.860 1091.670 1471.380 1091.810 ;
        RECT 1471.240 1055.770 1471.380 1091.670 ;
        RECT 1470.780 1055.630 1471.380 1055.770 ;
        RECT 1470.780 1000.610 1470.920 1055.630 ;
        RECT 1470.720 1000.290 1470.980 1000.610 ;
        RECT 1471.180 1000.290 1471.440 1000.610 ;
        RECT 1471.240 870.050 1471.380 1000.290 ;
        RECT 1471.180 869.730 1471.440 870.050 ;
        RECT 1470.720 869.050 1470.980 869.370 ;
        RECT 1470.780 844.970 1470.920 869.050 ;
        RECT 1470.320 844.830 1470.920 844.970 ;
        RECT 1470.320 787.170 1470.460 844.830 ;
        RECT 1469.860 787.030 1470.460 787.170 ;
        RECT 1469.860 786.490 1470.000 787.030 ;
        RECT 1469.860 786.350 1470.460 786.490 ;
        RECT 1470.320 724.530 1470.460 786.350 ;
        RECT 1470.260 724.210 1470.520 724.530 ;
        RECT 1471.180 724.210 1471.440 724.530 ;
        RECT 1471.240 699.450 1471.380 724.210 ;
        RECT 1470.780 699.310 1471.380 699.450 ;
        RECT 1470.780 628.845 1470.920 699.310 ;
        RECT 1470.710 628.475 1470.990 628.845 ;
        RECT 1470.250 627.795 1470.530 628.165 ;
        RECT 1470.320 573.230 1470.460 627.795 ;
        RECT 1470.260 572.910 1470.520 573.230 ;
        RECT 1470.720 572.570 1470.980 572.890 ;
        RECT 1470.780 548.750 1470.920 572.570 ;
        RECT 1470.720 548.430 1470.980 548.750 ;
        RECT 1470.720 547.750 1470.980 548.070 ;
        RECT 1470.780 494.090 1470.920 547.750 ;
        RECT 1470.320 493.950 1470.920 494.090 ;
        RECT 1470.320 469.610 1470.460 493.950 ;
        RECT 1470.320 469.470 1470.920 469.610 ;
        RECT 1470.780 469.190 1470.920 469.470 ;
        RECT 1470.720 468.870 1470.980 469.190 ;
        RECT 1470.720 420.930 1470.980 421.250 ;
        RECT 1470.780 386.820 1470.920 420.930 ;
        RECT 1470.780 386.680 1471.380 386.820 ;
        RECT 1471.240 385.970 1471.380 386.680 ;
        RECT 1470.320 385.830 1471.380 385.970 ;
        RECT 1470.320 362.430 1470.460 385.830 ;
        RECT 1470.260 362.110 1470.520 362.430 ;
        RECT 1471.180 362.110 1471.440 362.430 ;
        RECT 1471.240 331.150 1471.380 362.110 ;
        RECT 1469.800 330.830 1470.060 331.150 ;
        RECT 1471.180 330.830 1471.440 331.150 ;
        RECT 1469.860 258.810 1470.000 330.830 ;
        RECT 1469.860 258.670 1470.460 258.810 ;
        RECT 1470.320 210.530 1470.460 258.670 ;
        RECT 1470.320 210.390 1471.380 210.530 ;
        RECT 1471.240 206.450 1471.380 210.390 ;
        RECT 1470.780 206.310 1471.380 206.450 ;
        RECT 1470.780 144.830 1470.920 206.310 ;
        RECT 1469.800 144.510 1470.060 144.830 ;
        RECT 1470.720 144.510 1470.980 144.830 ;
        RECT 1469.860 62.550 1470.000 144.510 ;
        RECT 1469.800 62.230 1470.060 62.550 ;
        RECT 634.440 59.170 634.700 59.490 ;
        RECT 634.500 17.410 634.640 59.170 ;
        RECT 633.120 17.270 634.640 17.410 ;
        RECT 633.120 2.400 633.260 17.270 ;
        RECT 632.910 -4.800 633.470 2.400 ;
      LAYER via2 ;
        RECT 1470.710 1628.120 1470.990 1628.400 ;
        RECT 1471.630 1628.120 1471.910 1628.400 ;
        RECT 1469.790 1207.200 1470.070 1207.480 ;
        RECT 1470.710 1207.200 1470.990 1207.480 ;
        RECT 1469.790 1110.640 1470.070 1110.920 ;
        RECT 1470.710 1110.640 1470.990 1110.920 ;
        RECT 1470.710 628.520 1470.990 628.800 ;
        RECT 1470.250 627.840 1470.530 628.120 ;
      LAYER met3 ;
        RECT 1470.685 1628.410 1471.015 1628.425 ;
        RECT 1471.605 1628.410 1471.935 1628.425 ;
        RECT 1470.685 1628.110 1471.935 1628.410 ;
        RECT 1470.685 1628.095 1471.015 1628.110 ;
        RECT 1471.605 1628.095 1471.935 1628.110 ;
        RECT 1469.765 1207.490 1470.095 1207.505 ;
        RECT 1470.685 1207.490 1471.015 1207.505 ;
        RECT 1469.765 1207.190 1471.015 1207.490 ;
        RECT 1469.765 1207.175 1470.095 1207.190 ;
        RECT 1470.685 1207.175 1471.015 1207.190 ;
        RECT 1469.765 1110.930 1470.095 1110.945 ;
        RECT 1470.685 1110.930 1471.015 1110.945 ;
        RECT 1469.765 1110.630 1471.015 1110.930 ;
        RECT 1469.765 1110.615 1470.095 1110.630 ;
        RECT 1470.685 1110.615 1471.015 1110.630 ;
        RECT 1470.685 628.810 1471.015 628.825 ;
        RECT 1470.470 628.495 1471.015 628.810 ;
        RECT 1470.470 628.145 1470.770 628.495 ;
        RECT 1470.225 627.830 1470.770 628.145 ;
        RECT 1470.225 627.815 1470.555 627.830 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2392.530 1684.600 2392.850 1684.660 ;
        RECT 2415.990 1684.600 2416.310 1684.660 ;
        RECT 2392.530 1684.460 2416.310 1684.600 ;
        RECT 2392.530 1684.400 2392.850 1684.460 ;
        RECT 2415.990 1684.400 2416.310 1684.460 ;
      LAYER via ;
        RECT 2392.560 1684.400 2392.820 1684.660 ;
        RECT 2416.020 1684.400 2416.280 1684.660 ;
      LAYER met2 ;
        RECT 2392.480 1700.000 2392.760 1704.000 ;
        RECT 2392.620 1684.690 2392.760 1700.000 ;
        RECT 2392.560 1684.370 2392.820 1684.690 ;
        RECT 2416.020 1684.370 2416.280 1684.690 ;
        RECT 2416.080 3.130 2416.220 1684.370 ;
        RECT 2416.080 2.990 2417.600 3.130 ;
        RECT 2417.460 2.400 2417.600 2.990 ;
        RECT 2417.250 -4.800 2417.810 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2401.730 1683.920 2402.050 1683.980 ;
        RECT 2407.710 1683.920 2408.030 1683.980 ;
        RECT 2401.730 1683.780 2408.030 1683.920 ;
        RECT 2401.730 1683.720 2402.050 1683.780 ;
        RECT 2407.710 1683.720 2408.030 1683.780 ;
        RECT 2407.710 16.560 2408.030 16.620 ;
        RECT 2434.850 16.560 2435.170 16.620 ;
        RECT 2407.710 16.420 2435.170 16.560 ;
        RECT 2407.710 16.360 2408.030 16.420 ;
        RECT 2434.850 16.360 2435.170 16.420 ;
      LAYER via ;
        RECT 2401.760 1683.720 2402.020 1683.980 ;
        RECT 2407.740 1683.720 2408.000 1683.980 ;
        RECT 2407.740 16.360 2408.000 16.620 ;
        RECT 2434.880 16.360 2435.140 16.620 ;
      LAYER met2 ;
        RECT 2401.680 1700.000 2401.960 1704.000 ;
        RECT 2401.820 1684.010 2401.960 1700.000 ;
        RECT 2401.760 1683.690 2402.020 1684.010 ;
        RECT 2407.740 1683.690 2408.000 1684.010 ;
        RECT 2407.800 16.650 2407.940 1683.690 ;
        RECT 2407.740 16.330 2408.000 16.650 ;
        RECT 2434.880 16.330 2435.140 16.650 ;
        RECT 2434.940 2.400 2435.080 16.330 ;
        RECT 2434.730 -4.800 2435.290 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2410.930 1685.280 2411.250 1685.340 ;
        RECT 2414.150 1685.280 2414.470 1685.340 ;
        RECT 2410.930 1685.140 2414.470 1685.280 ;
        RECT 2410.930 1685.080 2411.250 1685.140 ;
        RECT 2414.150 1685.080 2414.470 1685.140 ;
        RECT 2414.150 19.280 2414.470 19.340 ;
        RECT 2452.790 19.280 2453.110 19.340 ;
        RECT 2414.150 19.140 2453.110 19.280 ;
        RECT 2414.150 19.080 2414.470 19.140 ;
        RECT 2452.790 19.080 2453.110 19.140 ;
      LAYER via ;
        RECT 2410.960 1685.080 2411.220 1685.340 ;
        RECT 2414.180 1685.080 2414.440 1685.340 ;
        RECT 2414.180 19.080 2414.440 19.340 ;
        RECT 2452.820 19.080 2453.080 19.340 ;
      LAYER met2 ;
        RECT 2410.880 1700.000 2411.160 1704.000 ;
        RECT 2411.020 1685.370 2411.160 1700.000 ;
        RECT 2410.960 1685.050 2411.220 1685.370 ;
        RECT 2414.180 1685.050 2414.440 1685.370 ;
        RECT 2414.240 19.370 2414.380 1685.050 ;
        RECT 2414.180 19.050 2414.440 19.370 ;
        RECT 2452.820 19.050 2453.080 19.370 ;
        RECT 2452.880 2.400 2453.020 19.050 ;
        RECT 2452.670 -4.800 2453.230 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2421.050 17.920 2421.370 17.980 ;
        RECT 2470.730 17.920 2471.050 17.980 ;
        RECT 2421.050 17.780 2471.050 17.920 ;
        RECT 2421.050 17.720 2421.370 17.780 ;
        RECT 2470.730 17.720 2471.050 17.780 ;
      LAYER via ;
        RECT 2421.080 17.720 2421.340 17.980 ;
        RECT 2470.760 17.720 2471.020 17.980 ;
      LAYER met2 ;
        RECT 2420.080 1700.410 2420.360 1704.000 ;
        RECT 2420.080 1700.270 2421.280 1700.410 ;
        RECT 2420.080 1700.000 2420.360 1700.270 ;
        RECT 2421.140 18.010 2421.280 1700.270 ;
        RECT 2421.080 17.690 2421.340 18.010 ;
        RECT 2470.760 17.690 2471.020 18.010 ;
        RECT 2470.820 2.400 2470.960 17.690 ;
        RECT 2470.610 -4.800 2471.170 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2429.330 1688.340 2429.650 1688.400 ;
        RECT 2445.890 1688.340 2446.210 1688.400 ;
        RECT 2429.330 1688.200 2446.210 1688.340 ;
        RECT 2429.330 1688.140 2429.650 1688.200 ;
        RECT 2445.890 1688.140 2446.210 1688.200 ;
        RECT 2445.890 18.940 2446.210 19.000 ;
        RECT 2488.670 18.940 2488.990 19.000 ;
        RECT 2445.890 18.800 2488.990 18.940 ;
        RECT 2445.890 18.740 2446.210 18.800 ;
        RECT 2488.670 18.740 2488.990 18.800 ;
      LAYER via ;
        RECT 2429.360 1688.140 2429.620 1688.400 ;
        RECT 2445.920 1688.140 2446.180 1688.400 ;
        RECT 2445.920 18.740 2446.180 19.000 ;
        RECT 2488.700 18.740 2488.960 19.000 ;
      LAYER met2 ;
        RECT 2429.280 1700.000 2429.560 1704.000 ;
        RECT 2429.420 1688.430 2429.560 1700.000 ;
        RECT 2429.360 1688.110 2429.620 1688.430 ;
        RECT 2445.920 1688.110 2446.180 1688.430 ;
        RECT 2445.980 19.030 2446.120 1688.110 ;
        RECT 2445.920 18.710 2446.180 19.030 ;
        RECT 2488.700 18.710 2488.960 19.030 ;
        RECT 2488.760 2.400 2488.900 18.710 ;
        RECT 2488.550 -4.800 2489.110 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2441.750 17.240 2442.070 17.300 ;
        RECT 2506.150 17.240 2506.470 17.300 ;
        RECT 2441.750 17.100 2506.470 17.240 ;
        RECT 2441.750 17.040 2442.070 17.100 ;
        RECT 2506.150 17.040 2506.470 17.100 ;
      LAYER via ;
        RECT 2441.780 17.040 2442.040 17.300 ;
        RECT 2506.180 17.040 2506.440 17.300 ;
      LAYER met2 ;
        RECT 2438.480 1701.090 2438.760 1704.000 ;
        RECT 2438.480 1700.950 2441.520 1701.090 ;
        RECT 2438.480 1700.000 2438.760 1700.950 ;
        RECT 2441.380 1688.850 2441.520 1700.950 ;
        RECT 2441.380 1688.710 2441.980 1688.850 ;
        RECT 2441.840 17.330 2441.980 1688.710 ;
        RECT 2441.780 17.010 2442.040 17.330 ;
        RECT 2506.180 17.010 2506.440 17.330 ;
        RECT 2506.240 2.400 2506.380 17.010 ;
        RECT 2506.030 -4.800 2506.590 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2449.110 16.220 2449.430 16.280 ;
        RECT 2524.090 16.220 2524.410 16.280 ;
        RECT 2449.110 16.080 2524.410 16.220 ;
        RECT 2449.110 16.020 2449.430 16.080 ;
        RECT 2524.090 16.020 2524.410 16.080 ;
      LAYER via ;
        RECT 2449.140 16.020 2449.400 16.280 ;
        RECT 2524.120 16.020 2524.380 16.280 ;
      LAYER met2 ;
        RECT 2447.680 1700.410 2447.960 1704.000 ;
        RECT 2447.680 1700.270 2449.340 1700.410 ;
        RECT 2447.680 1700.000 2447.960 1700.270 ;
        RECT 2449.200 16.310 2449.340 1700.270 ;
        RECT 2449.140 15.990 2449.400 16.310 ;
        RECT 2524.120 15.990 2524.380 16.310 ;
        RECT 2524.180 2.400 2524.320 15.990 ;
        RECT 2523.970 -4.800 2524.530 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2456.930 1688.340 2457.250 1688.400 ;
        RECT 2462.450 1688.340 2462.770 1688.400 ;
        RECT 2456.930 1688.200 2462.770 1688.340 ;
        RECT 2456.930 1688.140 2457.250 1688.200 ;
        RECT 2462.450 1688.140 2462.770 1688.200 ;
        RECT 2462.450 16.900 2462.770 16.960 ;
        RECT 2542.030 16.900 2542.350 16.960 ;
        RECT 2462.450 16.760 2542.350 16.900 ;
        RECT 2462.450 16.700 2462.770 16.760 ;
        RECT 2542.030 16.700 2542.350 16.760 ;
      LAYER via ;
        RECT 2456.960 1688.140 2457.220 1688.400 ;
        RECT 2462.480 1688.140 2462.740 1688.400 ;
        RECT 2462.480 16.700 2462.740 16.960 ;
        RECT 2542.060 16.700 2542.320 16.960 ;
      LAYER met2 ;
        RECT 2456.880 1700.000 2457.160 1704.000 ;
        RECT 2457.020 1688.430 2457.160 1700.000 ;
        RECT 2456.960 1688.110 2457.220 1688.430 ;
        RECT 2462.480 1688.110 2462.740 1688.430 ;
        RECT 2462.540 16.990 2462.680 1688.110 ;
        RECT 2462.480 16.670 2462.740 16.990 ;
        RECT 2542.060 16.670 2542.320 16.990 ;
        RECT 2542.120 2.400 2542.260 16.670 ;
        RECT 2541.910 -4.800 2542.470 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2469.350 19.960 2469.670 20.020 ;
        RECT 2559.970 19.960 2560.290 20.020 ;
        RECT 2469.350 19.820 2560.290 19.960 ;
        RECT 2469.350 19.760 2469.670 19.820 ;
        RECT 2559.970 19.760 2560.290 19.820 ;
      LAYER via ;
        RECT 2469.380 19.760 2469.640 20.020 ;
        RECT 2560.000 19.760 2560.260 20.020 ;
      LAYER met2 ;
        RECT 2466.080 1701.090 2466.360 1704.000 ;
        RECT 2466.080 1700.950 2469.120 1701.090 ;
        RECT 2466.080 1700.000 2466.360 1700.950 ;
        RECT 2468.980 1688.680 2469.120 1700.950 ;
        RECT 2468.980 1688.540 2469.580 1688.680 ;
        RECT 2469.440 20.050 2469.580 1688.540 ;
        RECT 2469.380 19.730 2469.640 20.050 ;
        RECT 2560.000 19.730 2560.260 20.050 ;
        RECT 2560.060 2.400 2560.200 19.730 ;
        RECT 2559.850 -4.800 2560.410 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2475.330 1688.340 2475.650 1688.400 ;
        RECT 2480.390 1688.340 2480.710 1688.400 ;
        RECT 2475.330 1688.200 2480.710 1688.340 ;
        RECT 2475.330 1688.140 2475.650 1688.200 ;
        RECT 2480.390 1688.140 2480.710 1688.200 ;
        RECT 2480.390 19.620 2480.710 19.680 ;
        RECT 2577.910 19.620 2578.230 19.680 ;
        RECT 2480.390 19.480 2578.230 19.620 ;
        RECT 2480.390 19.420 2480.710 19.480 ;
        RECT 2577.910 19.420 2578.230 19.480 ;
      LAYER via ;
        RECT 2475.360 1688.140 2475.620 1688.400 ;
        RECT 2480.420 1688.140 2480.680 1688.400 ;
        RECT 2480.420 19.420 2480.680 19.680 ;
        RECT 2577.940 19.420 2578.200 19.680 ;
      LAYER met2 ;
        RECT 2475.280 1700.000 2475.560 1704.000 ;
        RECT 2475.420 1688.430 2475.560 1700.000 ;
        RECT 2475.360 1688.110 2475.620 1688.430 ;
        RECT 2480.420 1688.110 2480.680 1688.430 ;
        RECT 2480.480 19.710 2480.620 1688.110 ;
        RECT 2480.420 19.390 2480.680 19.710 ;
        RECT 2577.940 19.390 2578.200 19.710 ;
        RECT 2578.000 2.400 2578.140 19.390 ;
        RECT 2577.790 -4.800 2578.350 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 813.810 60.080 814.130 60.140 ;
        RECT 1566.830 60.080 1567.150 60.140 ;
        RECT 813.810 59.940 1567.150 60.080 ;
        RECT 813.810 59.880 814.130 59.940 ;
        RECT 1566.830 59.880 1567.150 59.940 ;
      LAYER via ;
        RECT 813.840 59.880 814.100 60.140 ;
        RECT 1566.860 59.880 1567.120 60.140 ;
      LAYER met2 ;
        RECT 1566.320 1700.410 1566.600 1704.000 ;
        RECT 1566.320 1700.270 1567.060 1700.410 ;
        RECT 1566.320 1700.000 1566.600 1700.270 ;
        RECT 1566.920 60.170 1567.060 1700.270 ;
        RECT 813.840 59.850 814.100 60.170 ;
        RECT 1566.860 59.850 1567.120 60.170 ;
        RECT 813.900 16.730 814.040 59.850 ;
        RECT 811.600 16.590 814.040 16.730 ;
        RECT 811.600 2.400 811.740 16.590 ;
        RECT 811.390 -4.800 811.950 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2484.530 1688.340 2484.850 1688.400 ;
        RECT 2494.190 1688.340 2494.510 1688.400 ;
        RECT 2484.530 1688.200 2494.510 1688.340 ;
        RECT 2484.530 1688.140 2484.850 1688.200 ;
        RECT 2494.190 1688.140 2494.510 1688.200 ;
        RECT 2494.190 18.600 2494.510 18.660 ;
        RECT 2595.390 18.600 2595.710 18.660 ;
        RECT 2494.190 18.460 2595.710 18.600 ;
        RECT 2494.190 18.400 2494.510 18.460 ;
        RECT 2595.390 18.400 2595.710 18.460 ;
      LAYER via ;
        RECT 2484.560 1688.140 2484.820 1688.400 ;
        RECT 2494.220 1688.140 2494.480 1688.400 ;
        RECT 2494.220 18.400 2494.480 18.660 ;
        RECT 2595.420 18.400 2595.680 18.660 ;
      LAYER met2 ;
        RECT 2484.480 1700.000 2484.760 1704.000 ;
        RECT 2484.620 1688.430 2484.760 1700.000 ;
        RECT 2484.560 1688.110 2484.820 1688.430 ;
        RECT 2494.220 1688.110 2494.480 1688.430 ;
        RECT 2494.280 18.690 2494.420 1688.110 ;
        RECT 2494.220 18.370 2494.480 18.690 ;
        RECT 2595.420 18.370 2595.680 18.690 ;
        RECT 2595.480 2.400 2595.620 18.370 ;
        RECT 2595.270 -4.800 2595.830 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2493.730 1684.600 2494.050 1684.660 ;
        RECT 2497.410 1684.600 2497.730 1684.660 ;
        RECT 2493.730 1684.460 2497.730 1684.600 ;
        RECT 2493.730 1684.400 2494.050 1684.460 ;
        RECT 2497.410 1684.400 2497.730 1684.460 ;
        RECT 2497.410 18.260 2497.730 18.320 ;
        RECT 2613.330 18.260 2613.650 18.320 ;
        RECT 2497.410 18.120 2613.650 18.260 ;
        RECT 2497.410 18.060 2497.730 18.120 ;
        RECT 2613.330 18.060 2613.650 18.120 ;
      LAYER via ;
        RECT 2493.760 1684.400 2494.020 1684.660 ;
        RECT 2497.440 1684.400 2497.700 1684.660 ;
        RECT 2497.440 18.060 2497.700 18.320 ;
        RECT 2613.360 18.060 2613.620 18.320 ;
      LAYER met2 ;
        RECT 2493.680 1700.000 2493.960 1704.000 ;
        RECT 2493.820 1684.690 2493.960 1700.000 ;
        RECT 2493.760 1684.370 2494.020 1684.690 ;
        RECT 2497.440 1684.370 2497.700 1684.690 ;
        RECT 2497.500 18.350 2497.640 1684.370 ;
        RECT 2497.440 18.030 2497.700 18.350 ;
        RECT 2613.360 18.030 2613.620 18.350 ;
        RECT 2613.420 2.400 2613.560 18.030 ;
        RECT 2613.210 -4.800 2613.770 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2503.850 17.580 2504.170 17.640 ;
        RECT 2631.270 17.580 2631.590 17.640 ;
        RECT 2503.850 17.440 2631.590 17.580 ;
        RECT 2503.850 17.380 2504.170 17.440 ;
        RECT 2631.270 17.380 2631.590 17.440 ;
      LAYER via ;
        RECT 2503.880 17.380 2504.140 17.640 ;
        RECT 2631.300 17.380 2631.560 17.640 ;
      LAYER met2 ;
        RECT 2502.880 1700.410 2503.160 1704.000 ;
        RECT 2502.880 1700.270 2504.080 1700.410 ;
        RECT 2502.880 1700.000 2503.160 1700.270 ;
        RECT 2503.940 17.670 2504.080 1700.270 ;
        RECT 2503.880 17.350 2504.140 17.670 ;
        RECT 2631.300 17.350 2631.560 17.670 ;
        RECT 2631.360 2.400 2631.500 17.350 ;
        RECT 2631.150 -4.800 2631.710 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2512.130 1688.000 2512.450 1688.060 ;
        RECT 2517.650 1688.000 2517.970 1688.060 ;
        RECT 2512.130 1687.860 2517.970 1688.000 ;
        RECT 2512.130 1687.800 2512.450 1687.860 ;
        RECT 2517.650 1687.800 2517.970 1687.860 ;
        RECT 2517.650 24.720 2517.970 24.780 ;
        RECT 2648.750 24.720 2649.070 24.780 ;
        RECT 2517.650 24.580 2649.070 24.720 ;
        RECT 2517.650 24.520 2517.970 24.580 ;
        RECT 2648.750 24.520 2649.070 24.580 ;
      LAYER via ;
        RECT 2512.160 1687.800 2512.420 1688.060 ;
        RECT 2517.680 1687.800 2517.940 1688.060 ;
        RECT 2517.680 24.520 2517.940 24.780 ;
        RECT 2648.780 24.520 2649.040 24.780 ;
      LAYER met2 ;
        RECT 2512.080 1700.000 2512.360 1704.000 ;
        RECT 2512.220 1688.090 2512.360 1700.000 ;
        RECT 2512.160 1687.770 2512.420 1688.090 ;
        RECT 2517.680 1687.770 2517.940 1688.090 ;
        RECT 2517.740 24.810 2517.880 1687.770 ;
        RECT 2517.680 24.490 2517.940 24.810 ;
        RECT 2648.780 24.490 2649.040 24.810 ;
        RECT 2648.840 16.730 2648.980 24.490 ;
        RECT 2648.840 16.590 2649.440 16.730 ;
        RECT 2649.300 2.400 2649.440 16.590 ;
        RECT 2649.090 -4.800 2649.650 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2521.330 1689.020 2521.650 1689.080 ;
        RECT 2525.010 1689.020 2525.330 1689.080 ;
        RECT 2521.330 1688.880 2525.330 1689.020 ;
        RECT 2521.330 1688.820 2521.650 1688.880 ;
        RECT 2525.010 1688.820 2525.330 1688.880 ;
        RECT 2525.010 14.860 2525.330 14.920 ;
        RECT 2667.150 14.860 2667.470 14.920 ;
        RECT 2525.010 14.720 2667.470 14.860 ;
        RECT 2525.010 14.660 2525.330 14.720 ;
        RECT 2667.150 14.660 2667.470 14.720 ;
      LAYER via ;
        RECT 2521.360 1688.820 2521.620 1689.080 ;
        RECT 2525.040 1688.820 2525.300 1689.080 ;
        RECT 2525.040 14.660 2525.300 14.920 ;
        RECT 2667.180 14.660 2667.440 14.920 ;
      LAYER met2 ;
        RECT 2521.280 1700.000 2521.560 1704.000 ;
        RECT 2521.420 1689.110 2521.560 1700.000 ;
        RECT 2521.360 1688.790 2521.620 1689.110 ;
        RECT 2525.040 1688.790 2525.300 1689.110 ;
        RECT 2525.100 14.950 2525.240 1688.790 ;
        RECT 2525.040 14.630 2525.300 14.950 ;
        RECT 2667.180 14.630 2667.440 14.950 ;
        RECT 2667.240 2.400 2667.380 14.630 ;
        RECT 2667.030 -4.800 2667.590 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2531.450 24.040 2531.770 24.100 ;
        RECT 2684.630 24.040 2684.950 24.100 ;
        RECT 2531.450 23.900 2684.950 24.040 ;
        RECT 2531.450 23.840 2531.770 23.900 ;
        RECT 2684.630 23.840 2684.950 23.900 ;
      LAYER via ;
        RECT 2531.480 23.840 2531.740 24.100 ;
        RECT 2684.660 23.840 2684.920 24.100 ;
      LAYER met2 ;
        RECT 2530.480 1700.410 2530.760 1704.000 ;
        RECT 2530.480 1700.270 2531.680 1700.410 ;
        RECT 2530.480 1700.000 2530.760 1700.270 ;
        RECT 2531.540 24.130 2531.680 1700.270 ;
        RECT 2531.480 23.810 2531.740 24.130 ;
        RECT 2684.660 23.810 2684.920 24.130 ;
        RECT 2684.720 2.400 2684.860 23.810 ;
        RECT 2684.510 -4.800 2685.070 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2539.730 1689.020 2540.050 1689.080 ;
        RECT 2545.710 1689.020 2546.030 1689.080 ;
        RECT 2539.730 1688.880 2546.030 1689.020 ;
        RECT 2539.730 1688.820 2540.050 1688.880 ;
        RECT 2545.710 1688.820 2546.030 1688.880 ;
        RECT 2545.710 24.380 2546.030 24.440 ;
        RECT 2702.570 24.380 2702.890 24.440 ;
        RECT 2545.710 24.240 2702.890 24.380 ;
        RECT 2545.710 24.180 2546.030 24.240 ;
        RECT 2702.570 24.180 2702.890 24.240 ;
      LAYER via ;
        RECT 2539.760 1688.820 2540.020 1689.080 ;
        RECT 2545.740 1688.820 2546.000 1689.080 ;
        RECT 2545.740 24.180 2546.000 24.440 ;
        RECT 2702.600 24.180 2702.860 24.440 ;
      LAYER met2 ;
        RECT 2539.680 1700.000 2539.960 1704.000 ;
        RECT 2539.820 1689.110 2539.960 1700.000 ;
        RECT 2539.760 1688.790 2540.020 1689.110 ;
        RECT 2545.740 1688.790 2546.000 1689.110 ;
        RECT 2545.800 24.470 2545.940 1688.790 ;
        RECT 2545.740 24.150 2546.000 24.470 ;
        RECT 2702.600 24.150 2702.860 24.470 ;
        RECT 2702.660 2.400 2702.800 24.150 ;
        RECT 2702.450 -4.800 2703.010 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2548.930 1685.280 2549.250 1685.340 ;
        RECT 2701.650 1685.280 2701.970 1685.340 ;
        RECT 2548.930 1685.140 2701.970 1685.280 ;
        RECT 2548.930 1685.080 2549.250 1685.140 ;
        RECT 2701.650 1685.080 2701.970 1685.140 ;
        RECT 2701.650 16.220 2701.970 16.280 ;
        RECT 2720.510 16.220 2720.830 16.280 ;
        RECT 2701.650 16.080 2720.830 16.220 ;
        RECT 2701.650 16.020 2701.970 16.080 ;
        RECT 2720.510 16.020 2720.830 16.080 ;
      LAYER via ;
        RECT 2548.960 1685.080 2549.220 1685.340 ;
        RECT 2701.680 1685.080 2701.940 1685.340 ;
        RECT 2701.680 16.020 2701.940 16.280 ;
        RECT 2720.540 16.020 2720.800 16.280 ;
      LAYER met2 ;
        RECT 2548.880 1700.000 2549.160 1704.000 ;
        RECT 2549.020 1685.370 2549.160 1700.000 ;
        RECT 2548.960 1685.050 2549.220 1685.370 ;
        RECT 2701.680 1685.050 2701.940 1685.370 ;
        RECT 2701.740 16.310 2701.880 1685.050 ;
        RECT 2701.680 15.990 2701.940 16.310 ;
        RECT 2720.540 15.990 2720.800 16.310 ;
        RECT 2720.600 2.400 2720.740 15.990 ;
        RECT 2720.390 -4.800 2720.950 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2559.510 15.880 2559.830 15.940 ;
        RECT 2559.510 15.740 2694.520 15.880 ;
        RECT 2559.510 15.680 2559.830 15.740 ;
        RECT 2694.380 15.540 2694.520 15.740 ;
        RECT 2738.450 15.540 2738.770 15.600 ;
        RECT 2694.380 15.400 2738.770 15.540 ;
        RECT 2738.450 15.340 2738.770 15.400 ;
      LAYER via ;
        RECT 2559.540 15.680 2559.800 15.940 ;
        RECT 2738.480 15.340 2738.740 15.600 ;
      LAYER met2 ;
        RECT 2558.080 1700.410 2558.360 1704.000 ;
        RECT 2558.080 1700.270 2559.740 1700.410 ;
        RECT 2558.080 1700.000 2558.360 1700.270 ;
        RECT 2559.600 15.970 2559.740 1700.270 ;
        RECT 2559.540 15.650 2559.800 15.970 ;
        RECT 2738.480 15.310 2738.740 15.630 ;
        RECT 2738.540 2.400 2738.680 15.310 ;
        RECT 2738.330 -4.800 2738.890 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2567.330 1684.260 2567.650 1684.320 ;
        RECT 2714.990 1684.260 2715.310 1684.320 ;
        RECT 2567.330 1684.120 2715.310 1684.260 ;
        RECT 2567.330 1684.060 2567.650 1684.120 ;
        RECT 2714.990 1684.060 2715.310 1684.120 ;
        RECT 2755.930 15.540 2756.250 15.600 ;
        RECT 2739.000 15.400 2756.250 15.540 ;
        RECT 2714.990 14.520 2715.310 14.580 ;
        RECT 2739.000 14.520 2739.140 15.400 ;
        RECT 2755.930 15.340 2756.250 15.400 ;
        RECT 2714.990 14.380 2739.140 14.520 ;
        RECT 2714.990 14.320 2715.310 14.380 ;
      LAYER via ;
        RECT 2567.360 1684.060 2567.620 1684.320 ;
        RECT 2715.020 1684.060 2715.280 1684.320 ;
        RECT 2715.020 14.320 2715.280 14.580 ;
        RECT 2755.960 15.340 2756.220 15.600 ;
      LAYER met2 ;
        RECT 2567.280 1700.000 2567.560 1704.000 ;
        RECT 2567.420 1684.350 2567.560 1700.000 ;
        RECT 2567.360 1684.030 2567.620 1684.350 ;
        RECT 2715.020 1684.030 2715.280 1684.350 ;
        RECT 2715.080 14.610 2715.220 1684.030 ;
        RECT 2755.960 15.310 2756.220 15.630 ;
        RECT 2715.020 14.290 2715.280 14.610 ;
        RECT 2756.020 2.400 2756.160 15.310 ;
        RECT 2755.810 -4.800 2756.370 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 834.510 60.420 834.830 60.480 ;
        RECT 1573.730 60.420 1574.050 60.480 ;
        RECT 834.510 60.280 1574.050 60.420 ;
        RECT 834.510 60.220 834.830 60.280 ;
        RECT 1573.730 60.220 1574.050 60.280 ;
      LAYER via ;
        RECT 834.540 60.220 834.800 60.480 ;
        RECT 1573.760 60.220 1574.020 60.480 ;
      LAYER met2 ;
        RECT 1575.520 1700.410 1575.800 1704.000 ;
        RECT 1573.820 1700.270 1575.800 1700.410 ;
        RECT 1573.820 60.510 1573.960 1700.270 ;
        RECT 1575.520 1700.000 1575.800 1700.270 ;
        RECT 834.540 60.190 834.800 60.510 ;
        RECT 1573.760 60.190 1574.020 60.510 ;
        RECT 834.600 16.730 834.740 60.190 ;
        RECT 829.540 16.590 834.740 16.730 ;
        RECT 829.540 2.400 829.680 16.590 ;
        RECT 829.330 -4.800 829.890 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2600.985 1684.785 2601.155 1686.995 ;
      LAYER mcon ;
        RECT 2600.985 1686.825 2601.155 1686.995 ;
      LAYER met1 ;
        RECT 2576.530 1687.320 2576.850 1687.380 ;
        RECT 2576.530 1687.180 2597.460 1687.320 ;
        RECT 2576.530 1687.120 2576.850 1687.180 ;
        RECT 2597.320 1686.980 2597.460 1687.180 ;
        RECT 2600.925 1686.980 2601.215 1687.025 ;
        RECT 2597.320 1686.840 2601.215 1686.980 ;
        RECT 2600.925 1686.795 2601.215 1686.840 ;
        RECT 2600.925 1684.940 2601.215 1684.985 ;
        RECT 2728.790 1684.940 2729.110 1685.000 ;
        RECT 2600.925 1684.800 2729.110 1684.940 ;
        RECT 2600.925 1684.755 2601.215 1684.800 ;
        RECT 2728.790 1684.740 2729.110 1684.800 ;
        RECT 2728.790 16.220 2729.110 16.280 ;
        RECT 2773.870 16.220 2774.190 16.280 ;
        RECT 2728.790 16.080 2774.190 16.220 ;
        RECT 2728.790 16.020 2729.110 16.080 ;
        RECT 2773.870 16.020 2774.190 16.080 ;
      LAYER via ;
        RECT 2576.560 1687.120 2576.820 1687.380 ;
        RECT 2728.820 1684.740 2729.080 1685.000 ;
        RECT 2728.820 16.020 2729.080 16.280 ;
        RECT 2773.900 16.020 2774.160 16.280 ;
      LAYER met2 ;
        RECT 2576.480 1700.000 2576.760 1704.000 ;
        RECT 2576.620 1687.410 2576.760 1700.000 ;
        RECT 2576.560 1687.090 2576.820 1687.410 ;
        RECT 2728.820 1684.710 2729.080 1685.030 ;
        RECT 2728.880 16.310 2729.020 1684.710 ;
        RECT 2728.820 15.990 2729.080 16.310 ;
        RECT 2773.900 15.990 2774.160 16.310 ;
        RECT 2773.960 2.400 2774.100 15.990 ;
        RECT 2773.750 -4.800 2774.310 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2749.490 1686.640 2749.810 1686.700 ;
        RECT 2603.760 1686.500 2749.810 1686.640 ;
        RECT 2585.730 1686.300 2586.050 1686.360 ;
        RECT 2603.760 1686.300 2603.900 1686.500 ;
        RECT 2749.490 1686.440 2749.810 1686.500 ;
        RECT 2585.730 1686.160 2603.900 1686.300 ;
        RECT 2585.730 1686.100 2586.050 1686.160 ;
        RECT 2791.810 16.560 2792.130 16.620 ;
        RECT 2774.420 16.420 2792.130 16.560 ;
        RECT 2749.490 15.880 2749.810 15.940 ;
        RECT 2774.420 15.880 2774.560 16.420 ;
        RECT 2791.810 16.360 2792.130 16.420 ;
        RECT 2749.490 15.740 2774.560 15.880 ;
        RECT 2749.490 15.680 2749.810 15.740 ;
      LAYER via ;
        RECT 2585.760 1686.100 2586.020 1686.360 ;
        RECT 2749.520 1686.440 2749.780 1686.700 ;
        RECT 2749.520 15.680 2749.780 15.940 ;
        RECT 2791.840 16.360 2792.100 16.620 ;
      LAYER met2 ;
        RECT 2585.680 1700.000 2585.960 1704.000 ;
        RECT 2585.820 1686.390 2585.960 1700.000 ;
        RECT 2749.520 1686.410 2749.780 1686.730 ;
        RECT 2585.760 1686.070 2586.020 1686.390 ;
        RECT 2749.580 15.970 2749.720 1686.410 ;
        RECT 2791.840 16.330 2792.100 16.650 ;
        RECT 2749.520 15.650 2749.780 15.970 ;
        RECT 2791.900 2.400 2792.040 16.330 ;
        RECT 2791.690 -4.800 2792.250 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2594.930 1684.940 2595.250 1685.000 ;
        RECT 2600.450 1684.940 2600.770 1685.000 ;
        RECT 2594.930 1684.800 2600.770 1684.940 ;
        RECT 2594.930 1684.740 2595.250 1684.800 ;
        RECT 2600.450 1684.740 2600.770 1684.800 ;
        RECT 2600.450 19.960 2600.770 20.020 ;
        RECT 2809.750 19.960 2810.070 20.020 ;
        RECT 2600.450 19.820 2810.070 19.960 ;
        RECT 2600.450 19.760 2600.770 19.820 ;
        RECT 2809.750 19.760 2810.070 19.820 ;
      LAYER via ;
        RECT 2594.960 1684.740 2595.220 1685.000 ;
        RECT 2600.480 1684.740 2600.740 1685.000 ;
        RECT 2600.480 19.760 2600.740 20.020 ;
        RECT 2809.780 19.760 2810.040 20.020 ;
      LAYER met2 ;
        RECT 2594.880 1700.000 2595.160 1704.000 ;
        RECT 2595.020 1685.030 2595.160 1700.000 ;
        RECT 2594.960 1684.710 2595.220 1685.030 ;
        RECT 2600.480 1684.710 2600.740 1685.030 ;
        RECT 2600.540 20.050 2600.680 1684.710 ;
        RECT 2600.480 19.730 2600.740 20.050 ;
        RECT 2809.780 19.730 2810.040 20.050 ;
        RECT 2809.840 2.400 2809.980 19.730 ;
        RECT 2809.630 -4.800 2810.190 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2604.130 1689.700 2604.450 1689.760 ;
        RECT 2783.990 1689.700 2784.310 1689.760 ;
        RECT 2604.130 1689.560 2784.310 1689.700 ;
        RECT 2604.130 1689.500 2604.450 1689.560 ;
        RECT 2783.990 1689.500 2784.310 1689.560 ;
        RECT 2783.990 16.900 2784.310 16.960 ;
        RECT 2827.690 16.900 2828.010 16.960 ;
        RECT 2783.990 16.760 2828.010 16.900 ;
        RECT 2783.990 16.700 2784.310 16.760 ;
        RECT 2827.690 16.700 2828.010 16.760 ;
      LAYER via ;
        RECT 2604.160 1689.500 2604.420 1689.760 ;
        RECT 2784.020 1689.500 2784.280 1689.760 ;
        RECT 2784.020 16.700 2784.280 16.960 ;
        RECT 2827.720 16.700 2827.980 16.960 ;
      LAYER met2 ;
        RECT 2604.080 1700.000 2604.360 1704.000 ;
        RECT 2604.220 1689.790 2604.360 1700.000 ;
        RECT 2604.160 1689.470 2604.420 1689.790 ;
        RECT 2784.020 1689.470 2784.280 1689.790 ;
        RECT 2784.080 16.990 2784.220 1689.470 ;
        RECT 2784.020 16.670 2784.280 16.990 ;
        RECT 2827.720 16.670 2827.980 16.990 ;
        RECT 2827.780 2.400 2827.920 16.670 ;
        RECT 2827.570 -4.800 2828.130 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2614.710 18.600 2615.030 18.660 ;
        RECT 2845.170 18.600 2845.490 18.660 ;
        RECT 2614.710 18.460 2845.490 18.600 ;
        RECT 2614.710 18.400 2615.030 18.460 ;
        RECT 2845.170 18.400 2845.490 18.460 ;
      LAYER via ;
        RECT 2614.740 18.400 2615.000 18.660 ;
        RECT 2845.200 18.400 2845.460 18.660 ;
      LAYER met2 ;
        RECT 2613.280 1700.410 2613.560 1704.000 ;
        RECT 2613.280 1700.270 2614.940 1700.410 ;
        RECT 2613.280 1700.000 2613.560 1700.270 ;
        RECT 2614.800 18.690 2614.940 1700.270 ;
        RECT 2614.740 18.370 2615.000 18.690 ;
        RECT 2845.200 18.370 2845.460 18.690 ;
        RECT 2845.260 2.400 2845.400 18.370 ;
        RECT 2845.050 -4.800 2845.610 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2622.530 1683.920 2622.850 1683.980 ;
        RECT 2628.050 1683.920 2628.370 1683.980 ;
        RECT 2622.530 1683.780 2628.370 1683.920 ;
        RECT 2622.530 1683.720 2622.850 1683.780 ;
        RECT 2628.050 1683.720 2628.370 1683.780 ;
        RECT 2628.050 18.940 2628.370 19.000 ;
        RECT 2863.110 18.940 2863.430 19.000 ;
        RECT 2628.050 18.800 2863.430 18.940 ;
        RECT 2628.050 18.740 2628.370 18.800 ;
        RECT 2863.110 18.740 2863.430 18.800 ;
      LAYER via ;
        RECT 2622.560 1683.720 2622.820 1683.980 ;
        RECT 2628.080 1683.720 2628.340 1683.980 ;
        RECT 2628.080 18.740 2628.340 19.000 ;
        RECT 2863.140 18.740 2863.400 19.000 ;
      LAYER met2 ;
        RECT 2622.480 1700.000 2622.760 1704.000 ;
        RECT 2622.620 1684.010 2622.760 1700.000 ;
        RECT 2622.560 1683.690 2622.820 1684.010 ;
        RECT 2628.080 1683.690 2628.340 1684.010 ;
        RECT 2628.140 19.030 2628.280 1683.690 ;
        RECT 2628.080 18.710 2628.340 19.030 ;
        RECT 2863.140 18.710 2863.400 19.030 ;
        RECT 2863.200 2.400 2863.340 18.710 ;
        RECT 2862.990 -4.800 2863.550 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2657.565 1683.765 2657.735 1686.315 ;
      LAYER mcon ;
        RECT 2657.565 1686.145 2657.735 1686.315 ;
      LAYER met1 ;
        RECT 2657.505 1686.300 2657.795 1686.345 ;
        RECT 2790.890 1686.300 2791.210 1686.360 ;
        RECT 2657.505 1686.160 2791.210 1686.300 ;
        RECT 2657.505 1686.115 2657.795 1686.160 ;
        RECT 2790.890 1686.100 2791.210 1686.160 ;
        RECT 2631.730 1683.920 2632.050 1683.980 ;
        RECT 2657.505 1683.920 2657.795 1683.965 ;
        RECT 2631.730 1683.780 2637.480 1683.920 ;
        RECT 2631.730 1683.720 2632.050 1683.780 ;
        RECT 2637.340 1683.580 2637.480 1683.780 ;
        RECT 2649.760 1683.780 2657.795 1683.920 ;
        RECT 2649.760 1683.580 2649.900 1683.780 ;
        RECT 2657.505 1683.735 2657.795 1683.780 ;
        RECT 2637.340 1683.440 2649.900 1683.580 ;
        RECT 2790.890 20.640 2791.210 20.700 ;
        RECT 2881.050 20.640 2881.370 20.700 ;
        RECT 2790.890 20.500 2881.370 20.640 ;
        RECT 2790.890 20.440 2791.210 20.500 ;
        RECT 2881.050 20.440 2881.370 20.500 ;
      LAYER via ;
        RECT 2790.920 1686.100 2791.180 1686.360 ;
        RECT 2631.760 1683.720 2632.020 1683.980 ;
        RECT 2790.920 20.440 2791.180 20.700 ;
        RECT 2881.080 20.440 2881.340 20.700 ;
      LAYER met2 ;
        RECT 2631.680 1700.000 2631.960 1704.000 ;
        RECT 2631.820 1684.010 2631.960 1700.000 ;
        RECT 2790.920 1686.070 2791.180 1686.390 ;
        RECT 2631.760 1683.690 2632.020 1684.010 ;
        RECT 2790.980 20.730 2791.120 1686.070 ;
        RECT 2790.920 20.410 2791.180 20.730 ;
        RECT 2881.080 20.410 2881.340 20.730 ;
        RECT 2881.140 2.400 2881.280 20.410 ;
        RECT 2880.930 -4.800 2881.490 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2825.390 19.620 2825.710 19.680 ;
        RECT 2898.990 19.620 2899.310 19.680 ;
        RECT 2825.390 19.480 2899.310 19.620 ;
        RECT 2825.390 19.420 2825.710 19.480 ;
        RECT 2898.990 19.420 2899.310 19.480 ;
      LAYER via ;
        RECT 2825.420 19.420 2825.680 19.680 ;
        RECT 2899.020 19.420 2899.280 19.680 ;
      LAYER met2 ;
        RECT 2640.880 1700.000 2641.160 1704.000 ;
        RECT 2641.020 1686.925 2641.160 1700.000 ;
        RECT 2640.950 1686.555 2641.230 1686.925 ;
        RECT 2825.410 1686.555 2825.690 1686.925 ;
        RECT 2825.480 19.710 2825.620 1686.555 ;
        RECT 2825.420 19.390 2825.680 19.710 ;
        RECT 2899.020 19.390 2899.280 19.710 ;
        RECT 2899.080 2.400 2899.220 19.390 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
      LAYER via2 ;
        RECT 2640.950 1686.600 2641.230 1686.880 ;
        RECT 2825.410 1686.600 2825.690 1686.880 ;
      LAYER met3 ;
        RECT 2640.925 1686.890 2641.255 1686.905 ;
        RECT 2825.385 1686.890 2825.715 1686.905 ;
        RECT 2640.925 1686.590 2825.715 1686.890 ;
        RECT 2640.925 1686.575 2641.255 1686.590 ;
        RECT 2825.385 1686.575 2825.715 1686.590 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1580.170 1689.700 1580.490 1689.760 ;
        RECT 1583.390 1689.700 1583.710 1689.760 ;
        RECT 1580.170 1689.560 1583.710 1689.700 ;
        RECT 1580.170 1689.500 1580.490 1689.560 ;
        RECT 1583.390 1689.500 1583.710 1689.560 ;
        RECT 848.310 60.760 848.630 60.820 ;
        RECT 1580.170 60.760 1580.490 60.820 ;
        RECT 848.310 60.620 1580.490 60.760 ;
        RECT 848.310 60.560 848.630 60.620 ;
        RECT 1580.170 60.560 1580.490 60.620 ;
      LAYER via ;
        RECT 1580.200 1689.500 1580.460 1689.760 ;
        RECT 1583.420 1689.500 1583.680 1689.760 ;
        RECT 848.340 60.560 848.600 60.820 ;
        RECT 1580.200 60.560 1580.460 60.820 ;
      LAYER met2 ;
        RECT 1584.720 1700.410 1585.000 1704.000 ;
        RECT 1583.480 1700.270 1585.000 1700.410 ;
        RECT 1583.480 1689.790 1583.620 1700.270 ;
        RECT 1584.720 1700.000 1585.000 1700.270 ;
        RECT 1580.200 1689.470 1580.460 1689.790 ;
        RECT 1583.420 1689.470 1583.680 1689.790 ;
        RECT 1580.260 60.850 1580.400 1689.470 ;
        RECT 848.340 60.530 848.600 60.850 ;
        RECT 1580.200 60.530 1580.460 60.850 ;
        RECT 848.400 16.730 848.540 60.530 ;
        RECT 847.020 16.590 848.540 16.730 ;
        RECT 847.020 2.400 847.160 16.590 ;
        RECT 846.810 -4.800 847.370 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1587.990 1689.700 1588.310 1689.760 ;
        RECT 1591.670 1689.700 1591.990 1689.760 ;
        RECT 1587.990 1689.560 1591.990 1689.700 ;
        RECT 1587.990 1689.500 1588.310 1689.560 ;
        RECT 1591.670 1689.500 1591.990 1689.560 ;
        RECT 869.010 61.100 869.330 61.160 ;
        RECT 1587.990 61.100 1588.310 61.160 ;
        RECT 869.010 60.960 1588.310 61.100 ;
        RECT 869.010 60.900 869.330 60.960 ;
        RECT 1587.990 60.900 1588.310 60.960 ;
        RECT 864.870 2.960 865.190 3.020 ;
        RECT 869.010 2.960 869.330 3.020 ;
        RECT 864.870 2.820 869.330 2.960 ;
        RECT 864.870 2.760 865.190 2.820 ;
        RECT 869.010 2.760 869.330 2.820 ;
      LAYER via ;
        RECT 1588.020 1689.500 1588.280 1689.760 ;
        RECT 1591.700 1689.500 1591.960 1689.760 ;
        RECT 869.040 60.900 869.300 61.160 ;
        RECT 1588.020 60.900 1588.280 61.160 ;
        RECT 864.900 2.760 865.160 3.020 ;
        RECT 869.040 2.760 869.300 3.020 ;
      LAYER met2 ;
        RECT 1593.460 1700.410 1593.740 1704.000 ;
        RECT 1591.760 1700.270 1593.740 1700.410 ;
        RECT 1591.760 1689.790 1591.900 1700.270 ;
        RECT 1593.460 1700.000 1593.740 1700.270 ;
        RECT 1588.020 1689.470 1588.280 1689.790 ;
        RECT 1591.700 1689.470 1591.960 1689.790 ;
        RECT 1588.080 61.190 1588.220 1689.470 ;
        RECT 869.040 60.870 869.300 61.190 ;
        RECT 1588.020 60.870 1588.280 61.190 ;
        RECT 869.100 3.050 869.240 60.870 ;
        RECT 864.900 2.730 865.160 3.050 ;
        RECT 869.040 2.730 869.300 3.050 ;
        RECT 864.960 2.400 865.100 2.730 ;
        RECT 864.750 -4.800 865.310 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 882.810 61.440 883.130 61.500 ;
        RECT 1601.330 61.440 1601.650 61.500 ;
        RECT 882.810 61.300 1601.650 61.440 ;
        RECT 882.810 61.240 883.130 61.300 ;
        RECT 1601.330 61.240 1601.650 61.300 ;
      LAYER via ;
        RECT 882.840 61.240 883.100 61.500 ;
        RECT 1601.360 61.240 1601.620 61.500 ;
      LAYER met2 ;
        RECT 1602.660 1700.410 1602.940 1704.000 ;
        RECT 1601.420 1700.270 1602.940 1700.410 ;
        RECT 1601.420 61.530 1601.560 1700.270 ;
        RECT 1602.660 1700.000 1602.940 1700.270 ;
        RECT 882.840 61.210 883.100 61.530 ;
        RECT 1601.360 61.210 1601.620 61.530 ;
        RECT 882.900 2.400 883.040 61.210 ;
        RECT 882.690 -4.800 883.250 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1608.765 1360.765 1608.935 1400.715 ;
        RECT 1608.765 1256.045 1608.935 1304.155 ;
        RECT 1608.305 917.745 1608.475 932.195 ;
        RECT 1608.305 676.005 1608.475 717.655 ;
        RECT 1608.765 572.645 1608.935 594.235 ;
        RECT 1608.765 235.025 1608.935 255.935 ;
      LAYER mcon ;
        RECT 1608.765 1400.545 1608.935 1400.715 ;
        RECT 1608.765 1303.985 1608.935 1304.155 ;
        RECT 1608.305 932.025 1608.475 932.195 ;
        RECT 1608.305 717.485 1608.475 717.655 ;
        RECT 1608.765 594.065 1608.935 594.235 ;
        RECT 1608.765 255.765 1608.935 255.935 ;
      LAYER met1 ;
        RECT 1608.230 1628.500 1608.550 1628.560 ;
        RECT 1610.530 1628.500 1610.850 1628.560 ;
        RECT 1608.230 1628.360 1610.850 1628.500 ;
        RECT 1608.230 1628.300 1608.550 1628.360 ;
        RECT 1610.530 1628.300 1610.850 1628.360 ;
        RECT 1607.310 1580.220 1607.630 1580.280 ;
        RECT 1608.690 1580.220 1609.010 1580.280 ;
        RECT 1607.310 1580.080 1609.010 1580.220 ;
        RECT 1607.310 1580.020 1607.630 1580.080 ;
        RECT 1608.690 1580.020 1609.010 1580.080 ;
        RECT 1607.310 1556.080 1607.630 1556.140 ;
        RECT 1608.690 1556.080 1609.010 1556.140 ;
        RECT 1607.310 1555.940 1609.010 1556.080 ;
        RECT 1607.310 1555.880 1607.630 1555.940 ;
        RECT 1608.690 1555.880 1609.010 1555.940 ;
        RECT 1608.690 1463.060 1609.010 1463.320 ;
        RECT 1608.780 1462.640 1608.920 1463.060 ;
        RECT 1608.690 1462.380 1609.010 1462.640 ;
        RECT 1608.690 1400.700 1609.010 1400.760 ;
        RECT 1608.495 1400.560 1609.010 1400.700 ;
        RECT 1608.690 1400.500 1609.010 1400.560 ;
        RECT 1608.690 1360.920 1609.010 1360.980 ;
        RECT 1608.495 1360.780 1609.010 1360.920 ;
        RECT 1608.690 1360.720 1609.010 1360.780 ;
        RECT 1608.690 1304.140 1609.010 1304.200 ;
        RECT 1608.495 1304.000 1609.010 1304.140 ;
        RECT 1608.690 1303.940 1609.010 1304.000 ;
        RECT 1608.690 1256.200 1609.010 1256.260 ;
        RECT 1608.495 1256.060 1609.010 1256.200 ;
        RECT 1608.690 1256.000 1609.010 1256.060 ;
        RECT 1609.150 1173.240 1609.470 1173.300 ;
        RECT 1608.780 1173.100 1609.470 1173.240 ;
        RECT 1608.780 1172.960 1608.920 1173.100 ;
        RECT 1609.150 1173.040 1609.470 1173.100 ;
        RECT 1608.690 1172.700 1609.010 1172.960 ;
        RECT 1608.690 1080.080 1609.010 1080.140 ;
        RECT 1609.610 1080.080 1609.930 1080.140 ;
        RECT 1608.690 1079.940 1609.930 1080.080 ;
        RECT 1608.690 1079.880 1609.010 1079.940 ;
        RECT 1609.610 1079.880 1609.930 1079.940 ;
        RECT 1608.690 1007.320 1609.010 1007.380 ;
        RECT 1609.610 1007.320 1609.930 1007.380 ;
        RECT 1608.690 1007.180 1609.930 1007.320 ;
        RECT 1608.690 1007.120 1609.010 1007.180 ;
        RECT 1609.610 1007.120 1609.930 1007.180 ;
        RECT 1608.245 932.180 1608.535 932.225 ;
        RECT 1608.690 932.180 1609.010 932.240 ;
        RECT 1608.245 932.040 1609.010 932.180 ;
        RECT 1608.245 931.995 1608.535 932.040 ;
        RECT 1608.690 931.980 1609.010 932.040 ;
        RECT 1608.230 917.900 1608.550 917.960 ;
        RECT 1608.035 917.760 1608.550 917.900 ;
        RECT 1608.230 917.700 1608.550 917.760 ;
        RECT 1608.230 869.620 1608.550 869.680 ;
        RECT 1608.690 869.620 1609.010 869.680 ;
        RECT 1608.230 869.480 1609.010 869.620 ;
        RECT 1608.230 869.420 1608.550 869.480 ;
        RECT 1608.690 869.420 1609.010 869.480 ;
        RECT 1607.310 843.100 1607.630 843.160 ;
        RECT 1608.690 843.100 1609.010 843.160 ;
        RECT 1607.310 842.960 1609.010 843.100 ;
        RECT 1607.310 842.900 1607.630 842.960 ;
        RECT 1608.690 842.900 1609.010 842.960 ;
        RECT 1607.310 796.860 1607.630 796.920 ;
        RECT 1608.690 796.860 1609.010 796.920 ;
        RECT 1607.310 796.720 1609.010 796.860 ;
        RECT 1607.310 796.660 1607.630 796.720 ;
        RECT 1608.690 796.660 1609.010 796.720 ;
        RECT 1608.230 717.640 1608.550 717.700 ;
        RECT 1608.035 717.500 1608.550 717.640 ;
        RECT 1608.230 717.440 1608.550 717.500 ;
        RECT 1608.230 676.160 1608.550 676.220 ;
        RECT 1608.035 676.020 1608.550 676.160 ;
        RECT 1608.230 675.960 1608.550 676.020 ;
        RECT 1608.690 594.220 1609.010 594.280 ;
        RECT 1608.495 594.080 1609.010 594.220 ;
        RECT 1608.690 594.020 1609.010 594.080 ;
        RECT 1608.690 572.800 1609.010 572.860 ;
        RECT 1608.495 572.660 1609.010 572.800 ;
        RECT 1608.690 572.600 1609.010 572.660 ;
        RECT 1608.690 255.920 1609.010 255.980 ;
        RECT 1608.495 255.780 1609.010 255.920 ;
        RECT 1608.690 255.720 1609.010 255.780 ;
        RECT 1608.690 235.180 1609.010 235.240 ;
        RECT 1608.495 235.040 1609.010 235.180 ;
        RECT 1608.690 234.980 1609.010 235.040 ;
        RECT 1608.230 234.500 1608.550 234.560 ;
        RECT 1608.690 234.500 1609.010 234.560 ;
        RECT 1608.230 234.360 1609.010 234.500 ;
        RECT 1608.230 234.300 1608.550 234.360 ;
        RECT 1608.690 234.300 1609.010 234.360 ;
        RECT 1608.230 145.080 1608.550 145.140 ;
        RECT 1608.690 145.080 1609.010 145.140 ;
        RECT 1608.230 144.940 1609.010 145.080 ;
        RECT 1608.230 144.880 1608.550 144.940 ;
        RECT 1608.690 144.880 1609.010 144.940 ;
        RECT 903.510 61.780 903.830 61.840 ;
        RECT 1608.690 61.780 1609.010 61.840 ;
        RECT 903.510 61.640 1609.010 61.780 ;
        RECT 903.510 61.580 903.830 61.640 ;
        RECT 1608.690 61.580 1609.010 61.640 ;
        RECT 900.750 2.960 901.070 3.020 ;
        RECT 903.510 2.960 903.830 3.020 ;
        RECT 900.750 2.820 903.830 2.960 ;
        RECT 900.750 2.760 901.070 2.820 ;
        RECT 903.510 2.760 903.830 2.820 ;
      LAYER via ;
        RECT 1608.260 1628.300 1608.520 1628.560 ;
        RECT 1610.560 1628.300 1610.820 1628.560 ;
        RECT 1607.340 1580.020 1607.600 1580.280 ;
        RECT 1608.720 1580.020 1608.980 1580.280 ;
        RECT 1607.340 1555.880 1607.600 1556.140 ;
        RECT 1608.720 1555.880 1608.980 1556.140 ;
        RECT 1608.720 1463.060 1608.980 1463.320 ;
        RECT 1608.720 1462.380 1608.980 1462.640 ;
        RECT 1608.720 1400.500 1608.980 1400.760 ;
        RECT 1608.720 1360.720 1608.980 1360.980 ;
        RECT 1608.720 1303.940 1608.980 1304.200 ;
        RECT 1608.720 1256.000 1608.980 1256.260 ;
        RECT 1609.180 1173.040 1609.440 1173.300 ;
        RECT 1608.720 1172.700 1608.980 1172.960 ;
        RECT 1608.720 1079.880 1608.980 1080.140 ;
        RECT 1609.640 1079.880 1609.900 1080.140 ;
        RECT 1608.720 1007.120 1608.980 1007.380 ;
        RECT 1609.640 1007.120 1609.900 1007.380 ;
        RECT 1608.720 931.980 1608.980 932.240 ;
        RECT 1608.260 917.700 1608.520 917.960 ;
        RECT 1608.260 869.420 1608.520 869.680 ;
        RECT 1608.720 869.420 1608.980 869.680 ;
        RECT 1607.340 842.900 1607.600 843.160 ;
        RECT 1608.720 842.900 1608.980 843.160 ;
        RECT 1607.340 796.660 1607.600 796.920 ;
        RECT 1608.720 796.660 1608.980 796.920 ;
        RECT 1608.260 717.440 1608.520 717.700 ;
        RECT 1608.260 675.960 1608.520 676.220 ;
        RECT 1608.720 594.020 1608.980 594.280 ;
        RECT 1608.720 572.600 1608.980 572.860 ;
        RECT 1608.720 255.720 1608.980 255.980 ;
        RECT 1608.720 234.980 1608.980 235.240 ;
        RECT 1608.260 234.300 1608.520 234.560 ;
        RECT 1608.720 234.300 1608.980 234.560 ;
        RECT 1608.260 144.880 1608.520 145.140 ;
        RECT 1608.720 144.880 1608.980 145.140 ;
        RECT 903.540 61.580 903.800 61.840 ;
        RECT 1608.720 61.580 1608.980 61.840 ;
        RECT 900.780 2.760 901.040 3.020 ;
        RECT 903.540 2.760 903.800 3.020 ;
      LAYER met2 ;
        RECT 1611.860 1700.410 1612.140 1704.000 ;
        RECT 1609.700 1700.270 1612.140 1700.410 ;
        RECT 1609.700 1676.725 1609.840 1700.270 ;
        RECT 1611.860 1700.000 1612.140 1700.270 ;
        RECT 1609.630 1676.355 1609.910 1676.725 ;
        RECT 1610.550 1676.355 1610.830 1676.725 ;
        RECT 1610.620 1628.590 1610.760 1676.355 ;
        RECT 1608.260 1628.445 1608.520 1628.590 ;
        RECT 1607.330 1628.075 1607.610 1628.445 ;
        RECT 1608.250 1628.075 1608.530 1628.445 ;
        RECT 1610.560 1628.270 1610.820 1628.590 ;
        RECT 1607.400 1580.310 1607.540 1628.075 ;
        RECT 1608.780 1580.310 1608.920 1580.465 ;
        RECT 1607.340 1580.165 1607.600 1580.310 ;
        RECT 1607.330 1579.795 1607.610 1580.165 ;
        RECT 1608.250 1580.050 1608.530 1580.165 ;
        RECT 1608.720 1580.050 1608.980 1580.310 ;
        RECT 1608.250 1579.990 1608.980 1580.050 ;
        RECT 1608.250 1579.910 1608.920 1579.990 ;
        RECT 1608.250 1579.795 1608.530 1579.910 ;
        RECT 1607.400 1556.170 1607.540 1579.795 ;
        RECT 1607.340 1555.850 1607.600 1556.170 ;
        RECT 1608.720 1555.850 1608.980 1556.170 ;
        RECT 1608.780 1463.350 1608.920 1555.850 ;
        RECT 1608.720 1463.030 1608.980 1463.350 ;
        RECT 1608.720 1462.350 1608.980 1462.670 ;
        RECT 1608.780 1400.790 1608.920 1462.350 ;
        RECT 1608.720 1400.470 1608.980 1400.790 ;
        RECT 1608.720 1360.690 1608.980 1361.010 ;
        RECT 1608.780 1304.230 1608.920 1360.690 ;
        RECT 1608.720 1303.910 1608.980 1304.230 ;
        RECT 1608.720 1255.970 1608.980 1256.290 ;
        RECT 1608.780 1207.410 1608.920 1255.970 ;
        RECT 1608.780 1207.270 1609.380 1207.410 ;
        RECT 1609.240 1173.330 1609.380 1207.270 ;
        RECT 1609.180 1173.010 1609.440 1173.330 ;
        RECT 1608.720 1172.670 1608.980 1172.990 ;
        RECT 1608.780 1080.170 1608.920 1172.670 ;
        RECT 1608.720 1079.850 1608.980 1080.170 ;
        RECT 1609.640 1079.850 1609.900 1080.170 ;
        RECT 1609.700 1055.885 1609.840 1079.850 ;
        RECT 1608.710 1055.515 1608.990 1055.885 ;
        RECT 1609.630 1055.515 1609.910 1055.885 ;
        RECT 1608.780 1007.410 1608.920 1055.515 ;
        RECT 1608.720 1007.090 1608.980 1007.410 ;
        RECT 1609.640 1007.090 1609.900 1007.410 ;
        RECT 1609.700 959.325 1609.840 1007.090 ;
        RECT 1608.710 958.955 1608.990 959.325 ;
        RECT 1609.630 958.955 1609.910 959.325 ;
        RECT 1608.780 932.270 1608.920 958.955 ;
        RECT 1608.720 931.950 1608.980 932.270 ;
        RECT 1608.260 917.670 1608.520 917.990 ;
        RECT 1608.320 869.710 1608.460 917.670 ;
        RECT 1608.260 869.390 1608.520 869.710 ;
        RECT 1608.720 869.390 1608.980 869.710 ;
        RECT 1608.780 843.190 1608.920 869.390 ;
        RECT 1607.340 842.870 1607.600 843.190 ;
        RECT 1608.720 842.870 1608.980 843.190 ;
        RECT 1607.400 796.950 1607.540 842.870 ;
        RECT 1607.340 796.630 1607.600 796.950 ;
        RECT 1608.720 796.630 1608.980 796.950 ;
        RECT 1608.780 748.410 1608.920 796.630 ;
        RECT 1608.320 748.270 1608.920 748.410 ;
        RECT 1608.320 717.730 1608.460 748.270 ;
        RECT 1608.260 717.410 1608.520 717.730 ;
        RECT 1608.260 675.930 1608.520 676.250 ;
        RECT 1608.320 650.490 1608.460 675.930 ;
        RECT 1608.320 650.350 1608.920 650.490 ;
        RECT 1608.780 594.310 1608.920 650.350 ;
        RECT 1608.720 593.990 1608.980 594.310 ;
        RECT 1608.720 572.570 1608.980 572.890 ;
        RECT 1608.780 256.010 1608.920 572.570 ;
        RECT 1608.720 255.690 1608.980 256.010 ;
        RECT 1608.720 234.950 1608.980 235.270 ;
        RECT 1608.780 234.590 1608.920 234.950 ;
        RECT 1608.260 234.270 1608.520 234.590 ;
        RECT 1608.720 234.270 1608.980 234.590 ;
        RECT 1608.320 145.170 1608.460 234.270 ;
        RECT 1608.260 144.850 1608.520 145.170 ;
        RECT 1608.720 144.850 1608.980 145.170 ;
        RECT 1608.780 61.870 1608.920 144.850 ;
        RECT 903.540 61.550 903.800 61.870 ;
        RECT 1608.720 61.550 1608.980 61.870 ;
        RECT 903.600 3.050 903.740 61.550 ;
        RECT 900.780 2.730 901.040 3.050 ;
        RECT 903.540 2.730 903.800 3.050 ;
        RECT 900.840 2.400 900.980 2.730 ;
        RECT 900.630 -4.800 901.190 2.400 ;
      LAYER via2 ;
        RECT 1609.630 1676.400 1609.910 1676.680 ;
        RECT 1610.550 1676.400 1610.830 1676.680 ;
        RECT 1607.330 1628.120 1607.610 1628.400 ;
        RECT 1608.250 1628.120 1608.530 1628.400 ;
        RECT 1607.330 1579.840 1607.610 1580.120 ;
        RECT 1608.250 1579.840 1608.530 1580.120 ;
        RECT 1608.710 1055.560 1608.990 1055.840 ;
        RECT 1609.630 1055.560 1609.910 1055.840 ;
        RECT 1608.710 959.000 1608.990 959.280 ;
        RECT 1609.630 959.000 1609.910 959.280 ;
      LAYER met3 ;
        RECT 1609.605 1676.690 1609.935 1676.705 ;
        RECT 1610.525 1676.690 1610.855 1676.705 ;
        RECT 1609.605 1676.390 1610.855 1676.690 ;
        RECT 1609.605 1676.375 1609.935 1676.390 ;
        RECT 1610.525 1676.375 1610.855 1676.390 ;
        RECT 1607.305 1628.410 1607.635 1628.425 ;
        RECT 1608.225 1628.410 1608.555 1628.425 ;
        RECT 1607.305 1628.110 1608.555 1628.410 ;
        RECT 1607.305 1628.095 1607.635 1628.110 ;
        RECT 1608.225 1628.095 1608.555 1628.110 ;
        RECT 1607.305 1580.130 1607.635 1580.145 ;
        RECT 1608.225 1580.130 1608.555 1580.145 ;
        RECT 1607.305 1579.830 1608.555 1580.130 ;
        RECT 1607.305 1579.815 1607.635 1579.830 ;
        RECT 1608.225 1579.815 1608.555 1579.830 ;
        RECT 1608.685 1055.850 1609.015 1055.865 ;
        RECT 1609.605 1055.850 1609.935 1055.865 ;
        RECT 1608.685 1055.550 1609.935 1055.850 ;
        RECT 1608.685 1055.535 1609.015 1055.550 ;
        RECT 1609.605 1055.535 1609.935 1055.550 ;
        RECT 1608.685 959.290 1609.015 959.305 ;
        RECT 1609.605 959.290 1609.935 959.305 ;
        RECT 1608.685 958.990 1609.935 959.290 ;
        RECT 1608.685 958.975 1609.015 958.990 ;
        RECT 1609.605 958.975 1609.935 958.990 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1615.590 1678.140 1615.910 1678.200 ;
        RECT 1619.270 1678.140 1619.590 1678.200 ;
        RECT 1615.590 1678.000 1619.590 1678.140 ;
        RECT 1615.590 1677.940 1615.910 1678.000 ;
        RECT 1619.270 1677.940 1619.590 1678.000 ;
        RECT 924.210 62.120 924.530 62.180 ;
        RECT 1615.590 62.120 1615.910 62.180 ;
        RECT 924.210 61.980 1615.910 62.120 ;
        RECT 924.210 61.920 924.530 61.980 ;
        RECT 1615.590 61.920 1615.910 61.980 ;
      LAYER via ;
        RECT 1615.620 1677.940 1615.880 1678.200 ;
        RECT 1619.300 1677.940 1619.560 1678.200 ;
        RECT 924.240 61.920 924.500 62.180 ;
        RECT 1615.620 61.920 1615.880 62.180 ;
      LAYER met2 ;
        RECT 1621.060 1700.410 1621.340 1704.000 ;
        RECT 1619.360 1700.270 1621.340 1700.410 ;
        RECT 1619.360 1678.230 1619.500 1700.270 ;
        RECT 1621.060 1700.000 1621.340 1700.270 ;
        RECT 1615.620 1677.910 1615.880 1678.230 ;
        RECT 1619.300 1677.910 1619.560 1678.230 ;
        RECT 1615.680 62.210 1615.820 1677.910 ;
        RECT 924.240 61.890 924.500 62.210 ;
        RECT 1615.620 61.890 1615.880 62.210 ;
        RECT 924.300 29.650 924.440 61.890 ;
        RECT 918.780 29.510 924.440 29.650 ;
        RECT 918.780 2.400 918.920 29.510 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 938.010 58.380 938.330 58.440 ;
        RECT 1628.930 58.380 1629.250 58.440 ;
        RECT 938.010 58.240 1629.250 58.380 ;
        RECT 938.010 58.180 938.330 58.240 ;
        RECT 1628.930 58.180 1629.250 58.240 ;
      LAYER via ;
        RECT 938.040 58.180 938.300 58.440 ;
        RECT 1628.960 58.180 1629.220 58.440 ;
      LAYER met2 ;
        RECT 1630.260 1700.410 1630.540 1704.000 ;
        RECT 1629.020 1700.270 1630.540 1700.410 ;
        RECT 1629.020 58.470 1629.160 1700.270 ;
        RECT 1630.260 1700.000 1630.540 1700.270 ;
        RECT 938.040 58.150 938.300 58.470 ;
        RECT 1628.960 58.150 1629.220 58.470 ;
        RECT 938.100 17.410 938.240 58.150 ;
        RECT 936.260 17.270 938.240 17.410 ;
        RECT 936.260 2.400 936.400 17.270 ;
        RECT 936.050 -4.800 936.610 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1636.365 1360.765 1636.535 1400.715 ;
        RECT 1636.365 1256.045 1636.535 1304.155 ;
        RECT 1636.365 565.845 1636.535 613.955 ;
      LAYER mcon ;
        RECT 1636.365 1400.545 1636.535 1400.715 ;
        RECT 1636.365 1303.985 1636.535 1304.155 ;
        RECT 1636.365 613.785 1636.535 613.955 ;
      LAYER met1 ;
        RECT 1636.290 1659.440 1636.610 1659.500 ;
        RECT 1637.210 1659.440 1637.530 1659.500 ;
        RECT 1636.290 1659.300 1637.530 1659.440 ;
        RECT 1636.290 1659.240 1636.610 1659.300 ;
        RECT 1637.210 1659.240 1637.530 1659.300 ;
        RECT 1636.290 1607.900 1636.610 1608.160 ;
        RECT 1636.380 1607.480 1636.520 1607.900 ;
        RECT 1636.290 1607.220 1636.610 1607.480 ;
        RECT 1636.290 1586.820 1636.610 1587.080 ;
        RECT 1636.380 1586.400 1636.520 1586.820 ;
        RECT 1636.290 1586.140 1636.610 1586.400 ;
        RECT 1636.290 1463.060 1636.610 1463.320 ;
        RECT 1636.380 1462.640 1636.520 1463.060 ;
        RECT 1636.290 1462.380 1636.610 1462.640 ;
        RECT 1636.290 1400.700 1636.610 1400.760 ;
        RECT 1636.095 1400.560 1636.610 1400.700 ;
        RECT 1636.290 1400.500 1636.610 1400.560 ;
        RECT 1636.290 1360.920 1636.610 1360.980 ;
        RECT 1636.095 1360.780 1636.610 1360.920 ;
        RECT 1636.290 1360.720 1636.610 1360.780 ;
        RECT 1636.290 1304.140 1636.610 1304.200 ;
        RECT 1636.095 1304.000 1636.610 1304.140 ;
        RECT 1636.290 1303.940 1636.610 1304.000 ;
        RECT 1636.290 1256.200 1636.610 1256.260 ;
        RECT 1636.095 1256.060 1636.610 1256.200 ;
        RECT 1636.290 1256.000 1636.610 1256.060 ;
        RECT 1636.290 1104.220 1636.610 1104.280 ;
        RECT 1637.210 1104.220 1637.530 1104.280 ;
        RECT 1636.290 1104.080 1637.530 1104.220 ;
        RECT 1636.290 1104.020 1636.610 1104.080 ;
        RECT 1637.210 1104.020 1637.530 1104.080 ;
        RECT 1636.290 1014.460 1636.610 1014.520 ;
        RECT 1636.750 1014.460 1637.070 1014.520 ;
        RECT 1636.290 1014.320 1637.070 1014.460 ;
        RECT 1636.290 1014.260 1636.610 1014.320 ;
        RECT 1636.750 1014.260 1637.070 1014.320 ;
        RECT 1636.290 966.180 1636.610 966.240 ;
        RECT 1636.750 966.180 1637.070 966.240 ;
        RECT 1636.290 966.040 1637.070 966.180 ;
        RECT 1636.290 965.980 1636.610 966.040 ;
        RECT 1636.750 965.980 1637.070 966.040 ;
        RECT 1636.290 932.180 1636.610 932.240 ;
        RECT 1635.920 932.040 1636.610 932.180 ;
        RECT 1635.920 931.560 1636.060 932.040 ;
        RECT 1636.290 931.980 1636.610 932.040 ;
        RECT 1635.830 931.300 1636.150 931.560 ;
        RECT 1635.830 869.620 1636.150 869.680 ;
        RECT 1636.290 869.620 1636.610 869.680 ;
        RECT 1635.830 869.480 1636.610 869.620 ;
        RECT 1635.830 869.420 1636.150 869.480 ;
        RECT 1636.290 869.420 1636.610 869.480 ;
        RECT 1635.830 820.800 1636.150 821.060 ;
        RECT 1635.920 820.660 1636.060 820.800 ;
        RECT 1636.290 820.660 1636.610 820.720 ;
        RECT 1635.920 820.520 1636.610 820.660 ;
        RECT 1636.290 820.460 1636.610 820.520 ;
        RECT 1636.290 814.200 1636.610 814.260 ;
        RECT 1637.210 814.200 1637.530 814.260 ;
        RECT 1636.290 814.060 1637.530 814.200 ;
        RECT 1636.290 814.000 1636.610 814.060 ;
        RECT 1637.210 814.000 1637.530 814.060 ;
        RECT 1635.830 620.740 1636.150 620.800 ;
        RECT 1636.290 620.740 1636.610 620.800 ;
        RECT 1635.830 620.600 1636.610 620.740 ;
        RECT 1635.830 620.540 1636.150 620.600 ;
        RECT 1636.290 620.540 1636.610 620.600 ;
        RECT 1636.290 613.940 1636.610 614.000 ;
        RECT 1636.095 613.800 1636.610 613.940 ;
        RECT 1636.290 613.740 1636.610 613.800 ;
        RECT 1636.290 566.000 1636.610 566.060 ;
        RECT 1636.095 565.860 1636.610 566.000 ;
        RECT 1636.290 565.800 1636.610 565.860 ;
        RECT 1636.290 524.860 1636.610 524.920 ;
        RECT 1635.920 524.720 1636.610 524.860 ;
        RECT 1635.920 524.580 1636.060 524.720 ;
        RECT 1636.290 524.660 1636.610 524.720 ;
        RECT 1635.830 524.320 1636.150 524.580 ;
        RECT 1635.830 476.240 1636.150 476.300 ;
        RECT 1636.290 476.240 1636.610 476.300 ;
        RECT 1635.830 476.100 1636.610 476.240 ;
        RECT 1635.830 476.040 1636.150 476.100 ;
        RECT 1636.290 476.040 1636.610 476.100 ;
        RECT 1635.830 427.960 1636.150 428.020 ;
        RECT 1636.290 427.960 1636.610 428.020 ;
        RECT 1635.830 427.820 1636.610 427.960 ;
        RECT 1635.830 427.760 1636.150 427.820 ;
        RECT 1636.290 427.760 1636.610 427.820 ;
        RECT 1635.830 379.680 1636.150 379.740 ;
        RECT 1636.290 379.680 1636.610 379.740 ;
        RECT 1635.830 379.540 1636.610 379.680 ;
        RECT 1635.830 379.480 1636.150 379.540 ;
        RECT 1636.290 379.480 1636.610 379.540 ;
        RECT 1636.290 255.380 1636.610 255.640 ;
        RECT 1636.380 254.960 1636.520 255.380 ;
        RECT 1636.290 254.700 1636.610 254.960 ;
        RECT 1635.830 137.940 1636.150 138.000 ;
        RECT 1636.290 137.940 1636.610 138.000 ;
        RECT 1635.830 137.800 1636.610 137.940 ;
        RECT 1635.830 137.740 1636.150 137.800 ;
        RECT 1636.290 137.740 1636.610 137.800 ;
        RECT 958.710 58.040 959.030 58.100 ;
        RECT 1636.290 58.040 1636.610 58.100 ;
        RECT 958.710 57.900 1636.610 58.040 ;
        RECT 958.710 57.840 959.030 57.900 ;
        RECT 1636.290 57.840 1636.610 57.900 ;
      LAYER via ;
        RECT 1636.320 1659.240 1636.580 1659.500 ;
        RECT 1637.240 1659.240 1637.500 1659.500 ;
        RECT 1636.320 1607.900 1636.580 1608.160 ;
        RECT 1636.320 1607.220 1636.580 1607.480 ;
        RECT 1636.320 1586.820 1636.580 1587.080 ;
        RECT 1636.320 1586.140 1636.580 1586.400 ;
        RECT 1636.320 1463.060 1636.580 1463.320 ;
        RECT 1636.320 1462.380 1636.580 1462.640 ;
        RECT 1636.320 1400.500 1636.580 1400.760 ;
        RECT 1636.320 1360.720 1636.580 1360.980 ;
        RECT 1636.320 1303.940 1636.580 1304.200 ;
        RECT 1636.320 1256.000 1636.580 1256.260 ;
        RECT 1636.320 1104.020 1636.580 1104.280 ;
        RECT 1637.240 1104.020 1637.500 1104.280 ;
        RECT 1636.320 1014.260 1636.580 1014.520 ;
        RECT 1636.780 1014.260 1637.040 1014.520 ;
        RECT 1636.320 965.980 1636.580 966.240 ;
        RECT 1636.780 965.980 1637.040 966.240 ;
        RECT 1636.320 931.980 1636.580 932.240 ;
        RECT 1635.860 931.300 1636.120 931.560 ;
        RECT 1635.860 869.420 1636.120 869.680 ;
        RECT 1636.320 869.420 1636.580 869.680 ;
        RECT 1635.860 820.800 1636.120 821.060 ;
        RECT 1636.320 820.460 1636.580 820.720 ;
        RECT 1636.320 814.000 1636.580 814.260 ;
        RECT 1637.240 814.000 1637.500 814.260 ;
        RECT 1635.860 620.540 1636.120 620.800 ;
        RECT 1636.320 620.540 1636.580 620.800 ;
        RECT 1636.320 613.740 1636.580 614.000 ;
        RECT 1636.320 565.800 1636.580 566.060 ;
        RECT 1636.320 524.660 1636.580 524.920 ;
        RECT 1635.860 524.320 1636.120 524.580 ;
        RECT 1635.860 476.040 1636.120 476.300 ;
        RECT 1636.320 476.040 1636.580 476.300 ;
        RECT 1635.860 427.760 1636.120 428.020 ;
        RECT 1636.320 427.760 1636.580 428.020 ;
        RECT 1635.860 379.480 1636.120 379.740 ;
        RECT 1636.320 379.480 1636.580 379.740 ;
        RECT 1636.320 255.380 1636.580 255.640 ;
        RECT 1636.320 254.700 1636.580 254.960 ;
        RECT 1635.860 137.740 1636.120 138.000 ;
        RECT 1636.320 137.740 1636.580 138.000 ;
        RECT 958.740 57.840 959.000 58.100 ;
        RECT 1636.320 57.840 1636.580 58.100 ;
      LAYER met2 ;
        RECT 1639.460 1700.410 1639.740 1704.000 ;
        RECT 1637.300 1700.270 1639.740 1700.410 ;
        RECT 1637.300 1659.530 1637.440 1700.270 ;
        RECT 1639.460 1700.000 1639.740 1700.270 ;
        RECT 1636.320 1659.210 1636.580 1659.530 ;
        RECT 1637.240 1659.210 1637.500 1659.530 ;
        RECT 1636.380 1608.190 1636.520 1659.210 ;
        RECT 1636.320 1607.870 1636.580 1608.190 ;
        RECT 1636.320 1607.190 1636.580 1607.510 ;
        RECT 1636.380 1587.110 1636.520 1607.190 ;
        RECT 1636.320 1586.790 1636.580 1587.110 ;
        RECT 1636.320 1586.110 1636.580 1586.430 ;
        RECT 1636.380 1463.350 1636.520 1586.110 ;
        RECT 1636.320 1463.030 1636.580 1463.350 ;
        RECT 1636.320 1462.350 1636.580 1462.670 ;
        RECT 1636.380 1400.790 1636.520 1462.350 ;
        RECT 1636.320 1400.470 1636.580 1400.790 ;
        RECT 1636.320 1360.690 1636.580 1361.010 ;
        RECT 1636.380 1304.230 1636.520 1360.690 ;
        RECT 1636.320 1303.910 1636.580 1304.230 ;
        RECT 1636.320 1255.970 1636.580 1256.290 ;
        RECT 1636.380 1152.445 1636.520 1255.970 ;
        RECT 1636.310 1152.075 1636.590 1152.445 ;
        RECT 1637.230 1152.075 1637.510 1152.445 ;
        RECT 1637.300 1104.310 1637.440 1152.075 ;
        RECT 1636.320 1103.990 1636.580 1104.310 ;
        RECT 1637.240 1103.990 1637.500 1104.310 ;
        RECT 1636.380 1014.550 1636.520 1103.990 ;
        RECT 1636.320 1014.230 1636.580 1014.550 ;
        RECT 1636.780 1014.230 1637.040 1014.550 ;
        RECT 1636.840 966.270 1636.980 1014.230 ;
        RECT 1636.320 965.950 1636.580 966.270 ;
        RECT 1636.780 965.950 1637.040 966.270 ;
        RECT 1636.380 932.270 1636.520 965.950 ;
        RECT 1636.320 931.950 1636.580 932.270 ;
        RECT 1635.860 931.270 1636.120 931.590 ;
        RECT 1635.920 869.710 1636.060 931.270 ;
        RECT 1635.860 869.450 1636.120 869.710 ;
        RECT 1636.320 869.450 1636.580 869.710 ;
        RECT 1635.860 869.390 1636.580 869.450 ;
        RECT 1635.920 869.310 1636.520 869.390 ;
        RECT 1635.920 821.090 1636.060 869.310 ;
        RECT 1635.860 820.770 1636.120 821.090 ;
        RECT 1636.320 820.430 1636.580 820.750 ;
        RECT 1636.380 814.290 1636.520 820.430 ;
        RECT 1636.320 813.970 1636.580 814.290 ;
        RECT 1637.240 813.970 1637.500 814.290 ;
        RECT 1637.300 766.205 1637.440 813.970 ;
        RECT 1636.310 765.835 1636.590 766.205 ;
        RECT 1637.230 765.835 1637.510 766.205 ;
        RECT 1636.380 748.410 1636.520 765.835 ;
        RECT 1635.920 748.270 1636.520 748.410 ;
        RECT 1635.920 620.830 1636.060 748.270 ;
        RECT 1635.860 620.510 1636.120 620.830 ;
        RECT 1636.320 620.510 1636.580 620.830 ;
        RECT 1636.380 614.030 1636.520 620.510 ;
        RECT 1636.320 613.710 1636.580 614.030 ;
        RECT 1636.320 565.770 1636.580 566.090 ;
        RECT 1636.380 524.950 1636.520 565.770 ;
        RECT 1636.320 524.630 1636.580 524.950 ;
        RECT 1635.860 524.290 1636.120 524.610 ;
        RECT 1635.920 476.330 1636.060 524.290 ;
        RECT 1635.860 476.010 1636.120 476.330 ;
        RECT 1636.320 476.010 1636.580 476.330 ;
        RECT 1636.380 428.050 1636.520 476.010 ;
        RECT 1635.860 427.730 1636.120 428.050 ;
        RECT 1636.320 427.730 1636.580 428.050 ;
        RECT 1635.920 379.770 1636.060 427.730 ;
        RECT 1635.860 379.450 1636.120 379.770 ;
        RECT 1636.320 379.450 1636.580 379.770 ;
        RECT 1636.380 303.690 1636.520 379.450 ;
        RECT 1635.920 303.550 1636.520 303.690 ;
        RECT 1635.920 303.010 1636.060 303.550 ;
        RECT 1635.920 302.870 1636.520 303.010 ;
        RECT 1636.380 255.670 1636.520 302.870 ;
        RECT 1636.320 255.350 1636.580 255.670 ;
        RECT 1636.320 254.670 1636.580 254.990 ;
        RECT 1636.380 162.250 1636.520 254.670 ;
        RECT 1635.920 162.110 1636.520 162.250 ;
        RECT 1635.920 138.030 1636.060 162.110 ;
        RECT 1635.860 137.710 1636.120 138.030 ;
        RECT 1636.320 137.710 1636.580 138.030 ;
        RECT 1636.380 58.130 1636.520 137.710 ;
        RECT 958.740 57.810 959.000 58.130 ;
        RECT 1636.320 57.810 1636.580 58.130 ;
        RECT 958.800 17.410 958.940 57.810 ;
        RECT 954.200 17.270 958.940 17.410 ;
        RECT 954.200 2.400 954.340 17.270 ;
        RECT 953.990 -4.800 954.550 2.400 ;
      LAYER via2 ;
        RECT 1636.310 1152.120 1636.590 1152.400 ;
        RECT 1637.230 1152.120 1637.510 1152.400 ;
        RECT 1636.310 765.880 1636.590 766.160 ;
        RECT 1637.230 765.880 1637.510 766.160 ;
      LAYER met3 ;
        RECT 1636.285 1152.410 1636.615 1152.425 ;
        RECT 1637.205 1152.410 1637.535 1152.425 ;
        RECT 1636.285 1152.110 1637.535 1152.410 ;
        RECT 1636.285 1152.095 1636.615 1152.110 ;
        RECT 1637.205 1152.095 1637.535 1152.110 ;
        RECT 1636.285 766.170 1636.615 766.185 ;
        RECT 1637.205 766.170 1637.535 766.185 ;
        RECT 1636.285 765.870 1637.535 766.170 ;
        RECT 1636.285 765.855 1636.615 765.870 ;
        RECT 1637.205 765.855 1637.535 765.870 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1643.190 1678.140 1643.510 1678.200 ;
        RECT 1646.870 1678.140 1647.190 1678.200 ;
        RECT 1643.190 1678.000 1647.190 1678.140 ;
        RECT 1643.190 1677.940 1643.510 1678.000 ;
        RECT 1646.870 1677.940 1647.190 1678.000 ;
        RECT 972.510 57.700 972.830 57.760 ;
        RECT 1643.190 57.700 1643.510 57.760 ;
        RECT 972.510 57.560 1643.510 57.700 ;
        RECT 972.510 57.500 972.830 57.560 ;
        RECT 1643.190 57.500 1643.510 57.560 ;
      LAYER via ;
        RECT 1643.220 1677.940 1643.480 1678.200 ;
        RECT 1646.900 1677.940 1647.160 1678.200 ;
        RECT 972.540 57.500 972.800 57.760 ;
        RECT 1643.220 57.500 1643.480 57.760 ;
      LAYER met2 ;
        RECT 1648.660 1700.410 1648.940 1704.000 ;
        RECT 1646.960 1700.270 1648.940 1700.410 ;
        RECT 1646.960 1678.230 1647.100 1700.270 ;
        RECT 1648.660 1700.000 1648.940 1700.270 ;
        RECT 1643.220 1677.910 1643.480 1678.230 ;
        RECT 1646.900 1677.910 1647.160 1678.230 ;
        RECT 1643.280 57.790 1643.420 1677.910 ;
        RECT 972.540 57.470 972.800 57.790 ;
        RECT 1643.220 57.470 1643.480 57.790 ;
        RECT 972.600 17.410 972.740 57.470 ;
        RECT 972.140 17.270 972.740 17.410 ;
        RECT 972.140 2.400 972.280 17.270 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 650.970 26.760 651.290 26.820 ;
        RECT 1483.570 26.760 1483.890 26.820 ;
        RECT 650.970 26.620 1483.890 26.760 ;
        RECT 650.970 26.560 651.290 26.620 ;
        RECT 1483.570 26.560 1483.890 26.620 ;
      LAYER via ;
        RECT 651.000 26.560 651.260 26.820 ;
        RECT 1483.600 26.560 1483.860 26.820 ;
      LAYER met2 ;
        RECT 1483.520 1700.000 1483.800 1704.000 ;
        RECT 1483.660 26.850 1483.800 1700.000 ;
        RECT 651.000 26.530 651.260 26.850 ;
        RECT 1483.600 26.530 1483.860 26.850 ;
        RECT 651.060 2.400 651.200 26.530 ;
        RECT 650.850 -4.800 651.410 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 993.210 57.360 993.530 57.420 ;
        RECT 1656.070 57.360 1656.390 57.420 ;
        RECT 993.210 57.220 1656.390 57.360 ;
        RECT 993.210 57.160 993.530 57.220 ;
        RECT 1656.070 57.160 1656.390 57.220 ;
      LAYER via ;
        RECT 993.240 57.160 993.500 57.420 ;
        RECT 1656.100 57.160 1656.360 57.420 ;
      LAYER met2 ;
        RECT 1657.860 1700.410 1658.140 1704.000 ;
        RECT 1656.160 1700.270 1658.140 1700.410 ;
        RECT 1656.160 57.450 1656.300 1700.270 ;
        RECT 1657.860 1700.000 1658.140 1700.270 ;
        RECT 993.240 57.130 993.500 57.450 ;
        RECT 1656.100 57.130 1656.360 57.450 ;
        RECT 993.300 17.410 993.440 57.130 ;
        RECT 990.080 17.270 993.440 17.410 ;
        RECT 990.080 2.400 990.220 17.270 ;
        RECT 989.870 -4.800 990.430 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1663.965 945.285 1664.135 993.395 ;
      LAYER mcon ;
        RECT 1663.965 993.225 1664.135 993.395 ;
      LAYER met1 ;
        RECT 1663.430 1587.020 1663.750 1587.080 ;
        RECT 1664.350 1587.020 1664.670 1587.080 ;
        RECT 1663.430 1586.880 1664.670 1587.020 ;
        RECT 1663.430 1586.820 1663.750 1586.880 ;
        RECT 1664.350 1586.820 1664.670 1586.880 ;
        RECT 1663.430 1532.280 1663.750 1532.340 ;
        RECT 1664.350 1532.280 1664.670 1532.340 ;
        RECT 1663.430 1532.140 1664.670 1532.280 ;
        RECT 1663.430 1532.080 1663.750 1532.140 ;
        RECT 1664.350 1532.080 1664.670 1532.140 ;
        RECT 1663.890 1483.660 1664.210 1483.720 ;
        RECT 1664.810 1483.660 1665.130 1483.720 ;
        RECT 1663.890 1483.520 1665.130 1483.660 ;
        RECT 1663.890 1483.460 1664.210 1483.520 ;
        RECT 1664.810 1483.460 1665.130 1483.520 ;
        RECT 1664.350 1145.360 1664.670 1145.420 ;
        RECT 1665.270 1145.360 1665.590 1145.420 ;
        RECT 1664.350 1145.220 1665.590 1145.360 ;
        RECT 1664.350 1145.160 1664.670 1145.220 ;
        RECT 1665.270 1145.160 1665.590 1145.220 ;
        RECT 1663.430 1048.800 1663.750 1048.860 ;
        RECT 1664.350 1048.800 1664.670 1048.860 ;
        RECT 1663.430 1048.660 1664.670 1048.800 ;
        RECT 1663.430 1048.600 1663.750 1048.660 ;
        RECT 1664.350 1048.600 1664.670 1048.660 ;
        RECT 1663.890 993.380 1664.210 993.440 ;
        RECT 1663.695 993.240 1664.210 993.380 ;
        RECT 1663.890 993.180 1664.210 993.240 ;
        RECT 1663.890 945.440 1664.210 945.500 ;
        RECT 1663.695 945.300 1664.210 945.440 ;
        RECT 1663.890 945.240 1664.210 945.300 ;
        RECT 1663.890 911.100 1664.210 911.160 ;
        RECT 1663.520 910.960 1664.210 911.100 ;
        RECT 1663.520 910.820 1663.660 910.960 ;
        RECT 1663.890 910.900 1664.210 910.960 ;
        RECT 1663.430 910.560 1663.750 910.820 ;
        RECT 1663.430 862.480 1663.750 862.540 ;
        RECT 1663.890 862.480 1664.210 862.540 ;
        RECT 1663.430 862.340 1664.210 862.480 ;
        RECT 1663.430 862.280 1663.750 862.340 ;
        RECT 1663.890 862.280 1664.210 862.340 ;
        RECT 1663.890 593.340 1664.210 593.600 ;
        RECT 1663.980 592.920 1664.120 593.340 ;
        RECT 1663.890 592.660 1664.210 592.920 ;
        RECT 1663.890 400.220 1664.210 400.480 ;
        RECT 1663.980 399.800 1664.120 400.220 ;
        RECT 1663.890 399.540 1664.210 399.800 ;
        RECT 1663.890 241.980 1664.210 242.040 ;
        RECT 1663.520 241.840 1664.210 241.980 ;
        RECT 1663.520 241.360 1663.660 241.840 ;
        RECT 1663.890 241.780 1664.210 241.840 ;
        RECT 1663.430 241.100 1663.750 241.360 ;
        RECT 1663.430 210.360 1663.750 210.420 ;
        RECT 1664.350 210.360 1664.670 210.420 ;
        RECT 1663.430 210.220 1664.670 210.360 ;
        RECT 1663.430 210.160 1663.750 210.220 ;
        RECT 1664.350 210.160 1664.670 210.220 ;
        RECT 1007.470 57.020 1007.790 57.080 ;
        RECT 1664.350 57.020 1664.670 57.080 ;
        RECT 1007.470 56.880 1664.670 57.020 ;
        RECT 1007.470 56.820 1007.790 56.880 ;
        RECT 1664.350 56.820 1664.670 56.880 ;
      LAYER via ;
        RECT 1663.460 1586.820 1663.720 1587.080 ;
        RECT 1664.380 1586.820 1664.640 1587.080 ;
        RECT 1663.460 1532.080 1663.720 1532.340 ;
        RECT 1664.380 1532.080 1664.640 1532.340 ;
        RECT 1663.920 1483.460 1664.180 1483.720 ;
        RECT 1664.840 1483.460 1665.100 1483.720 ;
        RECT 1664.380 1145.160 1664.640 1145.420 ;
        RECT 1665.300 1145.160 1665.560 1145.420 ;
        RECT 1663.460 1048.600 1663.720 1048.860 ;
        RECT 1664.380 1048.600 1664.640 1048.860 ;
        RECT 1663.920 993.180 1664.180 993.440 ;
        RECT 1663.920 945.240 1664.180 945.500 ;
        RECT 1663.920 910.900 1664.180 911.160 ;
        RECT 1663.460 910.560 1663.720 910.820 ;
        RECT 1663.460 862.280 1663.720 862.540 ;
        RECT 1663.920 862.280 1664.180 862.540 ;
        RECT 1663.920 593.340 1664.180 593.600 ;
        RECT 1663.920 592.660 1664.180 592.920 ;
        RECT 1663.920 400.220 1664.180 400.480 ;
        RECT 1663.920 399.540 1664.180 399.800 ;
        RECT 1663.920 241.780 1664.180 242.040 ;
        RECT 1663.460 241.100 1663.720 241.360 ;
        RECT 1663.460 210.160 1663.720 210.420 ;
        RECT 1664.380 210.160 1664.640 210.420 ;
        RECT 1007.500 56.820 1007.760 57.080 ;
        RECT 1664.380 56.820 1664.640 57.080 ;
      LAYER met2 ;
        RECT 1667.060 1700.410 1667.340 1704.000 ;
        RECT 1665.820 1700.270 1667.340 1700.410 ;
        RECT 1665.820 1690.380 1665.960 1700.270 ;
        RECT 1667.060 1700.000 1667.340 1700.270 ;
        RECT 1663.980 1690.240 1665.960 1690.380 ;
        RECT 1663.980 1642.610 1664.120 1690.240 ;
        RECT 1663.520 1642.470 1664.120 1642.610 ;
        RECT 1663.520 1587.110 1663.660 1642.470 ;
        RECT 1663.460 1586.790 1663.720 1587.110 ;
        RECT 1664.380 1586.790 1664.640 1587.110 ;
        RECT 1664.440 1532.370 1664.580 1586.790 ;
        RECT 1663.460 1532.050 1663.720 1532.370 ;
        RECT 1664.380 1532.050 1664.640 1532.370 ;
        RECT 1663.520 1531.885 1663.660 1532.050 ;
        RECT 1663.450 1531.515 1663.730 1531.885 ;
        RECT 1664.830 1531.515 1665.110 1531.885 ;
        RECT 1664.900 1483.750 1665.040 1531.515 ;
        RECT 1663.920 1483.430 1664.180 1483.750 ;
        RECT 1664.840 1483.430 1665.100 1483.750 ;
        RECT 1663.980 1152.330 1664.120 1483.430 ;
        RECT 1663.980 1152.190 1664.580 1152.330 ;
        RECT 1664.440 1145.450 1664.580 1152.190 ;
        RECT 1664.380 1145.130 1664.640 1145.450 ;
        RECT 1665.300 1145.130 1665.560 1145.450 ;
        RECT 1665.360 1097.365 1665.500 1145.130 ;
        RECT 1663.910 1096.995 1664.190 1097.365 ;
        RECT 1665.290 1096.995 1665.570 1097.365 ;
        RECT 1663.980 1049.650 1664.120 1096.995 ;
        RECT 1663.980 1049.510 1664.580 1049.650 ;
        RECT 1664.440 1048.890 1664.580 1049.510 ;
        RECT 1663.460 1048.570 1663.720 1048.890 ;
        RECT 1664.380 1048.570 1664.640 1048.890 ;
        RECT 1663.520 1001.485 1663.660 1048.570 ;
        RECT 1663.450 1001.115 1663.730 1001.485 ;
        RECT 1663.910 1000.435 1664.190 1000.805 ;
        RECT 1663.980 993.470 1664.120 1000.435 ;
        RECT 1663.920 993.150 1664.180 993.470 ;
        RECT 1663.920 945.210 1664.180 945.530 ;
        RECT 1663.980 911.190 1664.120 945.210 ;
        RECT 1663.920 910.870 1664.180 911.190 ;
        RECT 1663.460 910.530 1663.720 910.850 ;
        RECT 1663.520 862.570 1663.660 910.530 ;
        RECT 1663.460 862.250 1663.720 862.570 ;
        RECT 1663.920 862.250 1664.180 862.570 ;
        RECT 1663.980 786.490 1664.120 862.250 ;
        RECT 1663.520 786.350 1664.120 786.490 ;
        RECT 1663.520 785.130 1663.660 786.350 ;
        RECT 1663.520 784.990 1664.120 785.130 ;
        RECT 1663.980 593.630 1664.120 784.990 ;
        RECT 1663.920 593.310 1664.180 593.630 ;
        RECT 1663.920 592.630 1664.180 592.950 ;
        RECT 1663.980 497.490 1664.120 592.630 ;
        RECT 1663.520 497.350 1664.120 497.490 ;
        RECT 1663.520 496.810 1663.660 497.350 ;
        RECT 1663.520 496.670 1664.120 496.810 ;
        RECT 1663.980 400.510 1664.120 496.670 ;
        RECT 1663.920 400.190 1664.180 400.510 ;
        RECT 1663.920 399.510 1664.180 399.830 ;
        RECT 1663.980 303.690 1664.120 399.510 ;
        RECT 1663.520 303.550 1664.120 303.690 ;
        RECT 1663.520 303.010 1663.660 303.550 ;
        RECT 1663.520 302.870 1664.120 303.010 ;
        RECT 1663.980 242.070 1664.120 302.870 ;
        RECT 1663.920 241.750 1664.180 242.070 ;
        RECT 1663.460 241.070 1663.720 241.390 ;
        RECT 1663.520 210.450 1663.660 241.070 ;
        RECT 1663.460 210.130 1663.720 210.450 ;
        RECT 1664.380 210.130 1664.640 210.450 ;
        RECT 1664.440 57.110 1664.580 210.130 ;
        RECT 1007.500 56.790 1007.760 57.110 ;
        RECT 1664.380 56.790 1664.640 57.110 ;
        RECT 1007.560 2.400 1007.700 56.790 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
      LAYER via2 ;
        RECT 1663.450 1531.560 1663.730 1531.840 ;
        RECT 1664.830 1531.560 1665.110 1531.840 ;
        RECT 1663.910 1097.040 1664.190 1097.320 ;
        RECT 1665.290 1097.040 1665.570 1097.320 ;
        RECT 1663.450 1001.160 1663.730 1001.440 ;
        RECT 1663.910 1000.480 1664.190 1000.760 ;
      LAYER met3 ;
        RECT 1663.425 1531.850 1663.755 1531.865 ;
        RECT 1664.805 1531.850 1665.135 1531.865 ;
        RECT 1663.425 1531.550 1665.135 1531.850 ;
        RECT 1663.425 1531.535 1663.755 1531.550 ;
        RECT 1664.805 1531.535 1665.135 1531.550 ;
        RECT 1663.885 1097.330 1664.215 1097.345 ;
        RECT 1665.265 1097.330 1665.595 1097.345 ;
        RECT 1663.885 1097.030 1665.595 1097.330 ;
        RECT 1663.885 1097.015 1664.215 1097.030 ;
        RECT 1665.265 1097.015 1665.595 1097.030 ;
        RECT 1663.425 1001.450 1663.755 1001.465 ;
        RECT 1663.425 1001.135 1663.970 1001.450 ;
        RECT 1663.670 1000.785 1663.970 1001.135 ;
        RECT 1663.670 1000.470 1664.215 1000.785 ;
        RECT 1663.885 1000.455 1664.215 1000.470 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1671.325 1483.505 1671.495 1490.815 ;
        RECT 1671.325 1413.805 1671.495 1448.995 ;
        RECT 1671.785 1365.865 1671.955 1400.715 ;
        RECT 1671.785 1256.385 1671.955 1304.155 ;
        RECT 1671.785 1220.685 1671.955 1255.875 ;
        RECT 1671.785 1062.245 1671.955 1097.095 ;
        RECT 1672.705 765.765 1672.875 807.075 ;
        RECT 1672.245 710.685 1672.415 758.795 ;
        RECT 1672.245 620.925 1672.415 669.375 ;
        RECT 1671.325 396.525 1671.495 427.635 ;
        RECT 1671.785 324.785 1671.955 372.555 ;
        RECT 1671.785 241.485 1671.955 324.275 ;
        RECT 1671.785 56.525 1671.955 89.675 ;
      LAYER mcon ;
        RECT 1671.325 1490.645 1671.495 1490.815 ;
        RECT 1671.325 1448.825 1671.495 1448.995 ;
        RECT 1671.785 1400.545 1671.955 1400.715 ;
        RECT 1671.785 1303.985 1671.955 1304.155 ;
        RECT 1671.785 1255.705 1671.955 1255.875 ;
        RECT 1671.785 1096.925 1671.955 1097.095 ;
        RECT 1672.705 806.905 1672.875 807.075 ;
        RECT 1672.245 758.625 1672.415 758.795 ;
        RECT 1672.245 669.205 1672.415 669.375 ;
        RECT 1671.325 427.465 1671.495 427.635 ;
        RECT 1671.785 372.385 1671.955 372.555 ;
        RECT 1671.785 324.105 1671.955 324.275 ;
        RECT 1671.785 89.505 1671.955 89.675 ;
      LAYER met1 ;
        RECT 1672.170 1642.440 1672.490 1642.500 ;
        RECT 1674.010 1642.440 1674.330 1642.500 ;
        RECT 1672.170 1642.300 1674.330 1642.440 ;
        RECT 1672.170 1642.240 1672.490 1642.300 ;
        RECT 1674.010 1642.240 1674.330 1642.300 ;
        RECT 1672.170 1587.360 1672.490 1587.420 ;
        RECT 1672.630 1587.360 1672.950 1587.420 ;
        RECT 1672.170 1587.220 1672.950 1587.360 ;
        RECT 1672.170 1587.160 1672.490 1587.220 ;
        RECT 1672.630 1587.160 1672.950 1587.220 ;
        RECT 1671.250 1490.800 1671.570 1490.860 ;
        RECT 1671.055 1490.660 1671.570 1490.800 ;
        RECT 1671.250 1490.600 1671.570 1490.660 ;
        RECT 1671.250 1483.660 1671.570 1483.720 ;
        RECT 1671.055 1483.520 1671.570 1483.660 ;
        RECT 1671.250 1483.460 1671.570 1483.520 ;
        RECT 1671.250 1448.980 1671.570 1449.040 ;
        RECT 1671.055 1448.840 1671.570 1448.980 ;
        RECT 1671.250 1448.780 1671.570 1448.840 ;
        RECT 1671.265 1413.960 1671.555 1414.005 ;
        RECT 1672.170 1413.960 1672.490 1414.020 ;
        RECT 1671.265 1413.820 1672.490 1413.960 ;
        RECT 1671.265 1413.775 1671.555 1413.820 ;
        RECT 1672.170 1413.760 1672.490 1413.820 ;
        RECT 1671.725 1400.700 1672.015 1400.745 ;
        RECT 1672.170 1400.700 1672.490 1400.760 ;
        RECT 1671.725 1400.560 1672.490 1400.700 ;
        RECT 1671.725 1400.515 1672.015 1400.560 ;
        RECT 1672.170 1400.500 1672.490 1400.560 ;
        RECT 1671.710 1366.020 1672.030 1366.080 ;
        RECT 1671.515 1365.880 1672.030 1366.020 ;
        RECT 1671.710 1365.820 1672.030 1365.880 ;
        RECT 1671.710 1317.880 1672.030 1318.140 ;
        RECT 1671.800 1317.400 1671.940 1317.880 ;
        RECT 1672.170 1317.400 1672.490 1317.460 ;
        RECT 1671.800 1317.260 1672.490 1317.400 ;
        RECT 1672.170 1317.200 1672.490 1317.260 ;
        RECT 1671.725 1304.140 1672.015 1304.185 ;
        RECT 1672.170 1304.140 1672.490 1304.200 ;
        RECT 1671.725 1304.000 1672.490 1304.140 ;
        RECT 1671.725 1303.955 1672.015 1304.000 ;
        RECT 1672.170 1303.940 1672.490 1304.000 ;
        RECT 1671.710 1256.540 1672.030 1256.600 ;
        RECT 1671.515 1256.400 1672.030 1256.540 ;
        RECT 1671.710 1256.340 1672.030 1256.400 ;
        RECT 1671.710 1255.860 1672.030 1255.920 ;
        RECT 1671.515 1255.720 1672.030 1255.860 ;
        RECT 1671.710 1255.660 1672.030 1255.720 ;
        RECT 1671.710 1220.840 1672.030 1220.900 ;
        RECT 1671.515 1220.700 1672.030 1220.840 ;
        RECT 1671.710 1220.640 1672.030 1220.700 ;
        RECT 1671.710 1159.980 1672.030 1160.040 ;
        RECT 1671.710 1159.840 1672.400 1159.980 ;
        RECT 1671.710 1159.780 1672.030 1159.840 ;
        RECT 1672.260 1159.360 1672.400 1159.840 ;
        RECT 1672.170 1159.100 1672.490 1159.360 ;
        RECT 1671.710 1097.080 1672.030 1097.140 ;
        RECT 1671.515 1096.940 1672.030 1097.080 ;
        RECT 1671.710 1096.880 1672.030 1096.940 ;
        RECT 1671.725 1062.400 1672.015 1062.445 ;
        RECT 1672.170 1062.400 1672.490 1062.460 ;
        RECT 1671.725 1062.260 1672.490 1062.400 ;
        RECT 1671.725 1062.215 1672.015 1062.260 ;
        RECT 1672.170 1062.200 1672.490 1062.260 ;
        RECT 1671.710 966.180 1672.030 966.240 ;
        RECT 1672.170 966.180 1672.490 966.240 ;
        RECT 1671.710 966.040 1672.490 966.180 ;
        RECT 1671.710 965.980 1672.030 966.040 ;
        RECT 1672.170 965.980 1672.490 966.040 ;
        RECT 1671.710 917.900 1672.030 917.960 ;
        RECT 1672.170 917.900 1672.490 917.960 ;
        RECT 1671.710 917.760 1672.490 917.900 ;
        RECT 1671.710 917.700 1672.030 917.760 ;
        RECT 1672.170 917.700 1672.490 917.760 ;
        RECT 1672.170 910.760 1672.490 910.820 ;
        RECT 1672.630 910.760 1672.950 910.820 ;
        RECT 1672.170 910.620 1672.950 910.760 ;
        RECT 1672.170 910.560 1672.490 910.620 ;
        RECT 1672.630 910.560 1672.950 910.620 ;
        RECT 1672.630 807.060 1672.950 807.120 ;
        RECT 1672.435 806.920 1672.950 807.060 ;
        RECT 1672.630 806.860 1672.950 806.920 ;
        RECT 1672.645 765.920 1672.935 765.965 ;
        RECT 1673.090 765.920 1673.410 765.980 ;
        RECT 1672.645 765.780 1673.410 765.920 ;
        RECT 1672.645 765.735 1672.935 765.780 ;
        RECT 1673.090 765.720 1673.410 765.780 ;
        RECT 1672.185 758.780 1672.475 758.825 ;
        RECT 1673.090 758.780 1673.410 758.840 ;
        RECT 1672.185 758.640 1673.410 758.780 ;
        RECT 1672.185 758.595 1672.475 758.640 ;
        RECT 1673.090 758.580 1673.410 758.640 ;
        RECT 1672.170 710.840 1672.490 710.900 ;
        RECT 1671.975 710.700 1672.490 710.840 ;
        RECT 1672.170 710.640 1672.490 710.700 ;
        RECT 1672.170 669.360 1672.490 669.420 ;
        RECT 1671.975 669.220 1672.490 669.360 ;
        RECT 1672.170 669.160 1672.490 669.220 ;
        RECT 1672.170 621.080 1672.490 621.140 ;
        RECT 1671.975 620.940 1672.490 621.080 ;
        RECT 1672.170 620.880 1672.490 620.940 ;
        RECT 1671.250 435.100 1671.570 435.160 ;
        RECT 1672.170 435.100 1672.490 435.160 ;
        RECT 1671.250 434.960 1672.490 435.100 ;
        RECT 1671.250 434.900 1671.570 434.960 ;
        RECT 1672.170 434.900 1672.490 434.960 ;
        RECT 1671.250 427.620 1671.570 427.680 ;
        RECT 1671.055 427.480 1671.570 427.620 ;
        RECT 1671.250 427.420 1671.570 427.480 ;
        RECT 1671.265 396.680 1671.555 396.725 ;
        RECT 1672.170 396.680 1672.490 396.740 ;
        RECT 1671.265 396.540 1672.490 396.680 ;
        RECT 1671.265 396.495 1671.555 396.540 ;
        RECT 1672.170 396.480 1672.490 396.540 ;
        RECT 1671.725 372.540 1672.015 372.585 ;
        RECT 1672.170 372.540 1672.490 372.600 ;
        RECT 1671.725 372.400 1672.490 372.540 ;
        RECT 1671.725 372.355 1672.015 372.400 ;
        RECT 1672.170 372.340 1672.490 372.400 ;
        RECT 1671.710 324.940 1672.030 325.000 ;
        RECT 1671.515 324.800 1672.030 324.940 ;
        RECT 1671.710 324.740 1672.030 324.800 ;
        RECT 1671.710 324.260 1672.030 324.320 ;
        RECT 1671.515 324.120 1672.030 324.260 ;
        RECT 1671.710 324.060 1672.030 324.120 ;
        RECT 1671.725 241.640 1672.015 241.685 ;
        RECT 1672.170 241.640 1672.490 241.700 ;
        RECT 1671.725 241.500 1672.490 241.640 ;
        RECT 1671.725 241.455 1672.015 241.500 ;
        RECT 1672.170 241.440 1672.490 241.500 ;
        RECT 1671.710 186.560 1672.030 186.620 ;
        RECT 1672.170 186.560 1672.490 186.620 ;
        RECT 1671.710 186.420 1672.490 186.560 ;
        RECT 1671.710 186.360 1672.030 186.420 ;
        RECT 1672.170 186.360 1672.490 186.420 ;
        RECT 1671.710 89.660 1672.030 89.720 ;
        RECT 1671.515 89.520 1672.030 89.660 ;
        RECT 1671.710 89.460 1672.030 89.520 ;
        RECT 1027.710 56.680 1028.030 56.740 ;
        RECT 1671.725 56.680 1672.015 56.725 ;
        RECT 1027.710 56.540 1672.015 56.680 ;
        RECT 1027.710 56.480 1028.030 56.540 ;
        RECT 1671.725 56.495 1672.015 56.540 ;
        RECT 1025.410 2.960 1025.730 3.020 ;
        RECT 1027.710 2.960 1028.030 3.020 ;
        RECT 1025.410 2.820 1028.030 2.960 ;
        RECT 1025.410 2.760 1025.730 2.820 ;
        RECT 1027.710 2.760 1028.030 2.820 ;
      LAYER via ;
        RECT 1672.200 1642.240 1672.460 1642.500 ;
        RECT 1674.040 1642.240 1674.300 1642.500 ;
        RECT 1672.200 1587.160 1672.460 1587.420 ;
        RECT 1672.660 1587.160 1672.920 1587.420 ;
        RECT 1671.280 1490.600 1671.540 1490.860 ;
        RECT 1671.280 1483.460 1671.540 1483.720 ;
        RECT 1671.280 1448.780 1671.540 1449.040 ;
        RECT 1672.200 1413.760 1672.460 1414.020 ;
        RECT 1672.200 1400.500 1672.460 1400.760 ;
        RECT 1671.740 1365.820 1672.000 1366.080 ;
        RECT 1671.740 1317.880 1672.000 1318.140 ;
        RECT 1672.200 1317.200 1672.460 1317.460 ;
        RECT 1672.200 1303.940 1672.460 1304.200 ;
        RECT 1671.740 1256.340 1672.000 1256.600 ;
        RECT 1671.740 1255.660 1672.000 1255.920 ;
        RECT 1671.740 1220.640 1672.000 1220.900 ;
        RECT 1671.740 1159.780 1672.000 1160.040 ;
        RECT 1672.200 1159.100 1672.460 1159.360 ;
        RECT 1671.740 1096.880 1672.000 1097.140 ;
        RECT 1672.200 1062.200 1672.460 1062.460 ;
        RECT 1671.740 965.980 1672.000 966.240 ;
        RECT 1672.200 965.980 1672.460 966.240 ;
        RECT 1671.740 917.700 1672.000 917.960 ;
        RECT 1672.200 917.700 1672.460 917.960 ;
        RECT 1672.200 910.560 1672.460 910.820 ;
        RECT 1672.660 910.560 1672.920 910.820 ;
        RECT 1672.660 806.860 1672.920 807.120 ;
        RECT 1673.120 765.720 1673.380 765.980 ;
        RECT 1673.120 758.580 1673.380 758.840 ;
        RECT 1672.200 710.640 1672.460 710.900 ;
        RECT 1672.200 669.160 1672.460 669.420 ;
        RECT 1672.200 620.880 1672.460 621.140 ;
        RECT 1671.280 434.900 1671.540 435.160 ;
        RECT 1672.200 434.900 1672.460 435.160 ;
        RECT 1671.280 427.420 1671.540 427.680 ;
        RECT 1672.200 396.480 1672.460 396.740 ;
        RECT 1672.200 372.340 1672.460 372.600 ;
        RECT 1671.740 324.740 1672.000 325.000 ;
        RECT 1671.740 324.060 1672.000 324.320 ;
        RECT 1672.200 241.440 1672.460 241.700 ;
        RECT 1671.740 186.360 1672.000 186.620 ;
        RECT 1672.200 186.360 1672.460 186.620 ;
        RECT 1671.740 89.460 1672.000 89.720 ;
        RECT 1027.740 56.480 1028.000 56.740 ;
        RECT 1025.440 2.760 1025.700 3.020 ;
        RECT 1027.740 2.760 1028.000 3.020 ;
      LAYER met2 ;
        RECT 1676.260 1701.090 1676.540 1704.000 ;
        RECT 1674.100 1700.950 1676.540 1701.090 ;
        RECT 1674.100 1642.530 1674.240 1700.950 ;
        RECT 1676.260 1700.000 1676.540 1700.950 ;
        RECT 1672.200 1642.210 1672.460 1642.530 ;
        RECT 1674.040 1642.210 1674.300 1642.530 ;
        RECT 1672.260 1587.450 1672.400 1642.210 ;
        RECT 1672.200 1587.130 1672.460 1587.450 ;
        RECT 1672.660 1587.130 1672.920 1587.450 ;
        RECT 1672.720 1556.250 1672.860 1587.130 ;
        RECT 1671.340 1556.110 1672.860 1556.250 ;
        RECT 1671.340 1490.890 1671.480 1556.110 ;
        RECT 1671.280 1490.570 1671.540 1490.890 ;
        RECT 1671.280 1483.430 1671.540 1483.750 ;
        RECT 1671.340 1449.070 1671.480 1483.430 ;
        RECT 1671.280 1448.750 1671.540 1449.070 ;
        RECT 1672.200 1413.730 1672.460 1414.050 ;
        RECT 1672.260 1400.790 1672.400 1413.730 ;
        RECT 1672.200 1400.470 1672.460 1400.790 ;
        RECT 1671.740 1365.790 1672.000 1366.110 ;
        RECT 1671.800 1318.170 1671.940 1365.790 ;
        RECT 1671.740 1317.850 1672.000 1318.170 ;
        RECT 1672.200 1317.170 1672.460 1317.490 ;
        RECT 1672.260 1304.230 1672.400 1317.170 ;
        RECT 1672.200 1303.910 1672.460 1304.230 ;
        RECT 1671.740 1256.310 1672.000 1256.630 ;
        RECT 1671.800 1255.950 1671.940 1256.310 ;
        RECT 1671.740 1255.630 1672.000 1255.950 ;
        RECT 1671.740 1220.610 1672.000 1220.930 ;
        RECT 1671.800 1160.070 1671.940 1220.610 ;
        RECT 1671.740 1159.750 1672.000 1160.070 ;
        RECT 1672.200 1159.070 1672.460 1159.390 ;
        RECT 1672.260 1134.650 1672.400 1159.070 ;
        RECT 1671.800 1134.510 1672.400 1134.650 ;
        RECT 1671.800 1097.170 1671.940 1134.510 ;
        RECT 1671.740 1096.850 1672.000 1097.170 ;
        RECT 1672.200 1062.170 1672.460 1062.490 ;
        RECT 1672.260 1048.970 1672.400 1062.170 ;
        RECT 1672.260 1048.830 1672.860 1048.970 ;
        RECT 1672.720 1027.890 1672.860 1048.830 ;
        RECT 1672.260 1027.750 1672.860 1027.890 ;
        RECT 1672.260 966.270 1672.400 1027.750 ;
        RECT 1671.740 965.950 1672.000 966.270 ;
        RECT 1672.200 965.950 1672.460 966.270 ;
        RECT 1671.800 917.990 1671.940 965.950 ;
        RECT 1671.740 917.670 1672.000 917.990 ;
        RECT 1672.200 917.670 1672.460 917.990 ;
        RECT 1672.260 910.850 1672.400 917.670 ;
        RECT 1672.200 910.530 1672.460 910.850 ;
        RECT 1672.660 910.530 1672.920 910.850 ;
        RECT 1672.720 807.150 1672.860 910.530 ;
        RECT 1672.660 806.830 1672.920 807.150 ;
        RECT 1673.120 765.690 1673.380 766.010 ;
        RECT 1673.180 758.870 1673.320 765.690 ;
        RECT 1673.120 758.550 1673.380 758.870 ;
        RECT 1672.200 710.610 1672.460 710.930 ;
        RECT 1672.260 669.450 1672.400 710.610 ;
        RECT 1672.200 669.130 1672.460 669.450 ;
        RECT 1672.200 620.850 1672.460 621.170 ;
        RECT 1672.260 596.770 1672.400 620.850 ;
        RECT 1672.260 596.630 1672.860 596.770 ;
        RECT 1672.720 554.610 1672.860 596.630 ;
        RECT 1672.260 554.470 1672.860 554.610 ;
        RECT 1672.260 497.490 1672.400 554.470 ;
        RECT 1672.260 497.350 1672.860 497.490 ;
        RECT 1672.720 482.530 1672.860 497.350 ;
        RECT 1672.260 482.390 1672.860 482.530 ;
        RECT 1672.260 435.190 1672.400 482.390 ;
        RECT 1671.280 434.870 1671.540 435.190 ;
        RECT 1672.200 434.870 1672.460 435.190 ;
        RECT 1671.340 427.710 1671.480 434.870 ;
        RECT 1671.280 427.390 1671.540 427.710 ;
        RECT 1672.200 396.450 1672.460 396.770 ;
        RECT 1672.260 372.630 1672.400 396.450 ;
        RECT 1672.200 372.310 1672.460 372.630 ;
        RECT 1671.740 324.710 1672.000 325.030 ;
        RECT 1671.800 324.350 1671.940 324.710 ;
        RECT 1671.740 324.030 1672.000 324.350 ;
        RECT 1672.200 241.410 1672.460 241.730 ;
        RECT 1672.260 186.650 1672.400 241.410 ;
        RECT 1671.740 186.330 1672.000 186.650 ;
        RECT 1672.200 186.330 1672.460 186.650 ;
        RECT 1671.800 89.750 1671.940 186.330 ;
        RECT 1671.740 89.430 1672.000 89.750 ;
        RECT 1027.740 56.450 1028.000 56.770 ;
        RECT 1027.800 3.050 1027.940 56.450 ;
        RECT 1025.440 2.730 1025.700 3.050 ;
        RECT 1027.740 2.730 1028.000 3.050 ;
        RECT 1025.500 2.400 1025.640 2.730 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1418.250 1686.300 1418.570 1686.360 ;
        RECT 1685.510 1686.300 1685.830 1686.360 ;
        RECT 1418.250 1686.160 1685.830 1686.300 ;
        RECT 1418.250 1686.100 1418.570 1686.160 ;
        RECT 1685.510 1686.100 1685.830 1686.160 ;
        RECT 1043.350 22.680 1043.670 22.740 ;
        RECT 1417.790 22.680 1418.110 22.740 ;
        RECT 1043.350 22.540 1418.110 22.680 ;
        RECT 1043.350 22.480 1043.670 22.540 ;
        RECT 1417.790 22.480 1418.110 22.540 ;
      LAYER via ;
        RECT 1418.280 1686.100 1418.540 1686.360 ;
        RECT 1685.540 1686.100 1685.800 1686.360 ;
        RECT 1043.380 22.480 1043.640 22.740 ;
        RECT 1417.820 22.480 1418.080 22.740 ;
      LAYER met2 ;
        RECT 1685.460 1700.000 1685.740 1704.000 ;
        RECT 1685.600 1686.390 1685.740 1700.000 ;
        RECT 1418.280 1686.070 1418.540 1686.390 ;
        RECT 1685.540 1686.070 1685.800 1686.390 ;
        RECT 1418.340 39.850 1418.480 1686.070 ;
        RECT 1417.880 39.710 1418.480 39.850 ;
        RECT 1417.880 22.770 1418.020 39.710 ;
        RECT 1043.380 22.450 1043.640 22.770 ;
        RECT 1417.820 22.450 1418.080 22.770 ;
        RECT 1043.440 2.400 1043.580 22.450 ;
        RECT 1043.230 -4.800 1043.790 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1424.690 1686.640 1425.010 1686.700 ;
        RECT 1694.710 1686.640 1695.030 1686.700 ;
        RECT 1424.690 1686.500 1695.030 1686.640 ;
        RECT 1424.690 1686.440 1425.010 1686.500 ;
        RECT 1694.710 1686.440 1695.030 1686.500 ;
        RECT 1061.290 22.340 1061.610 22.400 ;
        RECT 1424.690 22.340 1425.010 22.400 ;
        RECT 1061.290 22.200 1425.010 22.340 ;
        RECT 1061.290 22.140 1061.610 22.200 ;
        RECT 1424.690 22.140 1425.010 22.200 ;
      LAYER via ;
        RECT 1424.720 1686.440 1424.980 1686.700 ;
        RECT 1694.740 1686.440 1695.000 1686.700 ;
        RECT 1061.320 22.140 1061.580 22.400 ;
        RECT 1424.720 22.140 1424.980 22.400 ;
      LAYER met2 ;
        RECT 1694.660 1700.000 1694.940 1704.000 ;
        RECT 1694.800 1686.730 1694.940 1700.000 ;
        RECT 1424.720 1686.410 1424.980 1686.730 ;
        RECT 1694.740 1686.410 1695.000 1686.730 ;
        RECT 1424.780 22.430 1424.920 1686.410 ;
        RECT 1061.320 22.110 1061.580 22.430 ;
        RECT 1424.720 22.110 1424.980 22.430 ;
        RECT 1061.380 2.400 1061.520 22.110 ;
        RECT 1061.170 -4.800 1061.730 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1697.470 1666.240 1697.790 1666.300 ;
        RECT 1702.070 1666.240 1702.390 1666.300 ;
        RECT 1697.470 1666.100 1702.390 1666.240 ;
        RECT 1697.470 1666.040 1697.790 1666.100 ;
        RECT 1702.070 1666.040 1702.390 1666.100 ;
        RECT 1079.230 23.700 1079.550 23.760 ;
        RECT 1697.470 23.700 1697.790 23.760 ;
        RECT 1079.230 23.560 1697.790 23.700 ;
        RECT 1079.230 23.500 1079.550 23.560 ;
        RECT 1697.470 23.500 1697.790 23.560 ;
      LAYER via ;
        RECT 1697.500 1666.040 1697.760 1666.300 ;
        RECT 1702.100 1666.040 1702.360 1666.300 ;
        RECT 1079.260 23.500 1079.520 23.760 ;
        RECT 1697.500 23.500 1697.760 23.760 ;
      LAYER met2 ;
        RECT 1703.860 1700.410 1704.140 1704.000 ;
        RECT 1702.160 1700.270 1704.140 1700.410 ;
        RECT 1702.160 1666.330 1702.300 1700.270 ;
        RECT 1703.860 1700.000 1704.140 1700.270 ;
        RECT 1697.500 1666.010 1697.760 1666.330 ;
        RECT 1702.100 1666.010 1702.360 1666.330 ;
        RECT 1697.560 23.790 1697.700 1666.010 ;
        RECT 1079.260 23.470 1079.520 23.790 ;
        RECT 1697.500 23.470 1697.760 23.790 ;
        RECT 1079.320 2.400 1079.460 23.470 ;
        RECT 1079.110 -4.800 1079.670 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1713.060 1700.410 1713.340 1704.000 ;
        RECT 1711.360 1700.270 1713.340 1700.410 ;
        RECT 1711.360 24.325 1711.500 1700.270 ;
        RECT 1713.060 1700.000 1713.340 1700.270 ;
        RECT 1096.730 23.955 1097.010 24.325 ;
        RECT 1711.290 23.955 1711.570 24.325 ;
        RECT 1096.800 2.400 1096.940 23.955 ;
        RECT 1096.590 -4.800 1097.150 2.400 ;
      LAYER via2 ;
        RECT 1096.730 24.000 1097.010 24.280 ;
        RECT 1711.290 24.000 1711.570 24.280 ;
      LAYER met3 ;
        RECT 1096.705 24.290 1097.035 24.305 ;
        RECT 1711.265 24.290 1711.595 24.305 ;
        RECT 1096.705 23.990 1711.595 24.290 ;
        RECT 1096.705 23.975 1097.035 23.990 ;
        RECT 1711.265 23.975 1711.595 23.990 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1718.170 1661.140 1718.490 1661.200 ;
        RECT 1720.470 1661.140 1720.790 1661.200 ;
        RECT 1718.170 1661.000 1720.790 1661.140 ;
        RECT 1718.170 1660.940 1718.490 1661.000 ;
        RECT 1720.470 1660.940 1720.790 1661.000 ;
        RECT 1114.650 23.360 1114.970 23.420 ;
        RECT 1718.170 23.360 1718.490 23.420 ;
        RECT 1114.650 23.220 1718.490 23.360 ;
        RECT 1114.650 23.160 1114.970 23.220 ;
        RECT 1718.170 23.160 1718.490 23.220 ;
      LAYER via ;
        RECT 1718.200 1660.940 1718.460 1661.200 ;
        RECT 1720.500 1660.940 1720.760 1661.200 ;
        RECT 1114.680 23.160 1114.940 23.420 ;
        RECT 1718.200 23.160 1718.460 23.420 ;
      LAYER met2 ;
        RECT 1722.260 1700.410 1722.540 1704.000 ;
        RECT 1720.560 1700.270 1722.540 1700.410 ;
        RECT 1720.560 1661.230 1720.700 1700.270 ;
        RECT 1722.260 1700.000 1722.540 1700.270 ;
        RECT 1718.200 1660.910 1718.460 1661.230 ;
        RECT 1720.500 1660.910 1720.760 1661.230 ;
        RECT 1718.260 23.450 1718.400 1660.910 ;
        RECT 1114.680 23.130 1114.940 23.450 ;
        RECT 1718.200 23.130 1718.460 23.450 ;
        RECT 1114.740 2.400 1114.880 23.130 ;
        RECT 1114.530 -4.800 1115.090 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1725.070 1678.140 1725.390 1678.200 ;
        RECT 1729.670 1678.140 1729.990 1678.200 ;
        RECT 1725.070 1678.000 1729.990 1678.140 ;
        RECT 1725.070 1677.940 1725.390 1678.000 ;
        RECT 1729.670 1677.940 1729.990 1678.000 ;
        RECT 1132.590 23.020 1132.910 23.080 ;
        RECT 1725.070 23.020 1725.390 23.080 ;
        RECT 1132.590 22.880 1725.390 23.020 ;
        RECT 1132.590 22.820 1132.910 22.880 ;
        RECT 1725.070 22.820 1725.390 22.880 ;
      LAYER via ;
        RECT 1725.100 1677.940 1725.360 1678.200 ;
        RECT 1729.700 1677.940 1729.960 1678.200 ;
        RECT 1132.620 22.820 1132.880 23.080 ;
        RECT 1725.100 22.820 1725.360 23.080 ;
      LAYER met2 ;
        RECT 1731.460 1700.410 1731.740 1704.000 ;
        RECT 1729.760 1700.270 1731.740 1700.410 ;
        RECT 1729.760 1678.230 1729.900 1700.270 ;
        RECT 1731.460 1700.000 1731.740 1700.270 ;
        RECT 1725.100 1677.910 1725.360 1678.230 ;
        RECT 1729.700 1677.910 1729.960 1678.230 ;
        RECT 1725.160 23.110 1725.300 1677.910 ;
        RECT 1132.620 22.790 1132.880 23.110 ;
        RECT 1725.100 22.790 1725.360 23.110 ;
        RECT 1132.680 2.400 1132.820 22.790 ;
        RECT 1132.470 -4.800 1133.030 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1150.530 24.040 1150.850 24.100 ;
        RECT 1738.870 24.040 1739.190 24.100 ;
        RECT 1150.530 23.900 1739.190 24.040 ;
        RECT 1150.530 23.840 1150.850 23.900 ;
        RECT 1738.870 23.840 1739.190 23.900 ;
      LAYER via ;
        RECT 1150.560 23.840 1150.820 24.100 ;
        RECT 1738.900 23.840 1739.160 24.100 ;
      LAYER met2 ;
        RECT 1740.660 1700.410 1740.940 1704.000 ;
        RECT 1738.960 1700.270 1740.940 1700.410 ;
        RECT 1738.960 24.130 1739.100 1700.270 ;
        RECT 1740.660 1700.000 1740.940 1700.270 ;
        RECT 1150.560 23.810 1150.820 24.130 ;
        RECT 1738.900 23.810 1739.160 24.130 ;
        RECT 1150.620 2.400 1150.760 23.810 ;
        RECT 1150.410 -4.800 1150.970 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 668.910 27.100 669.230 27.160 ;
        RECT 1490.470 27.100 1490.790 27.160 ;
        RECT 668.910 26.960 1490.790 27.100 ;
        RECT 668.910 26.900 669.230 26.960 ;
        RECT 1490.470 26.900 1490.790 26.960 ;
      LAYER via ;
        RECT 668.940 26.900 669.200 27.160 ;
        RECT 1490.500 26.900 1490.760 27.160 ;
      LAYER met2 ;
        RECT 1492.720 1700.410 1493.000 1704.000 ;
        RECT 1490.560 1700.270 1493.000 1700.410 ;
        RECT 1490.560 27.190 1490.700 1700.270 ;
        RECT 1492.720 1700.000 1493.000 1700.270 ;
        RECT 668.940 26.870 669.200 27.190 ;
        RECT 1490.500 26.870 1490.760 27.190 ;
        RECT 669.000 2.400 669.140 26.870 ;
        RECT 668.790 -4.800 669.350 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1745.770 1678.140 1746.090 1678.200 ;
        RECT 1748.070 1678.140 1748.390 1678.200 ;
        RECT 1745.770 1678.000 1748.390 1678.140 ;
        RECT 1745.770 1677.940 1746.090 1678.000 ;
        RECT 1748.070 1677.940 1748.390 1678.000 ;
        RECT 1168.470 24.380 1168.790 24.440 ;
        RECT 1745.770 24.380 1746.090 24.440 ;
        RECT 1168.470 24.240 1746.090 24.380 ;
        RECT 1168.470 24.180 1168.790 24.240 ;
        RECT 1745.770 24.180 1746.090 24.240 ;
      LAYER via ;
        RECT 1745.800 1677.940 1746.060 1678.200 ;
        RECT 1748.100 1677.940 1748.360 1678.200 ;
        RECT 1168.500 24.180 1168.760 24.440 ;
        RECT 1745.800 24.180 1746.060 24.440 ;
      LAYER met2 ;
        RECT 1749.860 1700.410 1750.140 1704.000 ;
        RECT 1748.160 1700.270 1750.140 1700.410 ;
        RECT 1748.160 1678.230 1748.300 1700.270 ;
        RECT 1749.860 1700.000 1750.140 1700.270 ;
        RECT 1745.800 1677.910 1746.060 1678.230 ;
        RECT 1748.100 1677.910 1748.360 1678.230 ;
        RECT 1745.860 24.470 1746.000 1677.910 ;
        RECT 1168.500 24.150 1168.760 24.470 ;
        RECT 1745.800 24.150 1746.060 24.470 ;
        RECT 1168.560 2.400 1168.700 24.150 ;
        RECT 1168.350 -4.800 1168.910 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1752.670 1678.140 1752.990 1678.200 ;
        RECT 1757.270 1678.140 1757.590 1678.200 ;
        RECT 1752.670 1678.000 1757.590 1678.140 ;
        RECT 1752.670 1677.940 1752.990 1678.000 ;
        RECT 1757.270 1677.940 1757.590 1678.000 ;
        RECT 1185.950 24.720 1186.270 24.780 ;
        RECT 1752.670 24.720 1752.990 24.780 ;
        RECT 1185.950 24.580 1752.990 24.720 ;
        RECT 1185.950 24.520 1186.270 24.580 ;
        RECT 1752.670 24.520 1752.990 24.580 ;
      LAYER via ;
        RECT 1752.700 1677.940 1752.960 1678.200 ;
        RECT 1757.300 1677.940 1757.560 1678.200 ;
        RECT 1185.980 24.520 1186.240 24.780 ;
        RECT 1752.700 24.520 1752.960 24.780 ;
      LAYER met2 ;
        RECT 1759.060 1700.410 1759.340 1704.000 ;
        RECT 1757.360 1700.270 1759.340 1700.410 ;
        RECT 1757.360 1678.230 1757.500 1700.270 ;
        RECT 1759.060 1700.000 1759.340 1700.270 ;
        RECT 1752.700 1677.910 1752.960 1678.230 ;
        RECT 1757.300 1677.910 1757.560 1678.230 ;
        RECT 1752.760 24.810 1752.900 1677.910 ;
        RECT 1185.980 24.490 1186.240 24.810 ;
        RECT 1752.700 24.490 1752.960 24.810 ;
        RECT 1186.040 2.400 1186.180 24.490 ;
        RECT 1185.830 -4.800 1186.390 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1203.890 25.060 1204.210 25.120 ;
        RECT 1766.470 25.060 1766.790 25.120 ;
        RECT 1203.890 24.920 1766.790 25.060 ;
        RECT 1203.890 24.860 1204.210 24.920 ;
        RECT 1766.470 24.860 1766.790 24.920 ;
      LAYER via ;
        RECT 1203.920 24.860 1204.180 25.120 ;
        RECT 1766.500 24.860 1766.760 25.120 ;
      LAYER met2 ;
        RECT 1768.260 1700.410 1768.540 1704.000 ;
        RECT 1766.560 1700.270 1768.540 1700.410 ;
        RECT 1766.560 25.150 1766.700 1700.270 ;
        RECT 1768.260 1700.000 1768.540 1700.270 ;
        RECT 1203.920 24.830 1204.180 25.150 ;
        RECT 1766.500 24.830 1766.760 25.150 ;
        RECT 1203.980 2.400 1204.120 24.830 ;
        RECT 1203.770 -4.800 1204.330 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1773.370 1678.140 1773.690 1678.200 ;
        RECT 1775.670 1678.140 1775.990 1678.200 ;
        RECT 1773.370 1678.000 1775.990 1678.140 ;
        RECT 1773.370 1677.940 1773.690 1678.000 ;
        RECT 1775.670 1677.940 1775.990 1678.000 ;
        RECT 1221.830 25.400 1222.150 25.460 ;
        RECT 1773.370 25.400 1773.690 25.460 ;
        RECT 1221.830 25.260 1773.690 25.400 ;
        RECT 1221.830 25.200 1222.150 25.260 ;
        RECT 1773.370 25.200 1773.690 25.260 ;
      LAYER via ;
        RECT 1773.400 1677.940 1773.660 1678.200 ;
        RECT 1775.700 1677.940 1775.960 1678.200 ;
        RECT 1221.860 25.200 1222.120 25.460 ;
        RECT 1773.400 25.200 1773.660 25.460 ;
      LAYER met2 ;
        RECT 1777.460 1700.410 1777.740 1704.000 ;
        RECT 1775.760 1700.270 1777.740 1700.410 ;
        RECT 1775.760 1678.230 1775.900 1700.270 ;
        RECT 1777.460 1700.000 1777.740 1700.270 ;
        RECT 1773.400 1677.910 1773.660 1678.230 ;
        RECT 1775.700 1677.910 1775.960 1678.230 ;
        RECT 1773.460 25.490 1773.600 1677.910 ;
        RECT 1221.860 25.170 1222.120 25.490 ;
        RECT 1773.400 25.170 1773.660 25.490 ;
        RECT 1221.920 2.400 1222.060 25.170 ;
        RECT 1221.710 -4.800 1222.270 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1782.645 1587.205 1782.815 1676.455 ;
        RECT 1782.185 1352.265 1782.355 1366.715 ;
        RECT 1782.185 758.965 1782.355 806.735 ;
        RECT 1782.185 620.925 1782.355 669.375 ;
        RECT 1782.185 365.925 1782.355 414.035 ;
        RECT 1782.645 227.885 1782.815 317.475 ;
        RECT 1783.105 179.605 1783.275 203.915 ;
        RECT 1782.645 131.665 1782.815 155.635 ;
      LAYER mcon ;
        RECT 1782.645 1676.285 1782.815 1676.455 ;
        RECT 1782.185 1366.545 1782.355 1366.715 ;
        RECT 1782.185 806.565 1782.355 806.735 ;
        RECT 1782.185 669.205 1782.355 669.375 ;
        RECT 1782.185 413.865 1782.355 414.035 ;
        RECT 1782.645 317.305 1782.815 317.475 ;
        RECT 1783.105 203.745 1783.275 203.915 ;
        RECT 1782.645 155.465 1782.815 155.635 ;
      LAYER met1 ;
        RECT 1783.490 1692.080 1783.810 1692.140 ;
        RECT 1786.710 1692.080 1787.030 1692.140 ;
        RECT 1783.490 1691.940 1787.030 1692.080 ;
        RECT 1783.490 1691.880 1783.810 1691.940 ;
        RECT 1786.710 1691.880 1787.030 1691.940 ;
        RECT 1782.570 1683.580 1782.890 1683.640 ;
        RECT 1783.490 1683.580 1783.810 1683.640 ;
        RECT 1782.570 1683.440 1783.810 1683.580 ;
        RECT 1782.570 1683.380 1782.890 1683.440 ;
        RECT 1783.490 1683.380 1783.810 1683.440 ;
        RECT 1782.570 1676.440 1782.890 1676.500 ;
        RECT 1782.375 1676.300 1782.890 1676.440 ;
        RECT 1782.570 1676.240 1782.890 1676.300 ;
        RECT 1782.570 1587.360 1782.890 1587.420 ;
        RECT 1782.375 1587.220 1782.890 1587.360 ;
        RECT 1782.570 1587.160 1782.890 1587.220 ;
        RECT 1782.110 1448.780 1782.430 1449.040 ;
        RECT 1782.200 1448.640 1782.340 1448.780 ;
        RECT 1782.570 1448.640 1782.890 1448.700 ;
        RECT 1782.200 1448.500 1782.890 1448.640 ;
        RECT 1782.570 1448.440 1782.890 1448.500 ;
        RECT 1782.110 1387.100 1782.430 1387.160 ;
        RECT 1783.490 1387.100 1783.810 1387.160 ;
        RECT 1782.110 1386.960 1783.810 1387.100 ;
        RECT 1782.110 1386.900 1782.430 1386.960 ;
        RECT 1783.490 1386.900 1783.810 1386.960 ;
        RECT 1782.110 1366.700 1782.430 1366.760 ;
        RECT 1781.915 1366.560 1782.430 1366.700 ;
        RECT 1782.110 1366.500 1782.430 1366.560 ;
        RECT 1782.110 1352.420 1782.430 1352.480 ;
        RECT 1781.915 1352.280 1782.430 1352.420 ;
        RECT 1782.110 1352.220 1782.430 1352.280 ;
        RECT 1782.110 1318.220 1782.430 1318.480 ;
        RECT 1782.200 1317.740 1782.340 1318.220 ;
        RECT 1782.570 1317.740 1782.890 1317.800 ;
        RECT 1782.200 1317.600 1782.890 1317.740 ;
        RECT 1782.570 1317.540 1782.890 1317.600 ;
        RECT 1782.110 1290.200 1782.430 1290.260 ;
        RECT 1783.030 1290.200 1783.350 1290.260 ;
        RECT 1782.110 1290.060 1783.350 1290.200 ;
        RECT 1782.110 1290.000 1782.430 1290.060 ;
        RECT 1783.030 1290.000 1783.350 1290.060 ;
        RECT 1781.650 1241.920 1781.970 1241.980 ;
        RECT 1782.110 1241.920 1782.430 1241.980 ;
        RECT 1781.650 1241.780 1782.430 1241.920 ;
        RECT 1781.650 1241.720 1781.970 1241.780 ;
        RECT 1782.110 1241.720 1782.430 1241.780 ;
        RECT 1782.570 1193.300 1782.890 1193.360 ;
        RECT 1783.030 1193.300 1783.350 1193.360 ;
        RECT 1782.570 1193.160 1783.350 1193.300 ;
        RECT 1782.570 1193.100 1782.890 1193.160 ;
        RECT 1783.030 1193.100 1783.350 1193.160 ;
        RECT 1782.570 1063.080 1782.890 1063.140 ;
        RECT 1782.200 1062.940 1782.890 1063.080 ;
        RECT 1782.200 1062.800 1782.340 1062.940 ;
        RECT 1782.570 1062.880 1782.890 1062.940 ;
        RECT 1782.110 1062.540 1782.430 1062.800 ;
        RECT 1782.570 966.520 1782.890 966.580 ;
        RECT 1782.200 966.380 1782.890 966.520 ;
        RECT 1782.200 966.240 1782.340 966.380 ;
        RECT 1782.570 966.320 1782.890 966.380 ;
        RECT 1782.110 965.980 1782.430 966.240 ;
        RECT 1782.110 917.900 1782.430 917.960 ;
        RECT 1782.570 917.900 1782.890 917.960 ;
        RECT 1782.110 917.760 1782.890 917.900 ;
        RECT 1782.110 917.700 1782.430 917.760 ;
        RECT 1782.570 917.700 1782.890 917.760 ;
        RECT 1782.570 835.620 1782.890 835.680 ;
        RECT 1782.200 835.480 1782.890 835.620 ;
        RECT 1782.200 834.660 1782.340 835.480 ;
        RECT 1782.570 835.420 1782.890 835.480 ;
        RECT 1782.110 834.400 1782.430 834.660 ;
        RECT 1782.110 806.720 1782.430 806.780 ;
        RECT 1781.915 806.580 1782.430 806.720 ;
        RECT 1782.110 806.520 1782.430 806.580 ;
        RECT 1782.110 759.120 1782.430 759.180 ;
        RECT 1781.915 758.980 1782.430 759.120 ;
        RECT 1782.110 758.920 1782.430 758.980 ;
        RECT 1782.110 669.360 1782.430 669.420 ;
        RECT 1781.915 669.220 1782.430 669.360 ;
        RECT 1782.110 669.160 1782.430 669.220 ;
        RECT 1782.110 621.080 1782.430 621.140 ;
        RECT 1781.915 620.940 1782.430 621.080 ;
        RECT 1782.110 620.880 1782.430 620.940 ;
        RECT 1782.110 572.940 1782.430 573.200 ;
        RECT 1782.200 572.800 1782.340 572.940 ;
        RECT 1782.570 572.800 1782.890 572.860 ;
        RECT 1782.200 572.660 1782.890 572.800 ;
        RECT 1782.570 572.600 1782.890 572.660 ;
        RECT 1783.030 517.180 1783.350 517.440 ;
        RECT 1782.110 517.040 1782.430 517.100 ;
        RECT 1783.120 517.040 1783.260 517.180 ;
        RECT 1782.110 516.900 1783.260 517.040 ;
        RECT 1782.110 516.840 1782.430 516.900 ;
        RECT 1782.110 448.500 1782.430 448.760 ;
        RECT 1782.200 448.020 1782.340 448.500 ;
        RECT 1782.570 448.020 1782.890 448.080 ;
        RECT 1782.200 447.880 1782.890 448.020 ;
        RECT 1782.570 447.820 1782.890 447.880 ;
        RECT 1782.570 420.620 1782.890 420.880 ;
        RECT 1782.660 420.200 1782.800 420.620 ;
        RECT 1782.570 419.940 1782.890 420.200 ;
        RECT 1782.125 414.020 1782.415 414.065 ;
        RECT 1782.570 414.020 1782.890 414.080 ;
        RECT 1782.125 413.880 1782.890 414.020 ;
        RECT 1782.125 413.835 1782.415 413.880 ;
        RECT 1782.570 413.820 1782.890 413.880 ;
        RECT 1782.110 366.080 1782.430 366.140 ;
        RECT 1781.915 365.940 1782.430 366.080 ;
        RECT 1782.110 365.880 1782.430 365.940 ;
        RECT 1782.110 324.260 1782.430 324.320 ;
        RECT 1783.030 324.260 1783.350 324.320 ;
        RECT 1782.110 324.120 1783.350 324.260 ;
        RECT 1782.110 324.060 1782.430 324.120 ;
        RECT 1783.030 324.060 1783.350 324.120 ;
        RECT 1782.585 317.460 1782.875 317.505 ;
        RECT 1783.030 317.460 1783.350 317.520 ;
        RECT 1782.585 317.320 1783.350 317.460 ;
        RECT 1782.585 317.275 1782.875 317.320 ;
        RECT 1783.030 317.260 1783.350 317.320 ;
        RECT 1782.570 228.040 1782.890 228.100 ;
        RECT 1782.375 227.900 1782.890 228.040 ;
        RECT 1782.570 227.840 1782.890 227.900 ;
        RECT 1782.570 203.900 1782.890 203.960 ;
        RECT 1783.045 203.900 1783.335 203.945 ;
        RECT 1782.570 203.760 1783.335 203.900 ;
        RECT 1782.570 203.700 1782.890 203.760 ;
        RECT 1783.045 203.715 1783.335 203.760 ;
        RECT 1783.030 179.760 1783.350 179.820 ;
        RECT 1782.835 179.620 1783.350 179.760 ;
        RECT 1783.030 179.560 1783.350 179.620 ;
        RECT 1782.585 155.620 1782.875 155.665 ;
        RECT 1783.030 155.620 1783.350 155.680 ;
        RECT 1782.585 155.480 1783.350 155.620 ;
        RECT 1782.585 155.435 1782.875 155.480 ;
        RECT 1783.030 155.420 1783.350 155.480 ;
        RECT 1782.570 131.820 1782.890 131.880 ;
        RECT 1782.375 131.680 1782.890 131.820 ;
        RECT 1782.570 131.620 1782.890 131.680 ;
        RECT 1781.650 76.060 1781.970 76.120 ;
        RECT 1782.110 76.060 1782.430 76.120 ;
        RECT 1781.650 75.920 1782.430 76.060 ;
        RECT 1781.650 75.860 1781.970 75.920 ;
        RECT 1782.110 75.860 1782.430 75.920 ;
        RECT 1239.770 25.740 1240.090 25.800 ;
        RECT 1782.110 25.740 1782.430 25.800 ;
        RECT 1239.770 25.600 1782.430 25.740 ;
        RECT 1239.770 25.540 1240.090 25.600 ;
        RECT 1782.110 25.540 1782.430 25.600 ;
      LAYER via ;
        RECT 1783.520 1691.880 1783.780 1692.140 ;
        RECT 1786.740 1691.880 1787.000 1692.140 ;
        RECT 1782.600 1683.380 1782.860 1683.640 ;
        RECT 1783.520 1683.380 1783.780 1683.640 ;
        RECT 1782.600 1676.240 1782.860 1676.500 ;
        RECT 1782.600 1587.160 1782.860 1587.420 ;
        RECT 1782.140 1448.780 1782.400 1449.040 ;
        RECT 1782.600 1448.440 1782.860 1448.700 ;
        RECT 1782.140 1386.900 1782.400 1387.160 ;
        RECT 1783.520 1386.900 1783.780 1387.160 ;
        RECT 1782.140 1366.500 1782.400 1366.760 ;
        RECT 1782.140 1352.220 1782.400 1352.480 ;
        RECT 1782.140 1318.220 1782.400 1318.480 ;
        RECT 1782.600 1317.540 1782.860 1317.800 ;
        RECT 1782.140 1290.000 1782.400 1290.260 ;
        RECT 1783.060 1290.000 1783.320 1290.260 ;
        RECT 1781.680 1241.720 1781.940 1241.980 ;
        RECT 1782.140 1241.720 1782.400 1241.980 ;
        RECT 1782.600 1193.100 1782.860 1193.360 ;
        RECT 1783.060 1193.100 1783.320 1193.360 ;
        RECT 1782.600 1062.880 1782.860 1063.140 ;
        RECT 1782.140 1062.540 1782.400 1062.800 ;
        RECT 1782.600 966.320 1782.860 966.580 ;
        RECT 1782.140 965.980 1782.400 966.240 ;
        RECT 1782.140 917.700 1782.400 917.960 ;
        RECT 1782.600 917.700 1782.860 917.960 ;
        RECT 1782.600 835.420 1782.860 835.680 ;
        RECT 1782.140 834.400 1782.400 834.660 ;
        RECT 1782.140 806.520 1782.400 806.780 ;
        RECT 1782.140 758.920 1782.400 759.180 ;
        RECT 1782.140 669.160 1782.400 669.420 ;
        RECT 1782.140 620.880 1782.400 621.140 ;
        RECT 1782.140 572.940 1782.400 573.200 ;
        RECT 1782.600 572.600 1782.860 572.860 ;
        RECT 1783.060 517.180 1783.320 517.440 ;
        RECT 1782.140 516.840 1782.400 517.100 ;
        RECT 1782.140 448.500 1782.400 448.760 ;
        RECT 1782.600 447.820 1782.860 448.080 ;
        RECT 1782.600 420.620 1782.860 420.880 ;
        RECT 1782.600 419.940 1782.860 420.200 ;
        RECT 1782.600 413.820 1782.860 414.080 ;
        RECT 1782.140 365.880 1782.400 366.140 ;
        RECT 1782.140 324.060 1782.400 324.320 ;
        RECT 1783.060 324.060 1783.320 324.320 ;
        RECT 1783.060 317.260 1783.320 317.520 ;
        RECT 1782.600 227.840 1782.860 228.100 ;
        RECT 1782.600 203.700 1782.860 203.960 ;
        RECT 1783.060 179.560 1783.320 179.820 ;
        RECT 1783.060 155.420 1783.320 155.680 ;
        RECT 1782.600 131.620 1782.860 131.880 ;
        RECT 1781.680 75.860 1781.940 76.120 ;
        RECT 1782.140 75.860 1782.400 76.120 ;
        RECT 1239.800 25.540 1240.060 25.800 ;
        RECT 1782.140 25.540 1782.400 25.800 ;
      LAYER met2 ;
        RECT 1786.660 1700.000 1786.940 1704.000 ;
        RECT 1786.800 1692.170 1786.940 1700.000 ;
        RECT 1783.520 1691.850 1783.780 1692.170 ;
        RECT 1786.740 1691.850 1787.000 1692.170 ;
        RECT 1783.580 1683.670 1783.720 1691.850 ;
        RECT 1782.600 1683.350 1782.860 1683.670 ;
        RECT 1783.520 1683.350 1783.780 1683.670 ;
        RECT 1782.660 1676.530 1782.800 1683.350 ;
        RECT 1782.600 1676.210 1782.860 1676.530 ;
        RECT 1782.600 1587.130 1782.860 1587.450 ;
        RECT 1782.660 1521.570 1782.800 1587.130 ;
        RECT 1782.660 1521.430 1783.260 1521.570 ;
        RECT 1783.120 1449.490 1783.260 1521.430 ;
        RECT 1782.200 1449.350 1783.260 1449.490 ;
        RECT 1782.200 1449.070 1782.340 1449.350 ;
        RECT 1782.140 1448.750 1782.400 1449.070 ;
        RECT 1782.600 1448.410 1782.860 1448.730 ;
        RECT 1782.660 1442.125 1782.800 1448.410 ;
        RECT 1782.590 1441.755 1782.870 1442.125 ;
        RECT 1783.510 1441.755 1783.790 1442.125 ;
        RECT 1783.580 1387.190 1783.720 1441.755 ;
        RECT 1782.140 1386.870 1782.400 1387.190 ;
        RECT 1783.520 1386.870 1783.780 1387.190 ;
        RECT 1782.200 1366.790 1782.340 1386.870 ;
        RECT 1782.140 1366.470 1782.400 1366.790 ;
        RECT 1782.140 1352.190 1782.400 1352.510 ;
        RECT 1782.200 1318.510 1782.340 1352.190 ;
        RECT 1782.140 1318.190 1782.400 1318.510 ;
        RECT 1782.600 1317.510 1782.860 1317.830 ;
        RECT 1782.660 1297.850 1782.800 1317.510 ;
        RECT 1782.200 1297.710 1782.800 1297.850 ;
        RECT 1782.200 1290.290 1782.340 1297.710 ;
        RECT 1782.140 1289.970 1782.400 1290.290 ;
        RECT 1783.060 1289.970 1783.320 1290.290 ;
        RECT 1783.120 1242.205 1783.260 1289.970 ;
        RECT 1781.680 1241.690 1781.940 1242.010 ;
        RECT 1782.130 1241.835 1782.410 1242.205 ;
        RECT 1783.050 1241.835 1783.330 1242.205 ;
        RECT 1782.140 1241.690 1782.400 1241.835 ;
        RECT 1781.740 1193.925 1781.880 1241.690 ;
        RECT 1781.670 1193.555 1781.950 1193.925 ;
        RECT 1782.590 1193.555 1782.870 1193.925 ;
        RECT 1782.660 1193.390 1782.800 1193.555 ;
        RECT 1782.600 1193.070 1782.860 1193.390 ;
        RECT 1783.060 1193.070 1783.320 1193.390 ;
        RECT 1783.120 1169.330 1783.260 1193.070 ;
        RECT 1782.660 1169.190 1783.260 1169.330 ;
        RECT 1782.660 1063.170 1782.800 1169.190 ;
        RECT 1782.600 1062.850 1782.860 1063.170 ;
        RECT 1782.140 1062.685 1782.400 1062.830 ;
        RECT 1782.130 1062.315 1782.410 1062.685 ;
        RECT 1783.050 1062.315 1783.330 1062.685 ;
        RECT 1783.120 1024.490 1783.260 1062.315 ;
        RECT 1782.200 1024.350 1783.260 1024.490 ;
        RECT 1782.200 1013.610 1782.340 1024.350 ;
        RECT 1782.200 1013.470 1782.800 1013.610 ;
        RECT 1782.660 966.610 1782.800 1013.470 ;
        RECT 1782.600 966.290 1782.860 966.610 ;
        RECT 1782.140 965.950 1782.400 966.270 ;
        RECT 1782.200 917.990 1782.340 965.950 ;
        RECT 1782.140 917.670 1782.400 917.990 ;
        RECT 1782.600 917.670 1782.860 917.990 ;
        RECT 1782.660 835.710 1782.800 917.670 ;
        RECT 1782.600 835.390 1782.860 835.710 ;
        RECT 1782.140 834.370 1782.400 834.690 ;
        RECT 1782.200 806.810 1782.340 834.370 ;
        RECT 1782.140 806.490 1782.400 806.810 ;
        RECT 1782.140 758.890 1782.400 759.210 ;
        RECT 1782.200 724.725 1782.340 758.890 ;
        RECT 1782.130 724.355 1782.410 724.725 ;
        RECT 1782.130 723.675 1782.410 724.045 ;
        RECT 1782.200 670.325 1782.340 723.675 ;
        RECT 1782.130 669.955 1782.410 670.325 ;
        RECT 1782.130 669.275 1782.410 669.645 ;
        RECT 1782.140 669.130 1782.400 669.275 ;
        RECT 1782.140 620.850 1782.400 621.170 ;
        RECT 1782.200 573.230 1782.340 620.850 ;
        RECT 1782.140 572.910 1782.400 573.230 ;
        RECT 1782.600 572.570 1782.860 572.890 ;
        RECT 1782.660 524.010 1782.800 572.570 ;
        RECT 1782.660 523.870 1783.260 524.010 ;
        RECT 1783.120 517.470 1783.260 523.870 ;
        RECT 1783.060 517.150 1783.320 517.470 ;
        RECT 1782.140 516.810 1782.400 517.130 ;
        RECT 1782.200 470.405 1782.340 516.810 ;
        RECT 1782.130 470.035 1782.410 470.405 ;
        RECT 1782.130 469.355 1782.410 469.725 ;
        RECT 1782.200 448.790 1782.340 469.355 ;
        RECT 1782.140 448.470 1782.400 448.790 ;
        RECT 1782.600 447.790 1782.860 448.110 ;
        RECT 1782.660 420.910 1782.800 447.790 ;
        RECT 1782.600 420.590 1782.860 420.910 ;
        RECT 1782.600 419.910 1782.860 420.230 ;
        RECT 1782.660 414.110 1782.800 419.910 ;
        RECT 1782.600 413.790 1782.860 414.110 ;
        RECT 1782.140 365.850 1782.400 366.170 ;
        RECT 1782.200 324.350 1782.340 365.850 ;
        RECT 1782.140 324.030 1782.400 324.350 ;
        RECT 1783.060 324.030 1783.320 324.350 ;
        RECT 1783.120 317.550 1783.260 324.030 ;
        RECT 1783.060 317.230 1783.320 317.550 ;
        RECT 1782.600 227.810 1782.860 228.130 ;
        RECT 1782.660 203.990 1782.800 227.810 ;
        RECT 1782.600 203.670 1782.860 203.990 ;
        RECT 1783.060 179.530 1783.320 179.850 ;
        RECT 1783.120 155.710 1783.260 179.530 ;
        RECT 1783.060 155.390 1783.320 155.710 ;
        RECT 1782.600 131.590 1782.860 131.910 ;
        RECT 1782.660 124.285 1782.800 131.590 ;
        RECT 1781.670 123.915 1781.950 124.285 ;
        RECT 1782.590 123.915 1782.870 124.285 ;
        RECT 1781.740 76.150 1781.880 123.915 ;
        RECT 1781.680 75.830 1781.940 76.150 ;
        RECT 1782.140 75.830 1782.400 76.150 ;
        RECT 1782.200 25.830 1782.340 75.830 ;
        RECT 1239.800 25.510 1240.060 25.830 ;
        RECT 1782.140 25.510 1782.400 25.830 ;
        RECT 1239.860 2.400 1240.000 25.510 ;
        RECT 1239.650 -4.800 1240.210 2.400 ;
      LAYER via2 ;
        RECT 1782.590 1441.800 1782.870 1442.080 ;
        RECT 1783.510 1441.800 1783.790 1442.080 ;
        RECT 1782.130 1241.880 1782.410 1242.160 ;
        RECT 1783.050 1241.880 1783.330 1242.160 ;
        RECT 1781.670 1193.600 1781.950 1193.880 ;
        RECT 1782.590 1193.600 1782.870 1193.880 ;
        RECT 1782.130 1062.360 1782.410 1062.640 ;
        RECT 1783.050 1062.360 1783.330 1062.640 ;
        RECT 1782.130 724.400 1782.410 724.680 ;
        RECT 1782.130 723.720 1782.410 724.000 ;
        RECT 1782.130 670.000 1782.410 670.280 ;
        RECT 1782.130 669.320 1782.410 669.600 ;
        RECT 1782.130 470.080 1782.410 470.360 ;
        RECT 1782.130 469.400 1782.410 469.680 ;
        RECT 1781.670 123.960 1781.950 124.240 ;
        RECT 1782.590 123.960 1782.870 124.240 ;
      LAYER met3 ;
        RECT 1782.565 1442.090 1782.895 1442.105 ;
        RECT 1783.485 1442.090 1783.815 1442.105 ;
        RECT 1782.565 1441.790 1783.815 1442.090 ;
        RECT 1782.565 1441.775 1782.895 1441.790 ;
        RECT 1783.485 1441.775 1783.815 1441.790 ;
        RECT 1782.105 1242.170 1782.435 1242.185 ;
        RECT 1783.025 1242.170 1783.355 1242.185 ;
        RECT 1782.105 1241.870 1783.355 1242.170 ;
        RECT 1782.105 1241.855 1782.435 1241.870 ;
        RECT 1783.025 1241.855 1783.355 1241.870 ;
        RECT 1781.645 1193.890 1781.975 1193.905 ;
        RECT 1782.565 1193.890 1782.895 1193.905 ;
        RECT 1781.645 1193.590 1782.895 1193.890 ;
        RECT 1781.645 1193.575 1781.975 1193.590 ;
        RECT 1782.565 1193.575 1782.895 1193.590 ;
        RECT 1782.105 1062.650 1782.435 1062.665 ;
        RECT 1783.025 1062.650 1783.355 1062.665 ;
        RECT 1782.105 1062.350 1783.355 1062.650 ;
        RECT 1782.105 1062.335 1782.435 1062.350 ;
        RECT 1783.025 1062.335 1783.355 1062.350 ;
        RECT 1782.105 724.690 1782.435 724.705 ;
        RECT 1781.430 724.390 1782.435 724.690 ;
        RECT 1781.430 724.010 1781.730 724.390 ;
        RECT 1782.105 724.375 1782.435 724.390 ;
        RECT 1782.105 724.010 1782.435 724.025 ;
        RECT 1781.430 723.710 1782.435 724.010 ;
        RECT 1782.105 723.695 1782.435 723.710 ;
        RECT 1782.105 670.290 1782.435 670.305 ;
        RECT 1782.105 669.975 1782.650 670.290 ;
        RECT 1782.350 669.625 1782.650 669.975 ;
        RECT 1782.105 669.310 1782.650 669.625 ;
        RECT 1782.105 669.295 1782.435 669.310 ;
        RECT 1782.105 470.055 1782.435 470.385 ;
        RECT 1782.120 469.705 1782.420 470.055 ;
        RECT 1782.105 469.375 1782.435 469.705 ;
        RECT 1781.645 124.250 1781.975 124.265 ;
        RECT 1782.565 124.250 1782.895 124.265 ;
        RECT 1781.645 123.950 1782.895 124.250 ;
        RECT 1781.645 123.935 1781.975 123.950 ;
        RECT 1782.565 123.935 1782.895 123.950 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1257.250 26.080 1257.570 26.140 ;
        RECT 1794.070 26.080 1794.390 26.140 ;
        RECT 1257.250 25.940 1794.390 26.080 ;
        RECT 1257.250 25.880 1257.570 25.940 ;
        RECT 1794.070 25.880 1794.390 25.940 ;
      LAYER via ;
        RECT 1257.280 25.880 1257.540 26.140 ;
        RECT 1794.100 25.880 1794.360 26.140 ;
      LAYER met2 ;
        RECT 1795.860 1700.410 1796.140 1704.000 ;
        RECT 1794.160 1700.270 1796.140 1700.410 ;
        RECT 1794.160 26.170 1794.300 1700.270 ;
        RECT 1795.860 1700.000 1796.140 1700.270 ;
        RECT 1257.280 25.850 1257.540 26.170 ;
        RECT 1794.100 25.850 1794.360 26.170 ;
        RECT 1257.340 2.400 1257.480 25.850 ;
        RECT 1257.130 -4.800 1257.690 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1800.970 1678.140 1801.290 1678.200 ;
        RECT 1803.270 1678.140 1803.590 1678.200 ;
        RECT 1800.970 1678.000 1803.590 1678.140 ;
        RECT 1800.970 1677.940 1801.290 1678.000 ;
        RECT 1803.270 1677.940 1803.590 1678.000 ;
        RECT 1626.630 29.480 1626.950 29.540 ;
        RECT 1800.970 29.480 1801.290 29.540 ;
        RECT 1626.630 29.340 1801.290 29.480 ;
        RECT 1626.630 29.280 1626.950 29.340 ;
        RECT 1800.970 29.280 1801.290 29.340 ;
        RECT 1275.190 19.280 1275.510 19.340 ;
        RECT 1275.190 19.140 1583.620 19.280 ;
        RECT 1275.190 19.080 1275.510 19.140 ;
        RECT 1583.480 18.600 1583.620 19.140 ;
        RECT 1626.630 18.600 1626.950 18.660 ;
        RECT 1583.480 18.460 1626.950 18.600 ;
        RECT 1626.630 18.400 1626.950 18.460 ;
      LAYER via ;
        RECT 1801.000 1677.940 1801.260 1678.200 ;
        RECT 1803.300 1677.940 1803.560 1678.200 ;
        RECT 1626.660 29.280 1626.920 29.540 ;
        RECT 1801.000 29.280 1801.260 29.540 ;
        RECT 1275.220 19.080 1275.480 19.340 ;
        RECT 1626.660 18.400 1626.920 18.660 ;
      LAYER met2 ;
        RECT 1805.060 1700.410 1805.340 1704.000 ;
        RECT 1803.360 1700.270 1805.340 1700.410 ;
        RECT 1803.360 1678.230 1803.500 1700.270 ;
        RECT 1805.060 1700.000 1805.340 1700.270 ;
        RECT 1801.000 1677.910 1801.260 1678.230 ;
        RECT 1803.300 1677.910 1803.560 1678.230 ;
        RECT 1801.060 29.570 1801.200 1677.910 ;
        RECT 1626.660 29.250 1626.920 29.570 ;
        RECT 1801.000 29.250 1801.260 29.570 ;
        RECT 1275.220 19.050 1275.480 19.370 ;
        RECT 1275.280 2.400 1275.420 19.050 ;
        RECT 1626.720 18.690 1626.860 29.250 ;
        RECT 1626.660 18.370 1626.920 18.690 ;
        RECT 1275.070 -4.800 1275.630 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1808.330 1678.140 1808.650 1678.200 ;
        RECT 1812.470 1678.140 1812.790 1678.200 ;
        RECT 1808.330 1678.000 1812.790 1678.140 ;
        RECT 1808.330 1677.940 1808.650 1678.000 ;
        RECT 1812.470 1677.940 1812.790 1678.000 ;
        RECT 1808.330 46.480 1808.650 46.540 ;
        RECT 1626.720 46.340 1808.650 46.480 ;
        RECT 1612.830 45.800 1613.150 45.860 ;
        RECT 1626.720 45.800 1626.860 46.340 ;
        RECT 1808.330 46.280 1808.650 46.340 ;
        RECT 1612.830 45.660 1626.860 45.800 ;
        RECT 1612.830 45.600 1613.150 45.660 ;
        RECT 1293.130 19.620 1293.450 19.680 ;
        RECT 1612.830 19.620 1613.150 19.680 ;
        RECT 1293.130 19.480 1613.150 19.620 ;
        RECT 1293.130 19.420 1293.450 19.480 ;
        RECT 1612.830 19.420 1613.150 19.480 ;
      LAYER via ;
        RECT 1808.360 1677.940 1808.620 1678.200 ;
        RECT 1812.500 1677.940 1812.760 1678.200 ;
        RECT 1612.860 45.600 1613.120 45.860 ;
        RECT 1808.360 46.280 1808.620 46.540 ;
        RECT 1293.160 19.420 1293.420 19.680 ;
        RECT 1612.860 19.420 1613.120 19.680 ;
      LAYER met2 ;
        RECT 1814.260 1700.410 1814.540 1704.000 ;
        RECT 1812.560 1700.270 1814.540 1700.410 ;
        RECT 1812.560 1678.230 1812.700 1700.270 ;
        RECT 1814.260 1700.000 1814.540 1700.270 ;
        RECT 1808.360 1677.910 1808.620 1678.230 ;
        RECT 1812.500 1677.910 1812.760 1678.230 ;
        RECT 1808.420 46.570 1808.560 1677.910 ;
        RECT 1808.360 46.250 1808.620 46.570 ;
        RECT 1612.860 45.570 1613.120 45.890 ;
        RECT 1612.920 19.710 1613.060 45.570 ;
        RECT 1293.160 19.390 1293.420 19.710 ;
        RECT 1612.860 19.390 1613.120 19.710 ;
        RECT 1293.220 2.400 1293.360 19.390 ;
        RECT 1293.010 -4.800 1293.570 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1821.745 1061.905 1821.915 1064.115 ;
      LAYER mcon ;
        RECT 1821.745 1063.945 1821.915 1064.115 ;
      LAYER met1 ;
        RECT 1821.670 1064.100 1821.990 1064.160 ;
        RECT 1821.670 1063.960 1822.185 1064.100 ;
        RECT 1821.670 1063.900 1821.990 1063.960 ;
        RECT 1821.670 1062.060 1821.990 1062.120 ;
        RECT 1821.670 1061.920 1822.185 1062.060 ;
        RECT 1821.670 1061.860 1821.990 1061.920 ;
        RECT 1821.670 905.120 1821.990 905.380 ;
        RECT 1821.760 904.360 1821.900 905.120 ;
        RECT 1821.670 904.100 1821.990 904.360 ;
        RECT 1613.290 29.140 1613.610 29.200 ;
        RECT 1821.670 29.140 1821.990 29.200 ;
        RECT 1613.290 29.000 1821.990 29.140 ;
        RECT 1613.290 28.940 1613.610 29.000 ;
        RECT 1821.670 28.940 1821.990 29.000 ;
        RECT 1311.070 20.300 1311.390 20.360 ;
        RECT 1613.290 20.300 1613.610 20.360 ;
        RECT 1311.070 20.160 1613.610 20.300 ;
        RECT 1311.070 20.100 1311.390 20.160 ;
        RECT 1613.290 20.100 1613.610 20.160 ;
      LAYER via ;
        RECT 1821.700 1063.900 1821.960 1064.160 ;
        RECT 1821.700 1061.860 1821.960 1062.120 ;
        RECT 1821.700 905.120 1821.960 905.380 ;
        RECT 1821.700 904.100 1821.960 904.360 ;
        RECT 1613.320 28.940 1613.580 29.200 ;
        RECT 1821.700 28.940 1821.960 29.200 ;
        RECT 1311.100 20.100 1311.360 20.360 ;
        RECT 1613.320 20.100 1613.580 20.360 ;
      LAYER met2 ;
        RECT 1823.460 1700.410 1823.740 1704.000 ;
        RECT 1821.760 1700.270 1823.740 1700.410 ;
        RECT 1821.760 1064.190 1821.900 1700.270 ;
        RECT 1823.460 1700.000 1823.740 1700.270 ;
        RECT 1821.700 1063.870 1821.960 1064.190 ;
        RECT 1821.700 1061.830 1821.960 1062.150 ;
        RECT 1821.760 905.410 1821.900 1061.830 ;
        RECT 1821.700 905.090 1821.960 905.410 ;
        RECT 1821.700 904.070 1821.960 904.390 ;
        RECT 1821.760 29.230 1821.900 904.070 ;
        RECT 1613.320 28.910 1613.580 29.230 ;
        RECT 1821.700 28.910 1821.960 29.230 ;
        RECT 1613.380 20.390 1613.520 28.910 ;
        RECT 1311.100 20.070 1311.360 20.390 ;
        RECT 1613.320 20.070 1613.580 20.390 ;
        RECT 1311.160 2.400 1311.300 20.070 ;
        RECT 1310.950 -4.800 1311.510 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1829.565 593.045 1829.735 620.755 ;
      LAYER mcon ;
        RECT 1829.565 620.585 1829.735 620.755 ;
      LAYER met1 ;
        RECT 1829.030 1593.820 1829.350 1593.880 ;
        RECT 1829.490 1593.820 1829.810 1593.880 ;
        RECT 1829.030 1593.680 1829.810 1593.820 ;
        RECT 1829.030 1593.620 1829.350 1593.680 ;
        RECT 1829.490 1593.620 1829.810 1593.680 ;
        RECT 1829.030 1587.020 1829.350 1587.080 ;
        RECT 1829.490 1587.020 1829.810 1587.080 ;
        RECT 1829.030 1586.880 1829.810 1587.020 ;
        RECT 1829.030 1586.820 1829.350 1586.880 ;
        RECT 1829.490 1586.820 1829.810 1586.880 ;
        RECT 1829.490 1400.700 1829.810 1400.760 ;
        RECT 1829.950 1400.700 1830.270 1400.760 ;
        RECT 1829.490 1400.560 1830.270 1400.700 ;
        RECT 1829.490 1400.500 1829.810 1400.560 ;
        RECT 1829.950 1400.500 1830.270 1400.560 ;
        RECT 1828.570 983.180 1828.890 983.240 ;
        RECT 1829.490 983.180 1829.810 983.240 ;
        RECT 1828.570 983.040 1829.810 983.180 ;
        RECT 1828.570 982.980 1828.890 983.040 ;
        RECT 1829.490 982.980 1829.810 983.040 ;
        RECT 1828.570 910.760 1828.890 910.820 ;
        RECT 1829.490 910.760 1829.810 910.820 ;
        RECT 1828.570 910.620 1829.810 910.760 ;
        RECT 1828.570 910.560 1828.890 910.620 ;
        RECT 1829.490 910.560 1829.810 910.620 ;
        RECT 1829.950 676.500 1830.270 676.560 ;
        RECT 1829.580 676.360 1830.270 676.500 ;
        RECT 1829.580 676.220 1829.720 676.360 ;
        RECT 1829.950 676.300 1830.270 676.360 ;
        RECT 1829.490 675.960 1829.810 676.220 ;
        RECT 1829.490 628.220 1829.810 628.280 ;
        RECT 1829.950 628.220 1830.270 628.280 ;
        RECT 1829.490 628.080 1830.270 628.220 ;
        RECT 1829.490 628.020 1829.810 628.080 ;
        RECT 1829.950 628.020 1830.270 628.080 ;
        RECT 1829.490 620.740 1829.810 620.800 ;
        RECT 1829.295 620.600 1829.810 620.740 ;
        RECT 1829.490 620.540 1829.810 620.600 ;
        RECT 1829.490 593.200 1829.810 593.260 ;
        RECT 1829.295 593.060 1829.810 593.200 ;
        RECT 1829.490 593.000 1829.810 593.060 ;
        RECT 1829.490 400.220 1829.810 400.480 ;
        RECT 1829.580 399.800 1829.720 400.220 ;
        RECT 1829.490 399.540 1829.810 399.800 ;
        RECT 1828.570 113.800 1828.890 113.860 ;
        RECT 1829.950 113.800 1830.270 113.860 ;
        RECT 1828.570 113.660 1830.270 113.800 ;
        RECT 1828.570 113.600 1828.890 113.660 ;
        RECT 1829.950 113.600 1830.270 113.660 ;
        RECT 1438.030 52.600 1438.350 52.660 ;
        RECT 1828.570 52.600 1828.890 52.660 ;
        RECT 1438.030 52.460 1828.890 52.600 ;
        RECT 1438.030 52.400 1438.350 52.460 ;
        RECT 1828.570 52.400 1828.890 52.460 ;
        RECT 1329.010 17.580 1329.330 17.640 ;
        RECT 1438.030 17.580 1438.350 17.640 ;
        RECT 1329.010 17.440 1438.350 17.580 ;
        RECT 1329.010 17.380 1329.330 17.440 ;
        RECT 1438.030 17.380 1438.350 17.440 ;
      LAYER via ;
        RECT 1829.060 1593.620 1829.320 1593.880 ;
        RECT 1829.520 1593.620 1829.780 1593.880 ;
        RECT 1829.060 1586.820 1829.320 1587.080 ;
        RECT 1829.520 1586.820 1829.780 1587.080 ;
        RECT 1829.520 1400.500 1829.780 1400.760 ;
        RECT 1829.980 1400.500 1830.240 1400.760 ;
        RECT 1828.600 982.980 1828.860 983.240 ;
        RECT 1829.520 982.980 1829.780 983.240 ;
        RECT 1828.600 910.560 1828.860 910.820 ;
        RECT 1829.520 910.560 1829.780 910.820 ;
        RECT 1829.980 676.300 1830.240 676.560 ;
        RECT 1829.520 675.960 1829.780 676.220 ;
        RECT 1829.520 628.020 1829.780 628.280 ;
        RECT 1829.980 628.020 1830.240 628.280 ;
        RECT 1829.520 620.540 1829.780 620.800 ;
        RECT 1829.520 593.000 1829.780 593.260 ;
        RECT 1829.520 400.220 1829.780 400.480 ;
        RECT 1829.520 399.540 1829.780 399.800 ;
        RECT 1828.600 113.600 1828.860 113.860 ;
        RECT 1829.980 113.600 1830.240 113.860 ;
        RECT 1438.060 52.400 1438.320 52.660 ;
        RECT 1828.600 52.400 1828.860 52.660 ;
        RECT 1329.040 17.380 1329.300 17.640 ;
        RECT 1438.060 17.380 1438.320 17.640 ;
      LAYER met2 ;
        RECT 1832.660 1700.410 1832.940 1704.000 ;
        RECT 1830.040 1700.270 1832.940 1700.410 ;
        RECT 1830.040 1642.610 1830.180 1700.270 ;
        RECT 1832.660 1700.000 1832.940 1700.270 ;
        RECT 1829.580 1642.470 1830.180 1642.610 ;
        RECT 1829.580 1593.910 1829.720 1642.470 ;
        RECT 1829.060 1593.590 1829.320 1593.910 ;
        RECT 1829.520 1593.590 1829.780 1593.910 ;
        RECT 1829.120 1587.110 1829.260 1593.590 ;
        RECT 1829.060 1586.790 1829.320 1587.110 ;
        RECT 1829.520 1586.790 1829.780 1587.110 ;
        RECT 1829.580 1463.090 1829.720 1586.790 ;
        RECT 1829.120 1462.950 1829.720 1463.090 ;
        RECT 1829.120 1462.410 1829.260 1462.950 ;
        RECT 1829.120 1462.270 1829.720 1462.410 ;
        RECT 1829.580 1400.790 1829.720 1462.270 ;
        RECT 1829.520 1400.470 1829.780 1400.790 ;
        RECT 1829.980 1400.470 1830.240 1400.790 ;
        RECT 1830.040 1366.020 1830.180 1400.470 ;
        RECT 1829.580 1365.880 1830.180 1366.020 ;
        RECT 1829.580 1269.970 1829.720 1365.880 ;
        RECT 1829.120 1269.830 1829.720 1269.970 ;
        RECT 1829.120 1269.290 1829.260 1269.830 ;
        RECT 1829.120 1269.150 1829.720 1269.290 ;
        RECT 1829.580 983.270 1829.720 1269.150 ;
        RECT 1828.600 982.950 1828.860 983.270 ;
        RECT 1829.520 982.950 1829.780 983.270 ;
        RECT 1828.660 959.325 1828.800 982.950 ;
        RECT 1828.590 958.955 1828.870 959.325 ;
        RECT 1829.510 958.955 1829.790 959.325 ;
        RECT 1829.580 910.850 1829.720 958.955 ;
        RECT 1828.600 910.530 1828.860 910.850 ;
        RECT 1829.520 910.530 1829.780 910.850 ;
        RECT 1828.660 862.765 1828.800 910.530 ;
        RECT 1828.590 862.395 1828.870 862.765 ;
        RECT 1829.510 862.395 1829.790 862.765 ;
        RECT 1829.580 786.490 1829.720 862.395 ;
        RECT 1829.120 786.350 1829.720 786.490 ;
        RECT 1829.120 785.130 1829.260 786.350 ;
        RECT 1829.120 784.990 1829.720 785.130 ;
        RECT 1829.580 693.330 1829.720 784.990 ;
        RECT 1829.580 693.190 1830.180 693.330 ;
        RECT 1830.040 676.590 1830.180 693.190 ;
        RECT 1829.980 676.270 1830.240 676.590 ;
        RECT 1829.520 675.930 1829.780 676.250 ;
        RECT 1829.580 669.530 1829.720 675.930 ;
        RECT 1829.580 669.390 1830.180 669.530 ;
        RECT 1830.040 628.310 1830.180 669.390 ;
        RECT 1829.520 627.990 1829.780 628.310 ;
        RECT 1829.980 627.990 1830.240 628.310 ;
        RECT 1829.580 620.830 1829.720 627.990 ;
        RECT 1829.520 620.510 1829.780 620.830 ;
        RECT 1829.520 592.970 1829.780 593.290 ;
        RECT 1829.580 400.510 1829.720 592.970 ;
        RECT 1829.520 400.190 1829.780 400.510 ;
        RECT 1829.520 399.510 1829.780 399.830 ;
        RECT 1829.580 303.690 1829.720 399.510 ;
        RECT 1829.120 303.550 1829.720 303.690 ;
        RECT 1829.120 303.010 1829.260 303.550 ;
        RECT 1829.120 302.870 1829.720 303.010 ;
        RECT 1829.580 235.010 1829.720 302.870 ;
        RECT 1829.120 234.870 1829.720 235.010 ;
        RECT 1829.120 203.730 1829.260 234.870 ;
        RECT 1829.120 203.590 1829.720 203.730 ;
        RECT 1829.580 137.770 1829.720 203.590 ;
        RECT 1829.580 137.630 1830.180 137.770 ;
        RECT 1830.040 113.890 1830.180 137.630 ;
        RECT 1828.600 113.570 1828.860 113.890 ;
        RECT 1829.980 113.570 1830.240 113.890 ;
        RECT 1828.660 52.690 1828.800 113.570 ;
        RECT 1438.060 52.370 1438.320 52.690 ;
        RECT 1828.600 52.370 1828.860 52.690 ;
        RECT 1438.120 17.670 1438.260 52.370 ;
        RECT 1329.040 17.350 1329.300 17.670 ;
        RECT 1438.060 17.350 1438.320 17.670 ;
        RECT 1329.100 2.400 1329.240 17.350 ;
        RECT 1328.890 -4.800 1329.450 2.400 ;
      LAYER via2 ;
        RECT 1828.590 959.000 1828.870 959.280 ;
        RECT 1829.510 959.000 1829.790 959.280 ;
        RECT 1828.590 862.440 1828.870 862.720 ;
        RECT 1829.510 862.440 1829.790 862.720 ;
      LAYER met3 ;
        RECT 1828.565 959.290 1828.895 959.305 ;
        RECT 1829.485 959.290 1829.815 959.305 ;
        RECT 1828.565 958.990 1829.815 959.290 ;
        RECT 1828.565 958.975 1828.895 958.990 ;
        RECT 1829.485 958.975 1829.815 958.990 ;
        RECT 1828.565 862.730 1828.895 862.745 ;
        RECT 1829.485 862.730 1829.815 862.745 ;
        RECT 1828.565 862.430 1829.815 862.730 ;
        RECT 1828.565 862.415 1828.895 862.430 ;
        RECT 1829.485 862.415 1829.815 862.430 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1497.370 1669.640 1497.690 1669.700 ;
        RECT 1500.590 1669.640 1500.910 1669.700 ;
        RECT 1497.370 1669.500 1500.910 1669.640 ;
        RECT 1497.370 1669.440 1497.690 1669.500 ;
        RECT 1500.590 1669.440 1500.910 1669.500 ;
        RECT 686.390 27.440 686.710 27.500 ;
        RECT 1497.370 27.440 1497.690 27.500 ;
        RECT 686.390 27.300 1497.690 27.440 ;
        RECT 686.390 27.240 686.710 27.300 ;
        RECT 1497.370 27.240 1497.690 27.300 ;
      LAYER via ;
        RECT 1497.400 1669.440 1497.660 1669.700 ;
        RECT 1500.620 1669.440 1500.880 1669.700 ;
        RECT 686.420 27.240 686.680 27.500 ;
        RECT 1497.400 27.240 1497.660 27.500 ;
      LAYER met2 ;
        RECT 1501.920 1700.410 1502.200 1704.000 ;
        RECT 1500.680 1700.270 1502.200 1700.410 ;
        RECT 1500.680 1669.730 1500.820 1700.270 ;
        RECT 1501.920 1700.000 1502.200 1700.270 ;
        RECT 1497.400 1669.410 1497.660 1669.730 ;
        RECT 1500.620 1669.410 1500.880 1669.730 ;
        RECT 1497.460 27.530 1497.600 1669.410 ;
        RECT 686.420 27.210 686.680 27.530 ;
        RECT 1497.400 27.210 1497.660 27.530 ;
        RECT 686.480 2.400 686.620 27.210 ;
        RECT 686.270 -4.800 686.830 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1836.390 1642.440 1836.710 1642.500 ;
        RECT 1839.150 1642.440 1839.470 1642.500 ;
        RECT 1836.390 1642.300 1839.470 1642.440 ;
        RECT 1836.390 1642.240 1836.710 1642.300 ;
        RECT 1839.150 1642.240 1839.470 1642.300 ;
        RECT 1836.850 1545.880 1837.170 1545.940 ;
        RECT 1837.310 1545.880 1837.630 1545.940 ;
        RECT 1836.850 1545.740 1837.630 1545.880 ;
        RECT 1836.850 1545.680 1837.170 1545.740 ;
        RECT 1837.310 1545.680 1837.630 1545.740 ;
        RECT 1836.850 1463.060 1837.170 1463.320 ;
        RECT 1836.940 1462.640 1837.080 1463.060 ;
        RECT 1836.850 1462.380 1837.170 1462.640 ;
        RECT 1836.850 1366.500 1837.170 1366.760 ;
        RECT 1836.940 1366.080 1837.080 1366.500 ;
        RECT 1836.850 1365.820 1837.170 1366.080 ;
        RECT 1837.310 1173.240 1837.630 1173.300 ;
        RECT 1836.940 1173.100 1837.630 1173.240 ;
        RECT 1836.940 1172.960 1837.080 1173.100 ;
        RECT 1837.310 1173.040 1837.630 1173.100 ;
        RECT 1836.850 1172.700 1837.170 1172.960 ;
        RECT 1837.310 1076.680 1837.630 1076.740 ;
        RECT 1836.940 1076.540 1837.630 1076.680 ;
        RECT 1836.940 1076.400 1837.080 1076.540 ;
        RECT 1837.310 1076.480 1837.630 1076.540 ;
        RECT 1836.850 1076.140 1837.170 1076.400 ;
        RECT 1837.310 980.120 1837.630 980.180 ;
        RECT 1836.940 979.980 1837.630 980.120 ;
        RECT 1836.940 979.840 1837.080 979.980 ;
        RECT 1837.310 979.920 1837.630 979.980 ;
        RECT 1836.850 979.580 1837.170 979.840 ;
        RECT 1836.850 676.160 1837.170 676.220 ;
        RECT 1837.770 676.160 1838.090 676.220 ;
        RECT 1836.850 676.020 1838.090 676.160 ;
        RECT 1836.850 675.960 1837.170 676.020 ;
        RECT 1837.770 675.960 1838.090 676.020 ;
        RECT 1836.390 275.980 1836.710 276.040 ;
        RECT 1836.850 275.980 1837.170 276.040 ;
        RECT 1836.390 275.840 1837.170 275.980 ;
        RECT 1836.390 275.780 1836.710 275.840 ;
        RECT 1836.850 275.780 1837.170 275.840 ;
        RECT 1836.850 179.760 1837.170 179.820 ;
        RECT 1837.310 179.760 1837.630 179.820 ;
        RECT 1836.850 179.620 1837.630 179.760 ;
        RECT 1836.850 179.560 1837.170 179.620 ;
        RECT 1837.310 179.560 1837.630 179.620 ;
        RECT 1449.070 52.940 1449.390 53.000 ;
        RECT 1836.850 52.940 1837.170 53.000 ;
        RECT 1449.070 52.800 1837.170 52.940 ;
        RECT 1449.070 52.740 1449.390 52.800 ;
        RECT 1836.850 52.740 1837.170 52.800 ;
        RECT 1346.490 18.260 1346.810 18.320 ;
        RECT 1449.070 18.260 1449.390 18.320 ;
        RECT 1346.490 18.120 1449.390 18.260 ;
        RECT 1346.490 18.060 1346.810 18.120 ;
        RECT 1449.070 18.060 1449.390 18.120 ;
      LAYER via ;
        RECT 1836.420 1642.240 1836.680 1642.500 ;
        RECT 1839.180 1642.240 1839.440 1642.500 ;
        RECT 1836.880 1545.680 1837.140 1545.940 ;
        RECT 1837.340 1545.680 1837.600 1545.940 ;
        RECT 1836.880 1463.060 1837.140 1463.320 ;
        RECT 1836.880 1462.380 1837.140 1462.640 ;
        RECT 1836.880 1366.500 1837.140 1366.760 ;
        RECT 1836.880 1365.820 1837.140 1366.080 ;
        RECT 1837.340 1173.040 1837.600 1173.300 ;
        RECT 1836.880 1172.700 1837.140 1172.960 ;
        RECT 1837.340 1076.480 1837.600 1076.740 ;
        RECT 1836.880 1076.140 1837.140 1076.400 ;
        RECT 1837.340 979.920 1837.600 980.180 ;
        RECT 1836.880 979.580 1837.140 979.840 ;
        RECT 1836.880 675.960 1837.140 676.220 ;
        RECT 1837.800 675.960 1838.060 676.220 ;
        RECT 1836.420 275.780 1836.680 276.040 ;
        RECT 1836.880 275.780 1837.140 276.040 ;
        RECT 1836.880 179.560 1837.140 179.820 ;
        RECT 1837.340 179.560 1837.600 179.820 ;
        RECT 1449.100 52.740 1449.360 53.000 ;
        RECT 1836.880 52.740 1837.140 53.000 ;
        RECT 1346.520 18.060 1346.780 18.320 ;
        RECT 1449.100 18.060 1449.360 18.320 ;
      LAYER met2 ;
        RECT 1841.860 1701.090 1842.140 1704.000 ;
        RECT 1839.240 1700.950 1842.140 1701.090 ;
        RECT 1839.240 1642.530 1839.380 1700.950 ;
        RECT 1841.860 1700.000 1842.140 1700.950 ;
        RECT 1836.420 1642.210 1836.680 1642.530 ;
        RECT 1839.180 1642.210 1839.440 1642.530 ;
        RECT 1836.480 1641.930 1836.620 1642.210 ;
        RECT 1836.480 1641.790 1837.540 1641.930 ;
        RECT 1837.400 1545.970 1837.540 1641.790 ;
        RECT 1836.880 1545.650 1837.140 1545.970 ;
        RECT 1837.340 1545.650 1837.600 1545.970 ;
        RECT 1836.940 1463.350 1837.080 1545.650 ;
        RECT 1836.880 1463.030 1837.140 1463.350 ;
        RECT 1836.880 1462.350 1837.140 1462.670 ;
        RECT 1836.940 1366.790 1837.080 1462.350 ;
        RECT 1836.880 1366.470 1837.140 1366.790 ;
        RECT 1836.880 1365.790 1837.140 1366.110 ;
        RECT 1836.940 1269.970 1837.080 1365.790 ;
        RECT 1836.480 1269.830 1837.080 1269.970 ;
        RECT 1836.480 1269.290 1836.620 1269.830 ;
        RECT 1836.480 1269.150 1837.080 1269.290 ;
        RECT 1836.940 1207.410 1837.080 1269.150 ;
        RECT 1836.940 1207.270 1837.540 1207.410 ;
        RECT 1837.400 1173.330 1837.540 1207.270 ;
        RECT 1837.340 1173.010 1837.600 1173.330 ;
        RECT 1836.880 1172.670 1837.140 1172.990 ;
        RECT 1836.940 1110.850 1837.080 1172.670 ;
        RECT 1836.940 1110.710 1837.540 1110.850 ;
        RECT 1837.400 1076.770 1837.540 1110.710 ;
        RECT 1837.340 1076.450 1837.600 1076.770 ;
        RECT 1836.880 1076.110 1837.140 1076.430 ;
        RECT 1836.940 1014.290 1837.080 1076.110 ;
        RECT 1836.940 1014.150 1837.540 1014.290 ;
        RECT 1837.400 980.210 1837.540 1014.150 ;
        RECT 1837.340 979.890 1837.600 980.210 ;
        RECT 1836.880 979.550 1837.140 979.870 ;
        RECT 1836.940 677.125 1837.080 979.550 ;
        RECT 1836.870 676.755 1837.150 677.125 ;
        RECT 1836.870 676.075 1837.150 676.445 ;
        RECT 1836.880 675.930 1837.140 676.075 ;
        RECT 1837.800 675.930 1838.060 676.250 ;
        RECT 1837.860 628.165 1838.000 675.930 ;
        RECT 1836.870 627.795 1837.150 628.165 ;
        RECT 1837.790 627.795 1838.070 628.165 ;
        RECT 1836.940 497.490 1837.080 627.795 ;
        RECT 1836.480 497.350 1837.080 497.490 ;
        RECT 1836.480 496.810 1836.620 497.350 ;
        RECT 1836.480 496.670 1837.080 496.810 ;
        RECT 1836.940 400.420 1837.080 496.670 ;
        RECT 1836.940 400.280 1837.540 400.420 ;
        RECT 1837.400 399.740 1837.540 400.280 ;
        RECT 1836.940 399.600 1837.540 399.740 ;
        RECT 1836.940 277.285 1837.080 399.600 ;
        RECT 1836.870 276.915 1837.150 277.285 ;
        RECT 1836.410 276.235 1836.690 276.605 ;
        RECT 1836.480 276.070 1836.620 276.235 ;
        RECT 1836.420 275.750 1836.680 276.070 ;
        RECT 1836.880 275.750 1837.140 276.070 ;
        RECT 1836.940 228.325 1837.080 275.750 ;
        RECT 1836.870 227.955 1837.150 228.325 ;
        RECT 1837.330 227.275 1837.610 227.645 ;
        RECT 1837.400 179.850 1837.540 227.275 ;
        RECT 1836.880 179.530 1837.140 179.850 ;
        RECT 1837.340 179.530 1837.600 179.850 ;
        RECT 1836.940 159.530 1837.080 179.530 ;
        RECT 1836.940 159.390 1837.540 159.530 ;
        RECT 1837.400 155.450 1837.540 159.390 ;
        RECT 1836.480 155.310 1837.540 155.450 ;
        RECT 1836.480 130.970 1836.620 155.310 ;
        RECT 1836.480 130.830 1837.080 130.970 ;
        RECT 1836.940 53.030 1837.080 130.830 ;
        RECT 1449.100 52.710 1449.360 53.030 ;
        RECT 1836.880 52.710 1837.140 53.030 ;
        RECT 1449.160 18.350 1449.300 52.710 ;
        RECT 1346.520 18.030 1346.780 18.350 ;
        RECT 1449.100 18.030 1449.360 18.350 ;
        RECT 1346.580 2.400 1346.720 18.030 ;
        RECT 1346.370 -4.800 1346.930 2.400 ;
      LAYER via2 ;
        RECT 1836.870 676.800 1837.150 677.080 ;
        RECT 1836.870 676.120 1837.150 676.400 ;
        RECT 1836.870 627.840 1837.150 628.120 ;
        RECT 1837.790 627.840 1838.070 628.120 ;
        RECT 1836.870 276.960 1837.150 277.240 ;
        RECT 1836.410 276.280 1836.690 276.560 ;
        RECT 1836.870 228.000 1837.150 228.280 ;
        RECT 1837.330 227.320 1837.610 227.600 ;
      LAYER met3 ;
        RECT 1836.845 677.090 1837.175 677.105 ;
        RECT 1836.630 676.775 1837.175 677.090 ;
        RECT 1836.630 676.425 1836.930 676.775 ;
        RECT 1836.630 676.110 1837.175 676.425 ;
        RECT 1836.845 676.095 1837.175 676.110 ;
        RECT 1836.845 628.130 1837.175 628.145 ;
        RECT 1837.765 628.130 1838.095 628.145 ;
        RECT 1836.845 627.830 1838.095 628.130 ;
        RECT 1836.845 627.815 1837.175 627.830 ;
        RECT 1837.765 627.815 1838.095 627.830 ;
        RECT 1836.845 277.250 1837.175 277.265 ;
        RECT 1835.710 276.950 1837.175 277.250 ;
        RECT 1835.710 276.570 1836.010 276.950 ;
        RECT 1836.845 276.935 1837.175 276.950 ;
        RECT 1836.385 276.570 1836.715 276.585 ;
        RECT 1835.710 276.270 1836.715 276.570 ;
        RECT 1836.385 276.255 1836.715 276.270 ;
        RECT 1836.845 228.290 1837.175 228.305 ;
        RECT 1836.630 227.975 1837.175 228.290 ;
        RECT 1836.630 227.610 1836.930 227.975 ;
        RECT 1837.305 227.610 1837.635 227.625 ;
        RECT 1836.630 227.310 1837.635 227.610 ;
        RECT 1837.305 227.295 1837.635 227.310 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1582.930 29.820 1583.250 29.880 ;
        RECT 1849.270 29.820 1849.590 29.880 ;
        RECT 1582.930 29.680 1849.590 29.820 ;
        RECT 1582.930 29.620 1583.250 29.680 ;
        RECT 1849.270 29.620 1849.590 29.680 ;
        RECT 1364.430 18.940 1364.750 19.000 ;
        RECT 1582.930 18.940 1583.250 19.000 ;
        RECT 1364.430 18.800 1583.250 18.940 ;
        RECT 1364.430 18.740 1364.750 18.800 ;
        RECT 1582.930 18.740 1583.250 18.800 ;
      LAYER via ;
        RECT 1582.960 29.620 1583.220 29.880 ;
        RECT 1849.300 29.620 1849.560 29.880 ;
        RECT 1364.460 18.740 1364.720 19.000 ;
        RECT 1582.960 18.740 1583.220 19.000 ;
      LAYER met2 ;
        RECT 1851.060 1700.410 1851.340 1704.000 ;
        RECT 1849.360 1700.270 1851.340 1700.410 ;
        RECT 1849.360 29.910 1849.500 1700.270 ;
        RECT 1851.060 1700.000 1851.340 1700.270 ;
        RECT 1582.960 29.590 1583.220 29.910 ;
        RECT 1849.300 29.590 1849.560 29.910 ;
        RECT 1583.020 19.030 1583.160 29.590 ;
        RECT 1364.460 18.710 1364.720 19.030 ;
        RECT 1582.960 18.710 1583.220 19.030 ;
        RECT 1364.520 2.400 1364.660 18.710 ;
        RECT 1364.310 -4.800 1364.870 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1856.705 1545.385 1856.875 1587.035 ;
        RECT 1856.245 30.345 1856.415 48.195 ;
      LAYER mcon ;
        RECT 1856.705 1586.865 1856.875 1587.035 ;
        RECT 1856.245 48.025 1856.415 48.195 ;
      LAYER met1 ;
        RECT 1857.550 1642.780 1857.870 1642.840 ;
        RECT 1856.720 1642.640 1857.870 1642.780 ;
        RECT 1856.720 1642.500 1856.860 1642.640 ;
        RECT 1857.550 1642.580 1857.870 1642.640 ;
        RECT 1856.630 1642.240 1856.950 1642.500 ;
        RECT 1856.630 1593.820 1856.950 1593.880 ;
        RECT 1857.090 1593.820 1857.410 1593.880 ;
        RECT 1856.630 1593.680 1857.410 1593.820 ;
        RECT 1856.630 1593.620 1856.950 1593.680 ;
        RECT 1857.090 1593.620 1857.410 1593.680 ;
        RECT 1856.630 1587.020 1856.950 1587.080 ;
        RECT 1856.435 1586.880 1856.950 1587.020 ;
        RECT 1856.630 1586.820 1856.950 1586.880 ;
        RECT 1856.630 1545.540 1856.950 1545.600 ;
        RECT 1856.435 1545.400 1856.950 1545.540 ;
        RECT 1856.630 1545.340 1856.950 1545.400 ;
        RECT 1857.090 1400.700 1857.410 1400.760 ;
        RECT 1857.550 1400.700 1857.870 1400.760 ;
        RECT 1857.090 1400.560 1857.870 1400.700 ;
        RECT 1857.090 1400.500 1857.410 1400.560 ;
        RECT 1857.550 1400.500 1857.870 1400.560 ;
        RECT 1857.090 627.880 1857.410 627.940 ;
        RECT 1857.550 627.880 1857.870 627.940 ;
        RECT 1857.090 627.740 1857.870 627.880 ;
        RECT 1857.090 627.680 1857.410 627.740 ;
        RECT 1857.550 627.680 1857.870 627.740 ;
        RECT 1856.170 144.740 1856.490 144.800 ;
        RECT 1857.090 144.740 1857.410 144.800 ;
        RECT 1856.170 144.600 1857.410 144.740 ;
        RECT 1856.170 144.540 1856.490 144.600 ;
        RECT 1857.090 144.540 1857.410 144.600 ;
        RECT 1856.170 48.180 1856.490 48.240 ;
        RECT 1855.975 48.040 1856.490 48.180 ;
        RECT 1856.170 47.980 1856.490 48.040 ;
        RECT 1573.270 30.500 1573.590 30.560 ;
        RECT 1856.185 30.500 1856.475 30.545 ;
        RECT 1573.270 30.360 1856.475 30.500 ;
        RECT 1573.270 30.300 1573.590 30.360 ;
        RECT 1856.185 30.315 1856.475 30.360 ;
        RECT 1573.270 20.980 1573.590 21.040 ;
        RECT 1572.440 20.840 1573.590 20.980 ;
        RECT 1382.370 20.640 1382.690 20.700 ;
        RECT 1572.440 20.640 1572.580 20.840 ;
        RECT 1573.270 20.780 1573.590 20.840 ;
        RECT 1382.370 20.500 1572.580 20.640 ;
        RECT 1382.370 20.440 1382.690 20.500 ;
      LAYER via ;
        RECT 1857.580 1642.580 1857.840 1642.840 ;
        RECT 1856.660 1642.240 1856.920 1642.500 ;
        RECT 1856.660 1593.620 1856.920 1593.880 ;
        RECT 1857.120 1593.620 1857.380 1593.880 ;
        RECT 1856.660 1586.820 1856.920 1587.080 ;
        RECT 1856.660 1545.340 1856.920 1545.600 ;
        RECT 1857.120 1400.500 1857.380 1400.760 ;
        RECT 1857.580 1400.500 1857.840 1400.760 ;
        RECT 1857.120 627.680 1857.380 627.940 ;
        RECT 1857.580 627.680 1857.840 627.940 ;
        RECT 1856.200 144.540 1856.460 144.800 ;
        RECT 1857.120 144.540 1857.380 144.800 ;
        RECT 1856.200 47.980 1856.460 48.240 ;
        RECT 1573.300 30.300 1573.560 30.560 ;
        RECT 1382.400 20.440 1382.660 20.700 ;
        RECT 1573.300 20.780 1573.560 21.040 ;
      LAYER met2 ;
        RECT 1859.800 1701.090 1860.080 1704.000 ;
        RECT 1857.640 1700.950 1860.080 1701.090 ;
        RECT 1857.640 1642.870 1857.780 1700.950 ;
        RECT 1859.800 1700.000 1860.080 1700.950 ;
        RECT 1857.580 1642.550 1857.840 1642.870 ;
        RECT 1856.660 1642.210 1856.920 1642.530 ;
        RECT 1856.720 1618.130 1856.860 1642.210 ;
        RECT 1856.720 1617.990 1857.320 1618.130 ;
        RECT 1857.180 1593.910 1857.320 1617.990 ;
        RECT 1856.660 1593.590 1856.920 1593.910 ;
        RECT 1857.120 1593.590 1857.380 1593.910 ;
        RECT 1856.720 1587.110 1856.860 1593.590 ;
        RECT 1856.660 1586.790 1856.920 1587.110 ;
        RECT 1856.660 1545.310 1856.920 1545.630 ;
        RECT 1856.720 1521.570 1856.860 1545.310 ;
        RECT 1856.720 1521.430 1857.320 1521.570 ;
        RECT 1857.180 1462.410 1857.320 1521.430 ;
        RECT 1856.720 1462.270 1857.320 1462.410 ;
        RECT 1856.720 1461.050 1856.860 1462.270 ;
        RECT 1856.720 1460.910 1857.320 1461.050 ;
        RECT 1857.180 1400.790 1857.320 1460.910 ;
        RECT 1857.120 1400.470 1857.380 1400.790 ;
        RECT 1857.580 1400.470 1857.840 1400.790 ;
        RECT 1857.640 1365.850 1857.780 1400.470 ;
        RECT 1857.180 1365.710 1857.780 1365.850 ;
        RECT 1857.180 1269.970 1857.320 1365.710 ;
        RECT 1856.720 1269.830 1857.320 1269.970 ;
        RECT 1856.720 1269.290 1856.860 1269.830 ;
        RECT 1856.720 1269.150 1857.320 1269.290 ;
        RECT 1857.180 883.050 1857.320 1269.150 ;
        RECT 1856.720 882.910 1857.320 883.050 ;
        RECT 1856.720 881.690 1856.860 882.910 ;
        RECT 1856.720 881.550 1857.320 881.690 ;
        RECT 1857.180 786.490 1857.320 881.550 ;
        RECT 1856.720 786.350 1857.320 786.490 ;
        RECT 1856.720 785.130 1856.860 786.350 ;
        RECT 1856.720 784.990 1857.320 785.130 ;
        RECT 1857.180 690.610 1857.320 784.990 ;
        RECT 1856.720 690.470 1857.320 690.610 ;
        RECT 1856.720 688.570 1856.860 690.470 ;
        RECT 1856.720 688.430 1857.320 688.570 ;
        RECT 1857.180 627.970 1857.320 688.430 ;
        RECT 1857.120 627.650 1857.380 627.970 ;
        RECT 1857.580 627.650 1857.840 627.970 ;
        RECT 1857.640 593.370 1857.780 627.650 ;
        RECT 1857.180 593.230 1857.780 593.370 ;
        RECT 1857.180 497.490 1857.320 593.230 ;
        RECT 1856.720 497.350 1857.320 497.490 ;
        RECT 1856.720 496.810 1856.860 497.350 ;
        RECT 1856.720 496.670 1857.320 496.810 ;
        RECT 1857.180 303.690 1857.320 496.670 ;
        RECT 1856.720 303.550 1857.320 303.690 ;
        RECT 1856.720 303.010 1856.860 303.550 ;
        RECT 1856.720 302.870 1857.320 303.010 ;
        RECT 1857.180 235.010 1857.320 302.870 ;
        RECT 1856.720 234.870 1857.320 235.010 ;
        RECT 1856.720 203.730 1856.860 234.870 ;
        RECT 1856.720 203.590 1857.320 203.730 ;
        RECT 1857.180 144.830 1857.320 203.590 ;
        RECT 1856.200 144.510 1856.460 144.830 ;
        RECT 1857.120 144.510 1857.380 144.830 ;
        RECT 1856.260 96.970 1856.400 144.510 ;
        RECT 1856.260 96.830 1856.860 96.970 ;
        RECT 1856.720 62.290 1856.860 96.830 ;
        RECT 1856.720 62.150 1857.320 62.290 ;
        RECT 1857.180 48.690 1857.320 62.150 ;
        RECT 1856.260 48.550 1857.320 48.690 ;
        RECT 1856.260 48.270 1856.400 48.550 ;
        RECT 1856.200 47.950 1856.460 48.270 ;
        RECT 1573.300 30.270 1573.560 30.590 ;
        RECT 1573.360 21.070 1573.500 30.270 ;
        RECT 1573.300 20.750 1573.560 21.070 ;
        RECT 1382.400 20.410 1382.660 20.730 ;
        RECT 1382.460 2.400 1382.600 20.410 ;
        RECT 1382.250 -4.800 1382.810 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1399.850 30.840 1400.170 30.900 ;
        RECT 1863.990 30.840 1864.310 30.900 ;
        RECT 1399.850 30.700 1864.310 30.840 ;
        RECT 1399.850 30.640 1400.170 30.700 ;
        RECT 1863.990 30.640 1864.310 30.700 ;
      LAYER via ;
        RECT 1399.880 30.640 1400.140 30.900 ;
        RECT 1864.020 30.640 1864.280 30.900 ;
      LAYER met2 ;
        RECT 1869.000 1700.410 1869.280 1704.000 ;
        RECT 1867.300 1700.270 1869.280 1700.410 ;
        RECT 1867.300 1656.210 1867.440 1700.270 ;
        RECT 1869.000 1700.000 1869.280 1700.270 ;
        RECT 1864.080 1656.070 1867.440 1656.210 ;
        RECT 1864.080 30.930 1864.220 1656.070 ;
        RECT 1399.880 30.610 1400.140 30.930 ;
        RECT 1864.020 30.610 1864.280 30.930 ;
        RECT 1399.940 15.370 1400.080 30.610 ;
        RECT 1399.940 15.230 1400.540 15.370 ;
        RECT 1400.400 2.400 1400.540 15.230 ;
        RECT 1400.190 -4.800 1400.750 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1418.250 31.180 1418.570 31.240 ;
        RECT 1876.870 31.180 1877.190 31.240 ;
        RECT 1418.250 31.040 1877.190 31.180 ;
        RECT 1418.250 30.980 1418.570 31.040 ;
        RECT 1876.870 30.980 1877.190 31.040 ;
      LAYER via ;
        RECT 1418.280 30.980 1418.540 31.240 ;
        RECT 1876.900 30.980 1877.160 31.240 ;
      LAYER met2 ;
        RECT 1878.200 1700.410 1878.480 1704.000 ;
        RECT 1876.960 1700.270 1878.480 1700.410 ;
        RECT 1876.960 31.270 1877.100 1700.270 ;
        RECT 1878.200 1700.000 1878.480 1700.270 ;
        RECT 1418.280 30.950 1418.540 31.270 ;
        RECT 1876.900 30.950 1877.160 31.270 ;
        RECT 1418.340 2.400 1418.480 30.950 ;
        RECT 1418.130 -4.800 1418.690 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1885.225 1635.485 1885.395 1678.155 ;
        RECT 1884.765 1538.925 1884.935 1587.035 ;
        RECT 1884.765 1449.165 1884.935 1497.275 ;
        RECT 1884.765 772.905 1884.935 821.015 ;
        RECT 1884.305 31.365 1884.475 49.895 ;
      LAYER mcon ;
        RECT 1885.225 1677.985 1885.395 1678.155 ;
        RECT 1884.765 1586.865 1884.935 1587.035 ;
        RECT 1884.765 1497.105 1884.935 1497.275 ;
        RECT 1884.765 820.845 1884.935 821.015 ;
        RECT 1884.305 49.725 1884.475 49.895 ;
      LAYER met1 ;
        RECT 1885.150 1678.140 1885.470 1678.200 ;
        RECT 1884.955 1678.000 1885.470 1678.140 ;
        RECT 1885.150 1677.940 1885.470 1678.000 ;
        RECT 1885.150 1635.640 1885.470 1635.700 ;
        RECT 1884.955 1635.500 1885.470 1635.640 ;
        RECT 1885.150 1635.440 1885.470 1635.500 ;
        RECT 1884.690 1594.160 1885.010 1594.220 ;
        RECT 1885.150 1594.160 1885.470 1594.220 ;
        RECT 1884.690 1594.020 1885.470 1594.160 ;
        RECT 1884.690 1593.960 1885.010 1594.020 ;
        RECT 1885.150 1593.960 1885.470 1594.020 ;
        RECT 1884.690 1587.020 1885.010 1587.080 ;
        RECT 1884.495 1586.880 1885.010 1587.020 ;
        RECT 1884.690 1586.820 1885.010 1586.880 ;
        RECT 1884.690 1539.080 1885.010 1539.140 ;
        RECT 1884.495 1538.940 1885.010 1539.080 ;
        RECT 1884.690 1538.880 1885.010 1538.940 ;
        RECT 1884.690 1497.260 1885.010 1497.320 ;
        RECT 1884.495 1497.120 1885.010 1497.260 ;
        RECT 1884.690 1497.060 1885.010 1497.120 ;
        RECT 1884.690 1449.320 1885.010 1449.380 ;
        RECT 1884.495 1449.180 1885.010 1449.320 ;
        RECT 1884.690 1449.120 1885.010 1449.180 ;
        RECT 1884.690 1365.820 1885.010 1366.080 ;
        RECT 1884.780 1365.400 1884.920 1365.820 ;
        RECT 1884.690 1365.140 1885.010 1365.400 ;
        RECT 1884.690 1269.260 1885.010 1269.520 ;
        RECT 1884.780 1268.840 1884.920 1269.260 ;
        RECT 1884.690 1268.580 1885.010 1268.840 ;
        RECT 1884.690 1172.700 1885.010 1172.960 ;
        RECT 1884.780 1172.280 1884.920 1172.700 ;
        RECT 1884.690 1172.020 1885.010 1172.280 ;
        RECT 1884.690 1076.140 1885.010 1076.400 ;
        RECT 1884.780 1075.720 1884.920 1076.140 ;
        RECT 1884.690 1075.460 1885.010 1075.720 ;
        RECT 1884.690 979.580 1885.010 979.840 ;
        RECT 1884.780 979.160 1884.920 979.580 ;
        RECT 1884.690 978.900 1885.010 979.160 ;
        RECT 1884.690 845.480 1885.010 845.540 ;
        RECT 1885.610 845.480 1885.930 845.540 ;
        RECT 1884.690 845.340 1885.930 845.480 ;
        RECT 1884.690 845.280 1885.010 845.340 ;
        RECT 1885.610 845.280 1885.930 845.340 ;
        RECT 1884.690 821.000 1885.010 821.060 ;
        RECT 1884.495 820.860 1885.010 821.000 ;
        RECT 1884.690 820.800 1885.010 820.860 ;
        RECT 1884.690 773.060 1885.010 773.120 ;
        RECT 1884.495 772.920 1885.010 773.060 ;
        RECT 1884.690 772.860 1885.010 772.920 ;
        RECT 1884.690 689.900 1885.010 690.160 ;
        RECT 1884.780 689.480 1884.920 689.900 ;
        RECT 1884.690 689.220 1885.010 689.480 ;
        RECT 1884.690 400.220 1885.010 400.480 ;
        RECT 1884.780 399.800 1884.920 400.220 ;
        RECT 1884.690 399.540 1885.010 399.800 ;
        RECT 1884.690 338.540 1885.010 338.600 ;
        RECT 1884.320 338.400 1885.010 338.540 ;
        RECT 1884.320 338.260 1884.460 338.400 ;
        RECT 1884.690 338.340 1885.010 338.400 ;
        RECT 1884.230 338.000 1884.550 338.260 ;
        RECT 1884.230 193.360 1884.550 193.420 ;
        RECT 1884.690 193.360 1885.010 193.420 ;
        RECT 1884.230 193.220 1885.010 193.360 ;
        RECT 1884.230 193.160 1884.550 193.220 ;
        RECT 1884.690 193.160 1885.010 193.220 ;
        RECT 1884.230 137.940 1884.550 138.000 ;
        RECT 1885.150 137.940 1885.470 138.000 ;
        RECT 1884.230 137.800 1885.470 137.940 ;
        RECT 1884.230 137.740 1884.550 137.800 ;
        RECT 1885.150 137.740 1885.470 137.800 ;
        RECT 1884.245 49.880 1884.535 49.925 ;
        RECT 1885.150 49.880 1885.470 49.940 ;
        RECT 1884.245 49.740 1885.470 49.880 ;
        RECT 1884.245 49.695 1884.535 49.740 ;
        RECT 1885.150 49.680 1885.470 49.740 ;
        RECT 1435.730 31.520 1436.050 31.580 ;
        RECT 1884.245 31.520 1884.535 31.565 ;
        RECT 1435.730 31.380 1884.535 31.520 ;
        RECT 1435.730 31.320 1436.050 31.380 ;
        RECT 1884.245 31.335 1884.535 31.380 ;
      LAYER via ;
        RECT 1885.180 1677.940 1885.440 1678.200 ;
        RECT 1885.180 1635.440 1885.440 1635.700 ;
        RECT 1884.720 1593.960 1884.980 1594.220 ;
        RECT 1885.180 1593.960 1885.440 1594.220 ;
        RECT 1884.720 1586.820 1884.980 1587.080 ;
        RECT 1884.720 1538.880 1884.980 1539.140 ;
        RECT 1884.720 1497.060 1884.980 1497.320 ;
        RECT 1884.720 1449.120 1884.980 1449.380 ;
        RECT 1884.720 1365.820 1884.980 1366.080 ;
        RECT 1884.720 1365.140 1884.980 1365.400 ;
        RECT 1884.720 1269.260 1884.980 1269.520 ;
        RECT 1884.720 1268.580 1884.980 1268.840 ;
        RECT 1884.720 1172.700 1884.980 1172.960 ;
        RECT 1884.720 1172.020 1884.980 1172.280 ;
        RECT 1884.720 1076.140 1884.980 1076.400 ;
        RECT 1884.720 1075.460 1884.980 1075.720 ;
        RECT 1884.720 979.580 1884.980 979.840 ;
        RECT 1884.720 978.900 1884.980 979.160 ;
        RECT 1884.720 845.280 1884.980 845.540 ;
        RECT 1885.640 845.280 1885.900 845.540 ;
        RECT 1884.720 820.800 1884.980 821.060 ;
        RECT 1884.720 772.860 1884.980 773.120 ;
        RECT 1884.720 689.900 1884.980 690.160 ;
        RECT 1884.720 689.220 1884.980 689.480 ;
        RECT 1884.720 400.220 1884.980 400.480 ;
        RECT 1884.720 399.540 1884.980 399.800 ;
        RECT 1884.720 338.340 1884.980 338.600 ;
        RECT 1884.260 338.000 1884.520 338.260 ;
        RECT 1884.260 193.160 1884.520 193.420 ;
        RECT 1884.720 193.160 1884.980 193.420 ;
        RECT 1884.260 137.740 1884.520 138.000 ;
        RECT 1885.180 137.740 1885.440 138.000 ;
        RECT 1885.180 49.680 1885.440 49.940 ;
        RECT 1435.760 31.320 1436.020 31.580 ;
      LAYER met2 ;
        RECT 1887.400 1701.090 1887.680 1704.000 ;
        RECT 1885.240 1700.950 1887.680 1701.090 ;
        RECT 1885.240 1678.230 1885.380 1700.950 ;
        RECT 1887.400 1700.000 1887.680 1700.950 ;
        RECT 1885.180 1677.910 1885.440 1678.230 ;
        RECT 1885.180 1635.410 1885.440 1635.730 ;
        RECT 1885.240 1594.250 1885.380 1635.410 ;
        RECT 1884.720 1593.930 1884.980 1594.250 ;
        RECT 1885.180 1593.930 1885.440 1594.250 ;
        RECT 1884.780 1587.110 1884.920 1593.930 ;
        RECT 1884.720 1586.790 1884.980 1587.110 ;
        RECT 1884.720 1538.850 1884.980 1539.170 ;
        RECT 1884.780 1497.350 1884.920 1538.850 ;
        RECT 1884.720 1497.030 1884.980 1497.350 ;
        RECT 1884.720 1449.090 1884.980 1449.410 ;
        RECT 1884.780 1366.110 1884.920 1449.090 ;
        RECT 1884.720 1365.790 1884.980 1366.110 ;
        RECT 1884.720 1365.110 1884.980 1365.430 ;
        RECT 1884.780 1269.550 1884.920 1365.110 ;
        RECT 1884.720 1269.230 1884.980 1269.550 ;
        RECT 1884.720 1268.550 1884.980 1268.870 ;
        RECT 1884.780 1172.990 1884.920 1268.550 ;
        RECT 1884.720 1172.670 1884.980 1172.990 ;
        RECT 1884.720 1171.990 1884.980 1172.310 ;
        RECT 1884.780 1076.430 1884.920 1171.990 ;
        RECT 1884.720 1076.110 1884.980 1076.430 ;
        RECT 1884.720 1075.430 1884.980 1075.750 ;
        RECT 1884.780 979.870 1884.920 1075.430 ;
        RECT 1884.720 979.550 1884.980 979.870 ;
        RECT 1884.720 978.870 1884.980 979.190 ;
        RECT 1884.780 845.570 1884.920 978.870 ;
        RECT 1884.720 845.250 1884.980 845.570 ;
        RECT 1885.640 845.250 1885.900 845.570 ;
        RECT 1885.700 821.285 1885.840 845.250 ;
        RECT 1884.710 820.915 1884.990 821.285 ;
        RECT 1885.630 820.915 1885.910 821.285 ;
        RECT 1884.720 820.770 1884.980 820.915 ;
        RECT 1884.720 772.830 1884.980 773.150 ;
        RECT 1884.780 690.190 1884.920 772.830 ;
        RECT 1884.720 689.870 1884.980 690.190 ;
        RECT 1884.720 689.190 1884.980 689.510 ;
        RECT 1884.780 497.490 1884.920 689.190 ;
        RECT 1884.320 497.350 1884.920 497.490 ;
        RECT 1884.320 496.810 1884.460 497.350 ;
        RECT 1884.320 496.670 1884.920 496.810 ;
        RECT 1884.780 400.510 1884.920 496.670 ;
        RECT 1884.720 400.190 1884.980 400.510 ;
        RECT 1884.720 399.510 1884.980 399.830 ;
        RECT 1884.780 338.630 1884.920 399.510 ;
        RECT 1884.720 338.310 1884.980 338.630 ;
        RECT 1884.260 337.970 1884.520 338.290 ;
        RECT 1884.320 193.450 1884.460 337.970 ;
        RECT 1884.260 193.130 1884.520 193.450 ;
        RECT 1884.720 193.130 1884.980 193.450 ;
        RECT 1884.780 145.250 1884.920 193.130 ;
        RECT 1884.320 145.110 1884.920 145.250 ;
        RECT 1884.320 138.030 1884.460 145.110 ;
        RECT 1884.260 137.710 1884.520 138.030 ;
        RECT 1885.180 137.710 1885.440 138.030 ;
        RECT 1885.240 49.970 1885.380 137.710 ;
        RECT 1885.180 49.650 1885.440 49.970 ;
        RECT 1435.760 31.290 1436.020 31.610 ;
        RECT 1435.820 2.400 1435.960 31.290 ;
        RECT 1435.610 -4.800 1436.170 2.400 ;
      LAYER via2 ;
        RECT 1884.710 820.960 1884.990 821.240 ;
        RECT 1885.630 820.960 1885.910 821.240 ;
      LAYER met3 ;
        RECT 1884.685 821.250 1885.015 821.265 ;
        RECT 1885.605 821.250 1885.935 821.265 ;
        RECT 1884.685 820.950 1885.935 821.250 ;
        RECT 1884.685 820.935 1885.015 820.950 ;
        RECT 1885.605 820.935 1885.935 820.950 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1891.130 1678.140 1891.450 1678.200 ;
        RECT 1895.270 1678.140 1895.590 1678.200 ;
        RECT 1891.130 1678.000 1895.590 1678.140 ;
        RECT 1891.130 1677.940 1891.450 1678.000 ;
        RECT 1895.270 1677.940 1895.590 1678.000 ;
        RECT 1453.670 31.860 1453.990 31.920 ;
        RECT 1891.130 31.860 1891.450 31.920 ;
        RECT 1453.670 31.720 1891.450 31.860 ;
        RECT 1453.670 31.660 1453.990 31.720 ;
        RECT 1891.130 31.660 1891.450 31.720 ;
      LAYER via ;
        RECT 1891.160 1677.940 1891.420 1678.200 ;
        RECT 1895.300 1677.940 1895.560 1678.200 ;
        RECT 1453.700 31.660 1453.960 31.920 ;
        RECT 1891.160 31.660 1891.420 31.920 ;
      LAYER met2 ;
        RECT 1896.600 1700.410 1896.880 1704.000 ;
        RECT 1895.360 1700.270 1896.880 1700.410 ;
        RECT 1895.360 1678.230 1895.500 1700.270 ;
        RECT 1896.600 1700.000 1896.880 1700.270 ;
        RECT 1891.160 1677.910 1891.420 1678.230 ;
        RECT 1895.300 1677.910 1895.560 1678.230 ;
        RECT 1891.220 31.950 1891.360 1677.910 ;
        RECT 1453.700 31.630 1453.960 31.950 ;
        RECT 1891.160 31.630 1891.420 31.950 ;
        RECT 1453.760 2.400 1453.900 31.630 ;
        RECT 1453.550 -4.800 1454.110 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1471.610 26.420 1471.930 26.480 ;
        RECT 1904.470 26.420 1904.790 26.480 ;
        RECT 1471.610 26.280 1904.790 26.420 ;
        RECT 1471.610 26.220 1471.930 26.280 ;
        RECT 1904.470 26.220 1904.790 26.280 ;
      LAYER via ;
        RECT 1471.640 26.220 1471.900 26.480 ;
        RECT 1904.500 26.220 1904.760 26.480 ;
      LAYER met2 ;
        RECT 1905.800 1700.410 1906.080 1704.000 ;
        RECT 1904.560 1700.270 1906.080 1700.410 ;
        RECT 1904.560 26.510 1904.700 1700.270 ;
        RECT 1905.800 1700.000 1906.080 1700.270 ;
        RECT 1471.640 26.190 1471.900 26.510 ;
        RECT 1904.500 26.190 1904.760 26.510 ;
        RECT 1471.700 2.400 1471.840 26.190 ;
        RECT 1471.490 -4.800 1472.050 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1912.365 1587.545 1912.535 1635.315 ;
        RECT 1912.365 1538.925 1912.535 1587.035 ;
        RECT 1912.365 1352.605 1912.535 1400.715 ;
        RECT 1912.365 1256.045 1912.535 1304.155 ;
        RECT 1912.365 772.905 1912.535 838.355 ;
        RECT 1912.365 379.525 1912.535 434.775 ;
        RECT 1911.905 241.485 1912.075 255.595 ;
        RECT 1911.905 26.605 1912.075 65.535 ;
      LAYER mcon ;
        RECT 1912.365 1635.145 1912.535 1635.315 ;
        RECT 1912.365 1586.865 1912.535 1587.035 ;
        RECT 1912.365 1400.545 1912.535 1400.715 ;
        RECT 1912.365 1303.985 1912.535 1304.155 ;
        RECT 1912.365 838.185 1912.535 838.355 ;
        RECT 1912.365 434.605 1912.535 434.775 ;
        RECT 1911.905 255.425 1912.075 255.595 ;
        RECT 1911.905 65.365 1912.075 65.535 ;
      LAYER met1 ;
        RECT 1913.210 1683.580 1913.530 1683.640 ;
        RECT 1912.380 1683.440 1913.530 1683.580 ;
        RECT 1912.380 1683.300 1912.520 1683.440 ;
        RECT 1913.210 1683.380 1913.530 1683.440 ;
        RECT 1912.290 1683.040 1912.610 1683.300 ;
        RECT 1912.290 1635.300 1912.610 1635.360 ;
        RECT 1912.095 1635.160 1912.610 1635.300 ;
        RECT 1912.290 1635.100 1912.610 1635.160 ;
        RECT 1912.290 1587.700 1912.610 1587.760 ;
        RECT 1912.095 1587.560 1912.610 1587.700 ;
        RECT 1912.290 1587.500 1912.610 1587.560 ;
        RECT 1912.290 1587.020 1912.610 1587.080 ;
        RECT 1912.095 1586.880 1912.610 1587.020 ;
        RECT 1912.290 1586.820 1912.610 1586.880 ;
        RECT 1912.290 1539.080 1912.610 1539.140 ;
        RECT 1912.095 1538.940 1912.610 1539.080 ;
        RECT 1912.290 1538.880 1912.610 1538.940 ;
        RECT 1912.290 1490.120 1912.610 1490.180 ;
        RECT 1912.750 1490.120 1913.070 1490.180 ;
        RECT 1912.290 1489.980 1913.070 1490.120 ;
        RECT 1912.290 1489.920 1912.610 1489.980 ;
        RECT 1912.750 1489.920 1913.070 1489.980 ;
        RECT 1912.290 1400.700 1912.610 1400.760 ;
        RECT 1912.095 1400.560 1912.610 1400.700 ;
        RECT 1912.290 1400.500 1912.610 1400.560 ;
        RECT 1912.290 1352.760 1912.610 1352.820 ;
        RECT 1912.095 1352.620 1912.610 1352.760 ;
        RECT 1912.290 1352.560 1912.610 1352.620 ;
        RECT 1912.290 1304.140 1912.610 1304.200 ;
        RECT 1912.095 1304.000 1912.610 1304.140 ;
        RECT 1912.290 1303.940 1912.610 1304.000 ;
        RECT 1912.290 1256.200 1912.610 1256.260 ;
        RECT 1912.095 1256.060 1912.610 1256.200 ;
        RECT 1912.290 1256.000 1912.610 1256.060 ;
        RECT 1911.370 1159.300 1911.690 1159.360 ;
        RECT 1912.290 1159.300 1912.610 1159.360 ;
        RECT 1911.370 1159.160 1912.610 1159.300 ;
        RECT 1911.370 1159.100 1911.690 1159.160 ;
        RECT 1912.290 1159.100 1912.610 1159.160 ;
        RECT 1911.370 1062.740 1911.690 1062.800 ;
        RECT 1912.290 1062.740 1912.610 1062.800 ;
        RECT 1911.370 1062.600 1912.610 1062.740 ;
        RECT 1911.370 1062.540 1911.690 1062.600 ;
        RECT 1912.290 1062.540 1912.610 1062.600 ;
        RECT 1911.370 966.180 1911.690 966.240 ;
        RECT 1912.290 966.180 1912.610 966.240 ;
        RECT 1911.370 966.040 1912.610 966.180 ;
        RECT 1911.370 965.980 1911.690 966.040 ;
        RECT 1912.290 965.980 1912.610 966.040 ;
        RECT 1912.290 918.040 1912.610 918.300 ;
        RECT 1912.380 917.620 1912.520 918.040 ;
        RECT 1912.290 917.360 1912.610 917.620 ;
        RECT 1911.370 838.340 1911.690 838.400 ;
        RECT 1912.305 838.340 1912.595 838.385 ;
        RECT 1911.370 838.200 1912.595 838.340 ;
        RECT 1911.370 838.140 1911.690 838.200 ;
        RECT 1912.305 838.155 1912.595 838.200 ;
        RECT 1912.290 773.060 1912.610 773.120 ;
        RECT 1912.095 772.920 1912.610 773.060 ;
        RECT 1912.290 772.860 1912.610 772.920 ;
        RECT 1912.290 689.900 1912.610 690.160 ;
        RECT 1912.380 689.480 1912.520 689.900 ;
        RECT 1912.290 689.220 1912.610 689.480 ;
        RECT 1912.290 434.760 1912.610 434.820 ;
        RECT 1912.095 434.620 1912.610 434.760 ;
        RECT 1912.290 434.560 1912.610 434.620 ;
        RECT 1912.290 379.680 1912.610 379.740 ;
        RECT 1912.095 379.540 1912.610 379.680 ;
        RECT 1912.290 379.480 1912.610 379.540 ;
        RECT 1911.845 255.580 1912.135 255.625 ;
        RECT 1912.290 255.580 1912.610 255.640 ;
        RECT 1911.845 255.440 1912.610 255.580 ;
        RECT 1911.845 255.395 1912.135 255.440 ;
        RECT 1912.290 255.380 1912.610 255.440 ;
        RECT 1911.830 241.640 1912.150 241.700 ;
        RECT 1911.635 241.500 1912.150 241.640 ;
        RECT 1911.830 241.440 1912.150 241.500 ;
        RECT 1911.830 193.360 1912.150 193.420 ;
        RECT 1912.290 193.360 1912.610 193.420 ;
        RECT 1911.830 193.220 1912.610 193.360 ;
        RECT 1911.830 193.160 1912.150 193.220 ;
        RECT 1912.290 193.160 1912.610 193.220 ;
        RECT 1911.830 137.940 1912.150 138.000 ;
        RECT 1913.210 137.940 1913.530 138.000 ;
        RECT 1911.830 137.800 1913.530 137.940 ;
        RECT 1911.830 137.740 1912.150 137.800 ;
        RECT 1913.210 137.740 1913.530 137.800 ;
        RECT 1911.845 65.520 1912.135 65.565 ;
        RECT 1913.210 65.520 1913.530 65.580 ;
        RECT 1911.845 65.380 1913.530 65.520 ;
        RECT 1911.845 65.335 1912.135 65.380 ;
        RECT 1913.210 65.320 1913.530 65.380 ;
        RECT 1489.550 26.760 1489.870 26.820 ;
        RECT 1911.845 26.760 1912.135 26.805 ;
        RECT 1489.550 26.620 1912.135 26.760 ;
        RECT 1489.550 26.560 1489.870 26.620 ;
        RECT 1911.845 26.575 1912.135 26.620 ;
      LAYER via ;
        RECT 1913.240 1683.380 1913.500 1683.640 ;
        RECT 1912.320 1683.040 1912.580 1683.300 ;
        RECT 1912.320 1635.100 1912.580 1635.360 ;
        RECT 1912.320 1587.500 1912.580 1587.760 ;
        RECT 1912.320 1586.820 1912.580 1587.080 ;
        RECT 1912.320 1538.880 1912.580 1539.140 ;
        RECT 1912.320 1489.920 1912.580 1490.180 ;
        RECT 1912.780 1489.920 1913.040 1490.180 ;
        RECT 1912.320 1400.500 1912.580 1400.760 ;
        RECT 1912.320 1352.560 1912.580 1352.820 ;
        RECT 1912.320 1303.940 1912.580 1304.200 ;
        RECT 1912.320 1256.000 1912.580 1256.260 ;
        RECT 1911.400 1159.100 1911.660 1159.360 ;
        RECT 1912.320 1159.100 1912.580 1159.360 ;
        RECT 1911.400 1062.540 1911.660 1062.800 ;
        RECT 1912.320 1062.540 1912.580 1062.800 ;
        RECT 1911.400 965.980 1911.660 966.240 ;
        RECT 1912.320 965.980 1912.580 966.240 ;
        RECT 1912.320 918.040 1912.580 918.300 ;
        RECT 1912.320 917.360 1912.580 917.620 ;
        RECT 1911.400 838.140 1911.660 838.400 ;
        RECT 1912.320 772.860 1912.580 773.120 ;
        RECT 1912.320 689.900 1912.580 690.160 ;
        RECT 1912.320 689.220 1912.580 689.480 ;
        RECT 1912.320 434.560 1912.580 434.820 ;
        RECT 1912.320 379.480 1912.580 379.740 ;
        RECT 1912.320 255.380 1912.580 255.640 ;
        RECT 1911.860 241.440 1912.120 241.700 ;
        RECT 1911.860 193.160 1912.120 193.420 ;
        RECT 1912.320 193.160 1912.580 193.420 ;
        RECT 1911.860 137.740 1912.120 138.000 ;
        RECT 1913.240 137.740 1913.500 138.000 ;
        RECT 1913.240 65.320 1913.500 65.580 ;
        RECT 1489.580 26.560 1489.840 26.820 ;
      LAYER met2 ;
        RECT 1915.000 1700.410 1915.280 1704.000 ;
        RECT 1913.300 1700.270 1915.280 1700.410 ;
        RECT 1913.300 1683.670 1913.440 1700.270 ;
        RECT 1915.000 1700.000 1915.280 1700.270 ;
        RECT 1913.240 1683.350 1913.500 1683.670 ;
        RECT 1912.320 1683.010 1912.580 1683.330 ;
        RECT 1912.380 1635.390 1912.520 1683.010 ;
        RECT 1912.320 1635.070 1912.580 1635.390 ;
        RECT 1912.320 1587.470 1912.580 1587.790 ;
        RECT 1912.380 1587.110 1912.520 1587.470 ;
        RECT 1912.320 1586.790 1912.580 1587.110 ;
        RECT 1912.320 1538.850 1912.580 1539.170 ;
        RECT 1912.380 1490.210 1912.520 1538.850 ;
        RECT 1912.320 1489.890 1912.580 1490.210 ;
        RECT 1912.780 1489.890 1913.040 1490.210 ;
        RECT 1912.840 1462.410 1912.980 1489.890 ;
        RECT 1912.380 1462.270 1912.980 1462.410 ;
        RECT 1912.380 1400.790 1912.520 1462.270 ;
        RECT 1912.320 1400.470 1912.580 1400.790 ;
        RECT 1912.320 1352.530 1912.580 1352.850 ;
        RECT 1912.380 1304.230 1912.520 1352.530 ;
        RECT 1912.320 1303.910 1912.580 1304.230 ;
        RECT 1912.320 1255.970 1912.580 1256.290 ;
        RECT 1912.380 1207.525 1912.520 1255.970 ;
        RECT 1911.390 1207.155 1911.670 1207.525 ;
        RECT 1912.310 1207.155 1912.590 1207.525 ;
        RECT 1911.460 1159.390 1911.600 1207.155 ;
        RECT 1911.400 1159.070 1911.660 1159.390 ;
        RECT 1912.320 1159.070 1912.580 1159.390 ;
        RECT 1912.380 1110.965 1912.520 1159.070 ;
        RECT 1911.390 1110.595 1911.670 1110.965 ;
        RECT 1912.310 1110.595 1912.590 1110.965 ;
        RECT 1911.460 1062.830 1911.600 1110.595 ;
        RECT 1911.400 1062.510 1911.660 1062.830 ;
        RECT 1912.320 1062.510 1912.580 1062.830 ;
        RECT 1912.380 1014.405 1912.520 1062.510 ;
        RECT 1911.390 1014.035 1911.670 1014.405 ;
        RECT 1912.310 1014.035 1912.590 1014.405 ;
        RECT 1911.460 966.270 1911.600 1014.035 ;
        RECT 1911.400 965.950 1911.660 966.270 ;
        RECT 1912.320 965.950 1912.580 966.270 ;
        RECT 1912.380 918.330 1912.520 965.950 ;
        RECT 1912.320 918.010 1912.580 918.330 ;
        RECT 1912.320 917.330 1912.580 917.650 ;
        RECT 1912.380 911.045 1912.520 917.330 ;
        RECT 1911.390 910.675 1911.670 911.045 ;
        RECT 1912.310 910.675 1912.590 911.045 ;
        RECT 1911.460 838.430 1911.600 910.675 ;
        RECT 1911.400 838.110 1911.660 838.430 ;
        RECT 1912.320 772.830 1912.580 773.150 ;
        RECT 1912.380 690.190 1912.520 772.830 ;
        RECT 1912.320 689.870 1912.580 690.190 ;
        RECT 1912.320 689.190 1912.580 689.510 ;
        RECT 1912.380 497.490 1912.520 689.190 ;
        RECT 1911.920 497.350 1912.520 497.490 ;
        RECT 1911.920 496.810 1912.060 497.350 ;
        RECT 1911.920 496.670 1912.520 496.810 ;
        RECT 1912.380 434.850 1912.520 496.670 ;
        RECT 1912.320 434.530 1912.580 434.850 ;
        RECT 1912.320 379.450 1912.580 379.770 ;
        RECT 1912.380 255.670 1912.520 379.450 ;
        RECT 1912.320 255.350 1912.580 255.670 ;
        RECT 1911.860 241.410 1912.120 241.730 ;
        RECT 1911.920 193.450 1912.060 241.410 ;
        RECT 1911.860 193.130 1912.120 193.450 ;
        RECT 1912.320 193.130 1912.580 193.450 ;
        RECT 1912.380 145.250 1912.520 193.130 ;
        RECT 1911.920 145.110 1912.520 145.250 ;
        RECT 1911.920 138.030 1912.060 145.110 ;
        RECT 1911.860 137.710 1912.120 138.030 ;
        RECT 1913.240 137.710 1913.500 138.030 ;
        RECT 1913.300 65.610 1913.440 137.710 ;
        RECT 1913.240 65.290 1913.500 65.610 ;
        RECT 1489.580 26.530 1489.840 26.850 ;
        RECT 1489.640 2.400 1489.780 26.530 ;
        RECT 1489.430 -4.800 1489.990 2.400 ;
      LAYER via2 ;
        RECT 1911.390 1207.200 1911.670 1207.480 ;
        RECT 1912.310 1207.200 1912.590 1207.480 ;
        RECT 1911.390 1110.640 1911.670 1110.920 ;
        RECT 1912.310 1110.640 1912.590 1110.920 ;
        RECT 1911.390 1014.080 1911.670 1014.360 ;
        RECT 1912.310 1014.080 1912.590 1014.360 ;
        RECT 1911.390 910.720 1911.670 911.000 ;
        RECT 1912.310 910.720 1912.590 911.000 ;
      LAYER met3 ;
        RECT 1911.365 1207.490 1911.695 1207.505 ;
        RECT 1912.285 1207.490 1912.615 1207.505 ;
        RECT 1911.365 1207.190 1912.615 1207.490 ;
        RECT 1911.365 1207.175 1911.695 1207.190 ;
        RECT 1912.285 1207.175 1912.615 1207.190 ;
        RECT 1911.365 1110.930 1911.695 1110.945 ;
        RECT 1912.285 1110.930 1912.615 1110.945 ;
        RECT 1911.365 1110.630 1912.615 1110.930 ;
        RECT 1911.365 1110.615 1911.695 1110.630 ;
        RECT 1912.285 1110.615 1912.615 1110.630 ;
        RECT 1911.365 1014.370 1911.695 1014.385 ;
        RECT 1912.285 1014.370 1912.615 1014.385 ;
        RECT 1911.365 1014.070 1912.615 1014.370 ;
        RECT 1911.365 1014.055 1911.695 1014.070 ;
        RECT 1912.285 1014.055 1912.615 1014.070 ;
        RECT 1911.365 911.010 1911.695 911.025 ;
        RECT 1912.285 911.010 1912.615 911.025 ;
        RECT 1911.365 910.710 1912.615 911.010 ;
        RECT 1911.365 910.695 1911.695 910.710 ;
        RECT 1912.285 910.695 1912.615 910.710 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1507.030 27.100 1507.350 27.160 ;
        RECT 1919.190 27.100 1919.510 27.160 ;
        RECT 1507.030 26.960 1919.510 27.100 ;
        RECT 1507.030 26.900 1507.350 26.960 ;
        RECT 1919.190 26.900 1919.510 26.960 ;
      LAYER via ;
        RECT 1507.060 26.900 1507.320 27.160 ;
        RECT 1919.220 26.900 1919.480 27.160 ;
      LAYER met2 ;
        RECT 1924.200 1700.410 1924.480 1704.000 ;
        RECT 1922.500 1700.270 1924.480 1700.410 ;
        RECT 1922.500 1656.210 1922.640 1700.270 ;
        RECT 1924.200 1700.000 1924.480 1700.270 ;
        RECT 1919.280 1656.070 1922.640 1656.210 ;
        RECT 1919.280 27.190 1919.420 1656.070 ;
        RECT 1507.060 26.870 1507.320 27.190 ;
        RECT 1919.220 26.870 1919.480 27.190 ;
        RECT 1507.120 2.400 1507.260 26.870 ;
        RECT 1506.910 -4.800 1507.470 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 710.310 59.740 710.630 59.800 ;
        RECT 1512.090 59.740 1512.410 59.800 ;
        RECT 710.310 59.600 1512.410 59.740 ;
        RECT 710.310 59.540 710.630 59.600 ;
        RECT 1512.090 59.540 1512.410 59.600 ;
        RECT 704.330 20.980 704.650 21.040 ;
        RECT 710.310 20.980 710.630 21.040 ;
        RECT 704.330 20.840 710.630 20.980 ;
        RECT 704.330 20.780 704.650 20.840 ;
        RECT 710.310 20.780 710.630 20.840 ;
      LAYER via ;
        RECT 710.340 59.540 710.600 59.800 ;
        RECT 1512.120 59.540 1512.380 59.800 ;
        RECT 704.360 20.780 704.620 21.040 ;
        RECT 710.340 20.780 710.600 21.040 ;
      LAYER met2 ;
        RECT 1511.120 1700.410 1511.400 1704.000 ;
        RECT 1511.120 1700.270 1512.320 1700.410 ;
        RECT 1511.120 1700.000 1511.400 1700.270 ;
        RECT 1512.180 59.830 1512.320 1700.270 ;
        RECT 710.340 59.510 710.600 59.830 ;
        RECT 1512.120 59.510 1512.380 59.830 ;
        RECT 710.400 21.070 710.540 59.510 ;
        RECT 704.360 20.750 704.620 21.070 ;
        RECT 710.340 20.750 710.600 21.070 ;
        RECT 704.420 2.400 704.560 20.750 ;
        RECT 704.210 -4.800 704.770 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1524.970 32.200 1525.290 32.260 ;
        RECT 1932.070 32.200 1932.390 32.260 ;
        RECT 1524.970 32.060 1932.390 32.200 ;
        RECT 1524.970 32.000 1525.290 32.060 ;
        RECT 1932.070 32.000 1932.390 32.060 ;
      LAYER via ;
        RECT 1525.000 32.000 1525.260 32.260 ;
        RECT 1932.100 32.000 1932.360 32.260 ;
      LAYER met2 ;
        RECT 1933.400 1700.410 1933.680 1704.000 ;
        RECT 1932.160 1700.270 1933.680 1700.410 ;
        RECT 1932.160 32.290 1932.300 1700.270 ;
        RECT 1933.400 1700.000 1933.680 1700.270 ;
        RECT 1525.000 31.970 1525.260 32.290 ;
        RECT 1932.100 31.970 1932.360 32.290 ;
        RECT 1525.060 2.400 1525.200 31.970 ;
        RECT 1524.850 -4.800 1525.410 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1939.890 1607.900 1940.210 1608.160 ;
        RECT 1939.980 1607.080 1940.120 1607.900 ;
        RECT 1940.350 1607.080 1940.670 1607.140 ;
        RECT 1939.980 1606.940 1940.670 1607.080 ;
        RECT 1940.350 1606.880 1940.670 1606.940 ;
        RECT 1939.890 1269.260 1940.210 1269.520 ;
        RECT 1939.980 1268.840 1940.120 1269.260 ;
        RECT 1939.890 1268.580 1940.210 1268.840 ;
        RECT 1939.890 1172.700 1940.210 1172.960 ;
        RECT 1939.980 1172.280 1940.120 1172.700 ;
        RECT 1939.890 1172.020 1940.210 1172.280 ;
        RECT 1939.890 1076.140 1940.210 1076.400 ;
        RECT 1939.980 1075.720 1940.120 1076.140 ;
        RECT 1939.890 1075.460 1940.210 1075.720 ;
        RECT 1939.890 979.580 1940.210 979.840 ;
        RECT 1939.980 979.160 1940.120 979.580 ;
        RECT 1939.890 978.900 1940.210 979.160 ;
        RECT 1939.890 787.140 1940.210 787.400 ;
        RECT 1939.980 786.720 1940.120 787.140 ;
        RECT 1939.890 786.460 1940.210 786.720 ;
        RECT 1939.890 400.220 1940.210 400.480 ;
        RECT 1939.980 399.800 1940.120 400.220 ;
        RECT 1939.890 399.540 1940.210 399.800 ;
        RECT 1939.430 289.580 1939.750 289.640 ;
        RECT 1939.890 289.580 1940.210 289.640 ;
        RECT 1939.430 289.440 1940.210 289.580 ;
        RECT 1939.430 289.380 1939.750 289.440 ;
        RECT 1939.890 289.380 1940.210 289.440 ;
        RECT 1939.430 145.080 1939.750 145.140 ;
        RECT 1940.350 145.080 1940.670 145.140 ;
        RECT 1939.430 144.940 1940.670 145.080 ;
        RECT 1939.430 144.880 1939.750 144.940 ;
        RECT 1940.350 144.880 1940.670 144.940 ;
        RECT 1542.910 32.540 1543.230 32.600 ;
        RECT 1939.430 32.540 1939.750 32.600 ;
        RECT 1542.910 32.400 1939.750 32.540 ;
        RECT 1542.910 32.340 1543.230 32.400 ;
        RECT 1939.430 32.340 1939.750 32.400 ;
      LAYER via ;
        RECT 1939.920 1607.900 1940.180 1608.160 ;
        RECT 1940.380 1606.880 1940.640 1607.140 ;
        RECT 1939.920 1269.260 1940.180 1269.520 ;
        RECT 1939.920 1268.580 1940.180 1268.840 ;
        RECT 1939.920 1172.700 1940.180 1172.960 ;
        RECT 1939.920 1172.020 1940.180 1172.280 ;
        RECT 1939.920 1076.140 1940.180 1076.400 ;
        RECT 1939.920 1075.460 1940.180 1075.720 ;
        RECT 1939.920 979.580 1940.180 979.840 ;
        RECT 1939.920 978.900 1940.180 979.160 ;
        RECT 1939.920 787.140 1940.180 787.400 ;
        RECT 1939.920 786.460 1940.180 786.720 ;
        RECT 1939.920 400.220 1940.180 400.480 ;
        RECT 1939.920 399.540 1940.180 399.800 ;
        RECT 1939.460 289.380 1939.720 289.640 ;
        RECT 1939.920 289.380 1940.180 289.640 ;
        RECT 1939.460 144.880 1939.720 145.140 ;
        RECT 1940.380 144.880 1940.640 145.140 ;
        RECT 1542.940 32.340 1543.200 32.600 ;
        RECT 1939.460 32.340 1939.720 32.600 ;
      LAYER met2 ;
        RECT 1942.600 1701.090 1942.880 1704.000 ;
        RECT 1940.440 1700.950 1942.880 1701.090 ;
        RECT 1940.440 1656.210 1940.580 1700.950 ;
        RECT 1942.600 1700.000 1942.880 1700.950 ;
        RECT 1939.980 1656.070 1940.580 1656.210 ;
        RECT 1939.980 1608.190 1940.120 1656.070 ;
        RECT 1939.920 1607.870 1940.180 1608.190 ;
        RECT 1940.380 1606.850 1940.640 1607.170 ;
        RECT 1940.440 1463.090 1940.580 1606.850 ;
        RECT 1939.520 1462.950 1940.580 1463.090 ;
        RECT 1939.520 1462.410 1939.660 1462.950 ;
        RECT 1939.520 1462.270 1940.120 1462.410 ;
        RECT 1939.980 1269.550 1940.120 1462.270 ;
        RECT 1939.920 1269.230 1940.180 1269.550 ;
        RECT 1939.920 1268.550 1940.180 1268.870 ;
        RECT 1939.980 1172.990 1940.120 1268.550 ;
        RECT 1939.920 1172.670 1940.180 1172.990 ;
        RECT 1939.920 1171.990 1940.180 1172.310 ;
        RECT 1939.980 1076.430 1940.120 1171.990 ;
        RECT 1939.920 1076.110 1940.180 1076.430 ;
        RECT 1939.920 1075.430 1940.180 1075.750 ;
        RECT 1939.980 979.870 1940.120 1075.430 ;
        RECT 1939.920 979.550 1940.180 979.870 ;
        RECT 1939.920 978.870 1940.180 979.190 ;
        RECT 1939.980 883.730 1940.120 978.870 ;
        RECT 1939.520 883.590 1940.120 883.730 ;
        RECT 1939.520 883.050 1939.660 883.590 ;
        RECT 1939.520 882.910 1940.120 883.050 ;
        RECT 1939.980 787.430 1940.120 882.910 ;
        RECT 1939.920 787.110 1940.180 787.430 ;
        RECT 1939.920 786.430 1940.180 786.750 ;
        RECT 1939.980 594.050 1940.120 786.430 ;
        RECT 1939.520 593.910 1940.120 594.050 ;
        RECT 1939.520 593.370 1939.660 593.910 ;
        RECT 1939.520 593.230 1940.120 593.370 ;
        RECT 1939.980 483.890 1940.120 593.230 ;
        RECT 1939.980 483.750 1940.580 483.890 ;
        RECT 1940.440 483.325 1940.580 483.750 ;
        RECT 1940.370 482.955 1940.650 483.325 ;
        RECT 1939.910 482.275 1940.190 482.645 ;
        RECT 1939.980 400.510 1940.120 482.275 ;
        RECT 1939.920 400.190 1940.180 400.510 ;
        RECT 1939.920 399.510 1940.180 399.830 ;
        RECT 1939.980 303.690 1940.120 399.510 ;
        RECT 1939.520 303.550 1940.120 303.690 ;
        RECT 1939.520 303.010 1939.660 303.550 ;
        RECT 1939.520 302.870 1940.120 303.010 ;
        RECT 1939.980 289.670 1940.120 302.870 ;
        RECT 1939.460 289.350 1939.720 289.670 ;
        RECT 1939.920 289.350 1940.180 289.670 ;
        RECT 1939.520 192.850 1939.660 289.350 ;
        RECT 1939.520 192.710 1940.580 192.850 ;
        RECT 1940.440 145.170 1940.580 192.710 ;
        RECT 1939.460 144.850 1939.720 145.170 ;
        RECT 1940.380 144.850 1940.640 145.170 ;
        RECT 1939.520 111.250 1939.660 144.850 ;
        RECT 1939.060 111.110 1939.660 111.250 ;
        RECT 1939.060 109.890 1939.200 111.110 ;
        RECT 1939.060 109.750 1939.660 109.890 ;
        RECT 1939.520 32.630 1939.660 109.750 ;
        RECT 1542.940 32.310 1543.200 32.630 ;
        RECT 1939.460 32.310 1939.720 32.630 ;
        RECT 1543.000 2.400 1543.140 32.310 ;
        RECT 1542.790 -4.800 1543.350 2.400 ;
      LAYER via2 ;
        RECT 1940.370 483.000 1940.650 483.280 ;
        RECT 1939.910 482.320 1940.190 482.600 ;
      LAYER met3 ;
        RECT 1940.345 483.290 1940.675 483.305 ;
        RECT 1940.345 482.975 1940.890 483.290 ;
        RECT 1939.885 482.610 1940.215 482.625 ;
        RECT 1940.590 482.610 1940.890 482.975 ;
        RECT 1939.885 482.310 1940.890 482.610 ;
        RECT 1939.885 482.295 1940.215 482.310 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1560.850 32.880 1561.170 32.940 ;
        RECT 1946.790 32.880 1947.110 32.940 ;
        RECT 1560.850 32.740 1947.110 32.880 ;
        RECT 1560.850 32.680 1561.170 32.740 ;
        RECT 1946.790 32.680 1947.110 32.740 ;
      LAYER via ;
        RECT 1560.880 32.680 1561.140 32.940 ;
        RECT 1946.820 32.680 1947.080 32.940 ;
      LAYER met2 ;
        RECT 1951.800 1700.410 1952.080 1704.000 ;
        RECT 1949.180 1700.270 1952.080 1700.410 ;
        RECT 1949.180 1678.650 1949.320 1700.270 ;
        RECT 1951.800 1700.000 1952.080 1700.270 ;
        RECT 1946.880 1678.510 1949.320 1678.650 ;
        RECT 1946.880 32.970 1947.020 1678.510 ;
        RECT 1560.880 32.650 1561.140 32.970 ;
        RECT 1946.820 32.650 1947.080 32.970 ;
        RECT 1560.940 2.400 1561.080 32.650 ;
        RECT 1560.730 -4.800 1561.290 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1578.790 27.440 1579.110 27.500 ;
        RECT 1959.670 27.440 1959.990 27.500 ;
        RECT 1578.790 27.300 1959.990 27.440 ;
        RECT 1578.790 27.240 1579.110 27.300 ;
        RECT 1959.670 27.240 1959.990 27.300 ;
      LAYER via ;
        RECT 1578.820 27.240 1579.080 27.500 ;
        RECT 1959.700 27.240 1959.960 27.500 ;
      LAYER met2 ;
        RECT 1961.000 1700.410 1961.280 1704.000 ;
        RECT 1959.760 1700.270 1961.280 1700.410 ;
        RECT 1959.760 27.530 1959.900 1700.270 ;
        RECT 1961.000 1700.000 1961.280 1700.270 ;
        RECT 1578.820 27.210 1579.080 27.530 ;
        RECT 1959.700 27.210 1959.960 27.530 ;
        RECT 1578.880 2.400 1579.020 27.210 ;
        RECT 1578.670 -4.800 1579.230 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1596.270 22.680 1596.590 22.740 ;
        RECT 1967.490 22.680 1967.810 22.740 ;
        RECT 1596.270 22.540 1967.810 22.680 ;
        RECT 1596.270 22.480 1596.590 22.540 ;
        RECT 1967.490 22.480 1967.810 22.540 ;
      LAYER via ;
        RECT 1596.300 22.480 1596.560 22.740 ;
        RECT 1967.520 22.480 1967.780 22.740 ;
      LAYER met2 ;
        RECT 1970.200 1700.410 1970.480 1704.000 ;
        RECT 1967.580 1700.270 1970.480 1700.410 ;
        RECT 1967.580 22.770 1967.720 1700.270 ;
        RECT 1970.200 1700.000 1970.480 1700.270 ;
        RECT 1596.300 22.450 1596.560 22.770 ;
        RECT 1967.520 22.450 1967.780 22.770 ;
        RECT 1596.360 2.400 1596.500 22.450 ;
        RECT 1596.150 -4.800 1596.710 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1614.210 22.340 1614.530 22.400 ;
        RECT 1974.390 22.340 1974.710 22.400 ;
        RECT 1614.210 22.200 1974.710 22.340 ;
        RECT 1614.210 22.140 1614.530 22.200 ;
        RECT 1974.390 22.140 1974.710 22.200 ;
      LAYER via ;
        RECT 1614.240 22.140 1614.500 22.400 ;
        RECT 1974.420 22.140 1974.680 22.400 ;
      LAYER met2 ;
        RECT 1979.400 1700.410 1979.680 1704.000 ;
        RECT 1976.780 1700.270 1979.680 1700.410 ;
        RECT 1976.780 1678.650 1976.920 1700.270 ;
        RECT 1979.400 1700.000 1979.680 1700.270 ;
        RECT 1974.480 1678.510 1976.920 1678.650 ;
        RECT 1974.480 22.430 1974.620 1678.510 ;
        RECT 1614.240 22.110 1614.500 22.430 ;
        RECT 1974.420 22.110 1974.680 22.430 ;
        RECT 1614.300 2.400 1614.440 22.110 ;
        RECT 1614.090 -4.800 1614.650 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1987.270 1400.840 1987.590 1401.100 ;
        RECT 1987.360 1400.420 1987.500 1400.840 ;
        RECT 1987.270 1400.160 1987.590 1400.420 ;
        RECT 1632.150 22.000 1632.470 22.060 ;
        RECT 1987.270 22.000 1987.590 22.060 ;
        RECT 1632.150 21.860 1987.590 22.000 ;
        RECT 1632.150 21.800 1632.470 21.860 ;
        RECT 1987.270 21.800 1987.590 21.860 ;
      LAYER via ;
        RECT 1987.300 1400.840 1987.560 1401.100 ;
        RECT 1987.300 1400.160 1987.560 1400.420 ;
        RECT 1632.180 21.800 1632.440 22.060 ;
        RECT 1987.300 21.800 1987.560 22.060 ;
      LAYER met2 ;
        RECT 1988.600 1700.410 1988.880 1704.000 ;
        RECT 1987.360 1700.270 1988.880 1700.410 ;
        RECT 1987.360 1401.130 1987.500 1700.270 ;
        RECT 1988.600 1700.000 1988.880 1700.270 ;
        RECT 1987.300 1400.810 1987.560 1401.130 ;
        RECT 1987.300 1400.130 1987.560 1400.450 ;
        RECT 1987.360 22.090 1987.500 1400.130 ;
        RECT 1632.180 21.770 1632.440 22.090 ;
        RECT 1987.300 21.770 1987.560 22.090 ;
        RECT 1632.240 2.400 1632.380 21.770 ;
        RECT 1632.030 -4.800 1632.590 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1650.090 21.660 1650.410 21.720 ;
        RECT 1995.090 21.660 1995.410 21.720 ;
        RECT 1650.090 21.520 1995.410 21.660 ;
        RECT 1650.090 21.460 1650.410 21.520 ;
        RECT 1995.090 21.460 1995.410 21.520 ;
      LAYER via ;
        RECT 1650.120 21.460 1650.380 21.720 ;
        RECT 1995.120 21.460 1995.380 21.720 ;
      LAYER met2 ;
        RECT 1997.800 1700.410 1998.080 1704.000 ;
        RECT 1995.180 1700.270 1998.080 1700.410 ;
        RECT 1995.180 21.750 1995.320 1700.270 ;
        RECT 1997.800 1700.000 1998.080 1700.270 ;
        RECT 1650.120 21.430 1650.380 21.750 ;
        RECT 1995.120 21.430 1995.380 21.750 ;
        RECT 1650.180 2.400 1650.320 21.430 ;
        RECT 1649.970 -4.800 1650.530 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2001.605 1594.005 2001.775 1635.315 ;
        RECT 2002.525 1497.105 2002.695 1579.895 ;
        RECT 2002.525 1304.325 2002.695 1352.435 ;
        RECT 2002.525 1207.425 2002.695 1255.875 ;
        RECT 2002.525 786.505 2002.695 821.015 ;
        RECT 2002.525 689.605 2002.695 724.455 ;
        RECT 2002.525 476.085 2002.695 524.195 ;
        RECT 2002.985 227.885 2003.155 235.875 ;
        RECT 2003.445 185.725 2003.615 227.375 ;
      LAYER mcon ;
        RECT 2001.605 1635.145 2001.775 1635.315 ;
        RECT 2002.525 1579.725 2002.695 1579.895 ;
        RECT 2002.525 1352.265 2002.695 1352.435 ;
        RECT 2002.525 1255.705 2002.695 1255.875 ;
        RECT 2002.525 820.845 2002.695 821.015 ;
        RECT 2002.525 724.285 2002.695 724.455 ;
        RECT 2002.525 524.025 2002.695 524.195 ;
        RECT 2002.985 235.705 2003.155 235.875 ;
        RECT 2003.445 227.205 2003.615 227.375 ;
      LAYER met1 ;
        RECT 2001.530 1642.100 2001.850 1642.160 ;
        RECT 2002.910 1642.100 2003.230 1642.160 ;
        RECT 2001.530 1641.960 2003.230 1642.100 ;
        RECT 2001.530 1641.900 2001.850 1641.960 ;
        RECT 2002.910 1641.900 2003.230 1641.960 ;
        RECT 2001.530 1635.300 2001.850 1635.360 ;
        RECT 2001.335 1635.160 2001.850 1635.300 ;
        RECT 2001.530 1635.100 2001.850 1635.160 ;
        RECT 2001.545 1594.160 2001.835 1594.205 ;
        RECT 2002.450 1594.160 2002.770 1594.220 ;
        RECT 2001.545 1594.020 2002.770 1594.160 ;
        RECT 2001.545 1593.975 2001.835 1594.020 ;
        RECT 2002.450 1593.960 2002.770 1594.020 ;
        RECT 2002.450 1579.880 2002.770 1579.940 ;
        RECT 2002.255 1579.740 2002.770 1579.880 ;
        RECT 2002.450 1579.680 2002.770 1579.740 ;
        RECT 2002.450 1497.260 2002.770 1497.320 ;
        RECT 2002.255 1497.120 2002.770 1497.260 ;
        RECT 2002.450 1497.060 2002.770 1497.120 ;
        RECT 2002.450 1414.100 2002.770 1414.360 ;
        RECT 2002.540 1413.680 2002.680 1414.100 ;
        RECT 2002.450 1413.420 2002.770 1413.680 ;
        RECT 2001.990 1366.020 2002.310 1366.080 ;
        RECT 2002.910 1366.020 2003.230 1366.080 ;
        RECT 2001.990 1365.880 2003.230 1366.020 ;
        RECT 2001.990 1365.820 2002.310 1365.880 ;
        RECT 2002.910 1365.820 2003.230 1365.880 ;
        RECT 2002.465 1352.420 2002.755 1352.465 ;
        RECT 2002.910 1352.420 2003.230 1352.480 ;
        RECT 2002.465 1352.280 2003.230 1352.420 ;
        RECT 2002.465 1352.235 2002.755 1352.280 ;
        RECT 2002.910 1352.220 2003.230 1352.280 ;
        RECT 2002.450 1304.480 2002.770 1304.540 ;
        RECT 2002.255 1304.340 2002.770 1304.480 ;
        RECT 2002.450 1304.280 2002.770 1304.340 ;
        RECT 2001.990 1269.460 2002.310 1269.520 ;
        RECT 2002.910 1269.460 2003.230 1269.520 ;
        RECT 2001.990 1269.320 2003.230 1269.460 ;
        RECT 2001.990 1269.260 2002.310 1269.320 ;
        RECT 2002.910 1269.260 2003.230 1269.320 ;
        RECT 2002.465 1255.860 2002.755 1255.905 ;
        RECT 2002.910 1255.860 2003.230 1255.920 ;
        RECT 2002.465 1255.720 2003.230 1255.860 ;
        RECT 2002.465 1255.675 2002.755 1255.720 ;
        RECT 2002.910 1255.660 2003.230 1255.720 ;
        RECT 2002.450 1207.580 2002.770 1207.640 ;
        RECT 2002.255 1207.440 2002.770 1207.580 ;
        RECT 2002.450 1207.380 2002.770 1207.440 ;
        RECT 2001.990 1172.900 2002.310 1172.960 ;
        RECT 2002.910 1172.900 2003.230 1172.960 ;
        RECT 2001.990 1172.760 2003.230 1172.900 ;
        RECT 2001.990 1172.700 2002.310 1172.760 ;
        RECT 2002.910 1172.700 2003.230 1172.760 ;
        RECT 2001.990 1111.020 2002.310 1111.080 ;
        RECT 2002.450 1111.020 2002.770 1111.080 ;
        RECT 2001.990 1110.880 2002.770 1111.020 ;
        RECT 2001.990 1110.820 2002.310 1110.880 ;
        RECT 2002.450 1110.820 2002.770 1110.880 ;
        RECT 2001.530 1062.740 2001.850 1062.800 ;
        RECT 2002.910 1062.740 2003.230 1062.800 ;
        RECT 2001.530 1062.600 2003.230 1062.740 ;
        RECT 2001.530 1062.540 2001.850 1062.600 ;
        RECT 2002.910 1062.540 2003.230 1062.600 ;
        RECT 2002.450 1014.120 2002.770 1014.180 ;
        RECT 2002.910 1014.120 2003.230 1014.180 ;
        RECT 2002.450 1013.980 2003.230 1014.120 ;
        RECT 2002.450 1013.920 2002.770 1013.980 ;
        RECT 2002.910 1013.920 2003.230 1013.980 ;
        RECT 2001.990 835.280 2002.310 835.340 ;
        RECT 2002.910 835.280 2003.230 835.340 ;
        RECT 2001.990 835.140 2003.230 835.280 ;
        RECT 2001.990 835.080 2002.310 835.140 ;
        RECT 2002.910 835.080 2003.230 835.140 ;
        RECT 2002.450 821.000 2002.770 821.060 ;
        RECT 2002.255 820.860 2002.770 821.000 ;
        RECT 2002.450 820.800 2002.770 820.860 ;
        RECT 2002.450 786.660 2002.770 786.720 ;
        RECT 2002.255 786.520 2002.770 786.660 ;
        RECT 2002.450 786.460 2002.770 786.520 ;
        RECT 2001.990 738.380 2002.310 738.440 ;
        RECT 2002.910 738.380 2003.230 738.440 ;
        RECT 2001.990 738.240 2003.230 738.380 ;
        RECT 2001.990 738.180 2002.310 738.240 ;
        RECT 2002.910 738.180 2003.230 738.240 ;
        RECT 2002.450 724.440 2002.770 724.500 ;
        RECT 2002.255 724.300 2002.770 724.440 ;
        RECT 2002.450 724.240 2002.770 724.300 ;
        RECT 2002.450 689.760 2002.770 689.820 ;
        RECT 2002.255 689.620 2002.770 689.760 ;
        RECT 2002.450 689.560 2002.770 689.620 ;
        RECT 2002.450 628.220 2002.770 628.280 ;
        RECT 2002.910 628.220 2003.230 628.280 ;
        RECT 2002.450 628.080 2003.230 628.220 ;
        RECT 2002.450 628.020 2002.770 628.080 ;
        RECT 2002.910 628.020 2003.230 628.080 ;
        RECT 2001.990 579.940 2002.310 580.000 ;
        RECT 2002.450 579.940 2002.770 580.000 ;
        RECT 2001.990 579.800 2002.770 579.940 ;
        RECT 2001.990 579.740 2002.310 579.800 ;
        RECT 2002.450 579.740 2002.770 579.800 ;
        RECT 2002.450 524.180 2002.770 524.240 ;
        RECT 2002.255 524.040 2002.770 524.180 ;
        RECT 2002.450 523.980 2002.770 524.040 ;
        RECT 2002.465 476.240 2002.755 476.285 ;
        RECT 2002.910 476.240 2003.230 476.300 ;
        RECT 2002.465 476.100 2003.230 476.240 ;
        RECT 2002.465 476.055 2002.755 476.100 ;
        RECT 2002.910 476.040 2003.230 476.100 ;
        RECT 2002.450 338.200 2002.770 338.260 ;
        RECT 2002.910 338.200 2003.230 338.260 ;
        RECT 2002.450 338.060 2003.230 338.200 ;
        RECT 2002.450 338.000 2002.770 338.060 ;
        RECT 2002.910 338.000 2003.230 338.060 ;
        RECT 2002.910 235.860 2003.230 235.920 ;
        RECT 2002.715 235.720 2003.230 235.860 ;
        RECT 2002.910 235.660 2003.230 235.720 ;
        RECT 2002.910 228.040 2003.230 228.100 ;
        RECT 2002.715 227.900 2003.230 228.040 ;
        RECT 2002.910 227.840 2003.230 227.900 ;
        RECT 2003.370 227.360 2003.690 227.420 ;
        RECT 2003.175 227.220 2003.690 227.360 ;
        RECT 2003.370 227.160 2003.690 227.220 ;
        RECT 2003.370 185.880 2003.690 185.940 ;
        RECT 2003.175 185.740 2003.690 185.880 ;
        RECT 2003.370 185.680 2003.690 185.740 ;
        RECT 2002.450 144.400 2002.770 144.460 ;
        RECT 2003.370 144.400 2003.690 144.460 ;
        RECT 2002.450 144.260 2003.690 144.400 ;
        RECT 2002.450 144.200 2002.770 144.260 ;
        RECT 2003.370 144.200 2003.690 144.260 ;
        RECT 2002.450 62.460 2002.770 62.520 ;
        RECT 2002.080 62.320 2002.770 62.460 ;
        RECT 2002.080 62.180 2002.220 62.320 ;
        RECT 2002.450 62.260 2002.770 62.320 ;
        RECT 2001.990 61.920 2002.310 62.180 ;
        RECT 1668.030 21.320 1668.350 21.380 ;
        RECT 2001.990 21.320 2002.310 21.380 ;
        RECT 1668.030 21.180 2002.310 21.320 ;
        RECT 1668.030 21.120 1668.350 21.180 ;
        RECT 2001.990 21.120 2002.310 21.180 ;
      LAYER via ;
        RECT 2001.560 1641.900 2001.820 1642.160 ;
        RECT 2002.940 1641.900 2003.200 1642.160 ;
        RECT 2001.560 1635.100 2001.820 1635.360 ;
        RECT 2002.480 1593.960 2002.740 1594.220 ;
        RECT 2002.480 1579.680 2002.740 1579.940 ;
        RECT 2002.480 1497.060 2002.740 1497.320 ;
        RECT 2002.480 1414.100 2002.740 1414.360 ;
        RECT 2002.480 1413.420 2002.740 1413.680 ;
        RECT 2002.020 1365.820 2002.280 1366.080 ;
        RECT 2002.940 1365.820 2003.200 1366.080 ;
        RECT 2002.940 1352.220 2003.200 1352.480 ;
        RECT 2002.480 1304.280 2002.740 1304.540 ;
        RECT 2002.020 1269.260 2002.280 1269.520 ;
        RECT 2002.940 1269.260 2003.200 1269.520 ;
        RECT 2002.940 1255.660 2003.200 1255.920 ;
        RECT 2002.480 1207.380 2002.740 1207.640 ;
        RECT 2002.020 1172.700 2002.280 1172.960 ;
        RECT 2002.940 1172.700 2003.200 1172.960 ;
        RECT 2002.020 1110.820 2002.280 1111.080 ;
        RECT 2002.480 1110.820 2002.740 1111.080 ;
        RECT 2001.560 1062.540 2001.820 1062.800 ;
        RECT 2002.940 1062.540 2003.200 1062.800 ;
        RECT 2002.480 1013.920 2002.740 1014.180 ;
        RECT 2002.940 1013.920 2003.200 1014.180 ;
        RECT 2002.020 835.080 2002.280 835.340 ;
        RECT 2002.940 835.080 2003.200 835.340 ;
        RECT 2002.480 820.800 2002.740 821.060 ;
        RECT 2002.480 786.460 2002.740 786.720 ;
        RECT 2002.020 738.180 2002.280 738.440 ;
        RECT 2002.940 738.180 2003.200 738.440 ;
        RECT 2002.480 724.240 2002.740 724.500 ;
        RECT 2002.480 689.560 2002.740 689.820 ;
        RECT 2002.480 628.020 2002.740 628.280 ;
        RECT 2002.940 628.020 2003.200 628.280 ;
        RECT 2002.020 579.740 2002.280 580.000 ;
        RECT 2002.480 579.740 2002.740 580.000 ;
        RECT 2002.480 523.980 2002.740 524.240 ;
        RECT 2002.940 476.040 2003.200 476.300 ;
        RECT 2002.480 338.000 2002.740 338.260 ;
        RECT 2002.940 338.000 2003.200 338.260 ;
        RECT 2002.940 235.660 2003.200 235.920 ;
        RECT 2002.940 227.840 2003.200 228.100 ;
        RECT 2003.400 227.160 2003.660 227.420 ;
        RECT 2003.400 185.680 2003.660 185.940 ;
        RECT 2002.480 144.200 2002.740 144.460 ;
        RECT 2003.400 144.200 2003.660 144.460 ;
        RECT 2002.480 62.260 2002.740 62.520 ;
        RECT 2002.020 61.920 2002.280 62.180 ;
        RECT 1668.060 21.120 1668.320 21.380 ;
        RECT 2002.020 21.120 2002.280 21.380 ;
      LAYER met2 ;
        RECT 2007.000 1700.410 2007.280 1704.000 ;
        RECT 2004.380 1700.270 2007.280 1700.410 ;
        RECT 2004.380 1677.970 2004.520 1700.270 ;
        RECT 2007.000 1700.000 2007.280 1700.270 ;
        RECT 2003.000 1677.830 2004.520 1677.970 ;
        RECT 2003.000 1642.190 2003.140 1677.830 ;
        RECT 2001.560 1641.870 2001.820 1642.190 ;
        RECT 2002.940 1641.870 2003.200 1642.190 ;
        RECT 2001.620 1635.390 2001.760 1641.870 ;
        RECT 2001.560 1635.070 2001.820 1635.390 ;
        RECT 2002.480 1593.930 2002.740 1594.250 ;
        RECT 2002.540 1579.970 2002.680 1593.930 ;
        RECT 2002.480 1579.650 2002.740 1579.970 ;
        RECT 2002.480 1497.030 2002.740 1497.350 ;
        RECT 2002.540 1414.390 2002.680 1497.030 ;
        RECT 2002.480 1414.070 2002.740 1414.390 ;
        RECT 2002.480 1413.390 2002.740 1413.710 ;
        RECT 2002.540 1366.530 2002.680 1413.390 ;
        RECT 2002.080 1366.390 2002.680 1366.530 ;
        RECT 2002.080 1366.110 2002.220 1366.390 ;
        RECT 2002.020 1365.790 2002.280 1366.110 ;
        RECT 2002.940 1365.790 2003.200 1366.110 ;
        RECT 2003.000 1352.510 2003.140 1365.790 ;
        RECT 2002.940 1352.190 2003.200 1352.510 ;
        RECT 2002.480 1304.250 2002.740 1304.570 ;
        RECT 2002.540 1269.970 2002.680 1304.250 ;
        RECT 2002.080 1269.830 2002.680 1269.970 ;
        RECT 2002.080 1269.550 2002.220 1269.830 ;
        RECT 2002.020 1269.230 2002.280 1269.550 ;
        RECT 2002.940 1269.230 2003.200 1269.550 ;
        RECT 2003.000 1255.950 2003.140 1269.230 ;
        RECT 2002.940 1255.630 2003.200 1255.950 ;
        RECT 2002.480 1207.350 2002.740 1207.670 ;
        RECT 2002.540 1173.410 2002.680 1207.350 ;
        RECT 2002.080 1173.270 2002.680 1173.410 ;
        RECT 2002.080 1172.990 2002.220 1173.270 ;
        RECT 2002.020 1172.670 2002.280 1172.990 ;
        RECT 2002.940 1172.670 2003.200 1172.990 ;
        RECT 2003.000 1159.245 2003.140 1172.670 ;
        RECT 2002.010 1158.875 2002.290 1159.245 ;
        RECT 2002.930 1158.875 2003.210 1159.245 ;
        RECT 2002.080 1111.110 2002.220 1158.875 ;
        RECT 2001.550 1110.595 2001.830 1110.965 ;
        RECT 2002.020 1110.790 2002.280 1111.110 ;
        RECT 2002.480 1110.965 2002.740 1111.110 ;
        RECT 2002.470 1110.595 2002.750 1110.965 ;
        RECT 2001.620 1062.830 2001.760 1110.595 ;
        RECT 2001.560 1062.510 2001.820 1062.830 ;
        RECT 2002.940 1062.510 2003.200 1062.830 ;
        RECT 2003.000 1027.890 2003.140 1062.510 ;
        RECT 2002.540 1027.750 2003.140 1027.890 ;
        RECT 2002.540 1014.210 2002.680 1027.750 ;
        RECT 2002.480 1013.890 2002.740 1014.210 ;
        RECT 2002.940 1013.890 2003.200 1014.210 ;
        RECT 2003.000 835.370 2003.140 1013.890 ;
        RECT 2002.020 835.050 2002.280 835.370 ;
        RECT 2002.940 835.050 2003.200 835.370 ;
        RECT 2002.080 834.770 2002.220 835.050 ;
        RECT 2002.080 834.630 2002.680 834.770 ;
        RECT 2002.540 821.090 2002.680 834.630 ;
        RECT 2002.480 820.770 2002.740 821.090 ;
        RECT 2002.480 786.430 2002.740 786.750 ;
        RECT 2002.540 772.890 2002.680 786.430 ;
        RECT 2002.540 772.750 2003.140 772.890 ;
        RECT 2003.000 738.470 2003.140 772.750 ;
        RECT 2002.020 738.210 2002.280 738.470 ;
        RECT 2002.020 738.150 2002.680 738.210 ;
        RECT 2002.940 738.150 2003.200 738.470 ;
        RECT 2002.080 738.070 2002.680 738.150 ;
        RECT 2002.540 724.530 2002.680 738.070 ;
        RECT 2002.480 724.210 2002.740 724.530 ;
        RECT 2002.480 689.530 2002.740 689.850 ;
        RECT 2002.540 676.330 2002.680 689.530 ;
        RECT 2002.540 676.190 2003.140 676.330 ;
        RECT 2003.000 628.310 2003.140 676.190 ;
        RECT 2002.480 627.990 2002.740 628.310 ;
        RECT 2002.940 627.990 2003.200 628.310 ;
        RECT 2002.540 580.030 2002.680 627.990 ;
        RECT 2002.020 579.710 2002.280 580.030 ;
        RECT 2002.480 579.710 2002.740 580.030 ;
        RECT 2002.080 555.290 2002.220 579.710 ;
        RECT 2002.080 555.150 2002.680 555.290 ;
        RECT 2002.540 524.270 2002.680 555.150 ;
        RECT 2002.480 523.950 2002.740 524.270 ;
        RECT 2002.940 476.010 2003.200 476.330 ;
        RECT 2003.000 338.290 2003.140 476.010 ;
        RECT 2002.480 337.970 2002.740 338.290 ;
        RECT 2002.940 337.970 2003.200 338.290 ;
        RECT 2002.540 303.690 2002.680 337.970 ;
        RECT 2002.540 303.550 2003.140 303.690 ;
        RECT 2003.000 235.950 2003.140 303.550 ;
        RECT 2002.940 235.630 2003.200 235.950 ;
        RECT 2002.940 227.810 2003.200 228.130 ;
        RECT 2003.000 227.530 2003.140 227.810 ;
        RECT 2003.000 227.450 2003.600 227.530 ;
        RECT 2003.000 227.390 2003.660 227.450 ;
        RECT 2003.400 227.130 2003.660 227.390 ;
        RECT 2003.400 185.650 2003.660 185.970 ;
        RECT 2003.460 144.490 2003.600 185.650 ;
        RECT 2002.480 144.170 2002.740 144.490 ;
        RECT 2003.400 144.170 2003.660 144.490 ;
        RECT 2002.540 62.550 2002.680 144.170 ;
        RECT 2002.480 62.230 2002.740 62.550 ;
        RECT 2002.020 61.890 2002.280 62.210 ;
        RECT 2002.080 21.410 2002.220 61.890 ;
        RECT 1668.060 21.090 1668.320 21.410 ;
        RECT 2002.020 21.090 2002.280 21.410 ;
        RECT 1668.120 2.400 1668.260 21.090 ;
        RECT 1667.910 -4.800 1668.470 2.400 ;
      LAYER via2 ;
        RECT 2002.010 1158.920 2002.290 1159.200 ;
        RECT 2002.930 1158.920 2003.210 1159.200 ;
        RECT 2001.550 1110.640 2001.830 1110.920 ;
        RECT 2002.470 1110.640 2002.750 1110.920 ;
      LAYER met3 ;
        RECT 2001.985 1159.210 2002.315 1159.225 ;
        RECT 2002.905 1159.210 2003.235 1159.225 ;
        RECT 2001.985 1158.910 2003.235 1159.210 ;
        RECT 2001.985 1158.895 2002.315 1158.910 ;
        RECT 2002.905 1158.895 2003.235 1158.910 ;
        RECT 2001.525 1110.930 2001.855 1110.945 ;
        RECT 2002.445 1110.930 2002.775 1110.945 ;
        RECT 2001.525 1110.630 2002.775 1110.930 ;
        RECT 2001.525 1110.615 2001.855 1110.630 ;
        RECT 2002.445 1110.615 2002.775 1110.630 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1685.510 20.980 1685.830 21.040 ;
        RECT 2015.330 20.980 2015.650 21.040 ;
        RECT 1685.510 20.840 2015.650 20.980 ;
        RECT 1685.510 20.780 1685.830 20.840 ;
        RECT 2015.330 20.780 2015.650 20.840 ;
      LAYER via ;
        RECT 1685.540 20.780 1685.800 21.040 ;
        RECT 2015.360 20.780 2015.620 21.040 ;
      LAYER met2 ;
        RECT 2016.200 1700.410 2016.480 1704.000 ;
        RECT 2015.420 1700.270 2016.480 1700.410 ;
        RECT 2015.420 21.070 2015.560 1700.270 ;
        RECT 2016.200 1700.000 2016.480 1700.270 ;
        RECT 1685.540 20.750 1685.800 21.070 ;
        RECT 2015.360 20.750 2015.620 21.070 ;
        RECT 1685.600 2.400 1685.740 20.750 ;
        RECT 1685.390 -4.800 1685.950 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 724.110 66.200 724.430 66.260 ;
        RECT 1518.530 66.200 1518.850 66.260 ;
        RECT 724.110 66.060 1518.850 66.200 ;
        RECT 724.110 66.000 724.430 66.060 ;
        RECT 1518.530 66.000 1518.850 66.060 ;
      LAYER via ;
        RECT 724.140 66.000 724.400 66.260 ;
        RECT 1518.560 66.000 1518.820 66.260 ;
      LAYER met2 ;
        RECT 1520.320 1700.410 1520.600 1704.000 ;
        RECT 1518.620 1700.270 1520.600 1700.410 ;
        RECT 1518.620 66.290 1518.760 1700.270 ;
        RECT 1520.320 1700.000 1520.600 1700.270 ;
        RECT 724.140 65.970 724.400 66.290 ;
        RECT 1518.560 65.970 1518.820 66.290 ;
        RECT 724.200 16.730 724.340 65.970 ;
        RECT 722.360 16.590 724.340 16.730 ;
        RECT 722.360 2.400 722.500 16.590 ;
        RECT 722.150 -4.800 722.710 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1703.450 23.700 1703.770 23.760 ;
        RECT 2022.690 23.700 2023.010 23.760 ;
        RECT 1703.450 23.560 2023.010 23.700 ;
        RECT 1703.450 23.500 1703.770 23.560 ;
        RECT 2022.690 23.500 2023.010 23.560 ;
      LAYER via ;
        RECT 1703.480 23.500 1703.740 23.760 ;
        RECT 2022.720 23.500 2022.980 23.760 ;
      LAYER met2 ;
        RECT 2025.400 1700.410 2025.680 1704.000 ;
        RECT 2022.780 1700.270 2025.680 1700.410 ;
        RECT 2022.780 23.790 2022.920 1700.270 ;
        RECT 2025.400 1700.000 2025.680 1700.270 ;
        RECT 1703.480 23.470 1703.740 23.790 ;
        RECT 2022.720 23.470 2022.980 23.790 ;
        RECT 1703.540 2.400 1703.680 23.470 ;
        RECT 1703.330 -4.800 1703.890 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2029.590 1678.140 2029.910 1678.200 ;
        RECT 2033.270 1678.140 2033.590 1678.200 ;
        RECT 2029.590 1678.000 2033.590 1678.140 ;
        RECT 2029.590 1677.940 2029.910 1678.000 ;
        RECT 2033.270 1677.940 2033.590 1678.000 ;
        RECT 1721.390 23.360 1721.710 23.420 ;
        RECT 2029.590 23.360 2029.910 23.420 ;
        RECT 1721.390 23.220 2029.910 23.360 ;
        RECT 1721.390 23.160 1721.710 23.220 ;
        RECT 2029.590 23.160 2029.910 23.220 ;
      LAYER via ;
        RECT 2029.620 1677.940 2029.880 1678.200 ;
        RECT 2033.300 1677.940 2033.560 1678.200 ;
        RECT 1721.420 23.160 1721.680 23.420 ;
        RECT 2029.620 23.160 2029.880 23.420 ;
      LAYER met2 ;
        RECT 2034.600 1700.410 2034.880 1704.000 ;
        RECT 2033.360 1700.270 2034.880 1700.410 ;
        RECT 2033.360 1678.230 2033.500 1700.270 ;
        RECT 2034.600 1700.000 2034.880 1700.270 ;
        RECT 2029.620 1677.910 2029.880 1678.230 ;
        RECT 2033.300 1677.910 2033.560 1678.230 ;
        RECT 2029.680 23.450 2029.820 1677.910 ;
        RECT 1721.420 23.130 1721.680 23.450 ;
        RECT 2029.620 23.130 2029.880 23.450 ;
        RECT 1721.480 2.400 1721.620 23.130 ;
        RECT 1721.270 -4.800 1721.830 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1739.330 24.040 1739.650 24.100 ;
        RECT 2042.470 24.040 2042.790 24.100 ;
        RECT 1739.330 23.900 2042.790 24.040 ;
        RECT 1739.330 23.840 1739.650 23.900 ;
        RECT 2042.470 23.840 2042.790 23.900 ;
      LAYER via ;
        RECT 1739.360 23.840 1739.620 24.100 ;
        RECT 2042.500 23.840 2042.760 24.100 ;
      LAYER met2 ;
        RECT 2043.800 1700.410 2044.080 1704.000 ;
        RECT 2042.560 1700.270 2044.080 1700.410 ;
        RECT 2042.560 24.130 2042.700 1700.270 ;
        RECT 2043.800 1700.000 2044.080 1700.270 ;
        RECT 1739.360 23.810 1739.620 24.130 ;
        RECT 2042.500 23.810 2042.760 24.130 ;
        RECT 1739.420 2.400 1739.560 23.810 ;
        RECT 1739.210 -4.800 1739.770 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1756.810 24.380 1757.130 24.440 ;
        RECT 2050.290 24.380 2050.610 24.440 ;
        RECT 1756.810 24.240 2050.610 24.380 ;
        RECT 1756.810 24.180 1757.130 24.240 ;
        RECT 2050.290 24.180 2050.610 24.240 ;
      LAYER via ;
        RECT 1756.840 24.180 1757.100 24.440 ;
        RECT 2050.320 24.180 2050.580 24.440 ;
      LAYER met2 ;
        RECT 2053.000 1700.410 2053.280 1704.000 ;
        RECT 2050.380 1700.270 2053.280 1700.410 ;
        RECT 2050.380 24.470 2050.520 1700.270 ;
        RECT 2053.000 1700.000 2053.280 1700.270 ;
        RECT 1756.840 24.150 1757.100 24.470 ;
        RECT 2050.320 24.150 2050.580 24.470 ;
        RECT 1756.900 2.400 1757.040 24.150 ;
        RECT 1756.690 -4.800 1757.250 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1774.750 30.160 1775.070 30.220 ;
        RECT 2056.730 30.160 2057.050 30.220 ;
        RECT 1774.750 30.020 2057.050 30.160 ;
        RECT 1774.750 29.960 1775.070 30.020 ;
        RECT 2056.730 29.960 2057.050 30.020 ;
      LAYER via ;
        RECT 1774.780 29.960 1775.040 30.220 ;
        RECT 2056.760 29.960 2057.020 30.220 ;
      LAYER met2 ;
        RECT 2062.200 1700.410 2062.480 1704.000 ;
        RECT 2059.580 1700.270 2062.480 1700.410 ;
        RECT 2059.580 1677.970 2059.720 1700.270 ;
        RECT 2062.200 1700.000 2062.480 1700.270 ;
        RECT 2056.820 1677.830 2059.720 1677.970 ;
        RECT 2056.820 30.250 2056.960 1677.830 ;
        RECT 1774.780 29.930 1775.040 30.250 ;
        RECT 2056.760 29.930 2057.020 30.250 ;
        RECT 1774.840 2.400 1774.980 29.930 ;
        RECT 1774.630 -4.800 1775.190 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1792.690 24.720 1793.010 24.780 ;
        RECT 2070.530 24.720 2070.850 24.780 ;
        RECT 1792.690 24.580 2070.850 24.720 ;
        RECT 1792.690 24.520 1793.010 24.580 ;
        RECT 2070.530 24.520 2070.850 24.580 ;
      LAYER via ;
        RECT 1792.720 24.520 1792.980 24.780 ;
        RECT 2070.560 24.520 2070.820 24.780 ;
      LAYER met2 ;
        RECT 2071.400 1700.410 2071.680 1704.000 ;
        RECT 2070.620 1700.270 2071.680 1700.410 ;
        RECT 2070.620 24.810 2070.760 1700.270 ;
        RECT 2071.400 1700.000 2071.680 1700.270 ;
        RECT 1792.720 24.490 1792.980 24.810 ;
        RECT 2070.560 24.490 2070.820 24.810 ;
        RECT 1792.780 2.400 1792.920 24.490 ;
        RECT 1792.570 -4.800 1793.130 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1810.630 29.480 1810.950 29.540 ;
        RECT 2077.890 29.480 2078.210 29.540 ;
        RECT 1810.630 29.340 2078.210 29.480 ;
        RECT 1810.630 29.280 1810.950 29.340 ;
        RECT 2077.890 29.280 2078.210 29.340 ;
      LAYER via ;
        RECT 1810.660 29.280 1810.920 29.540 ;
        RECT 2077.920 29.280 2078.180 29.540 ;
      LAYER met2 ;
        RECT 2080.600 1700.410 2080.880 1704.000 ;
        RECT 2077.980 1700.270 2080.880 1700.410 ;
        RECT 2077.980 29.570 2078.120 1700.270 ;
        RECT 2080.600 1700.000 2080.880 1700.270 ;
        RECT 1810.660 29.250 1810.920 29.570 ;
        RECT 2077.920 29.250 2078.180 29.570 ;
        RECT 1810.720 2.400 1810.860 29.250 ;
        RECT 1810.510 -4.800 1811.070 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2084.405 1594.005 2084.575 1642.115 ;
        RECT 2084.405 1497.445 2084.575 1545.555 ;
        RECT 2084.405 1352.605 2084.575 1400.715 ;
        RECT 2084.405 1256.045 2084.575 1304.155 ;
        RECT 2084.405 241.825 2084.575 289.595 ;
      LAYER mcon ;
        RECT 2084.405 1641.945 2084.575 1642.115 ;
        RECT 2084.405 1545.385 2084.575 1545.555 ;
        RECT 2084.405 1400.545 2084.575 1400.715 ;
        RECT 2084.405 1303.985 2084.575 1304.155 ;
        RECT 2084.405 289.425 2084.575 289.595 ;
      LAYER met1 ;
        RECT 2083.870 1656.040 2084.190 1656.100 ;
        RECT 2084.790 1656.040 2085.110 1656.100 ;
        RECT 2083.870 1655.900 2085.110 1656.040 ;
        RECT 2083.870 1655.840 2084.190 1655.900 ;
        RECT 2084.790 1655.840 2085.110 1655.900 ;
        RECT 2084.345 1642.100 2084.635 1642.145 ;
        RECT 2084.790 1642.100 2085.110 1642.160 ;
        RECT 2084.345 1641.960 2085.110 1642.100 ;
        RECT 2084.345 1641.915 2084.635 1641.960 ;
        RECT 2084.790 1641.900 2085.110 1641.960 ;
        RECT 2084.330 1594.160 2084.650 1594.220 ;
        RECT 2084.135 1594.020 2084.650 1594.160 ;
        RECT 2084.330 1593.960 2084.650 1594.020 ;
        RECT 2083.870 1559.140 2084.190 1559.200 ;
        RECT 2084.790 1559.140 2085.110 1559.200 ;
        RECT 2083.870 1559.000 2085.110 1559.140 ;
        RECT 2083.870 1558.940 2084.190 1559.000 ;
        RECT 2084.790 1558.940 2085.110 1559.000 ;
        RECT 2084.345 1545.540 2084.635 1545.585 ;
        RECT 2084.790 1545.540 2085.110 1545.600 ;
        RECT 2084.345 1545.400 2085.110 1545.540 ;
        RECT 2084.345 1545.355 2084.635 1545.400 ;
        RECT 2084.790 1545.340 2085.110 1545.400 ;
        RECT 2084.330 1497.600 2084.650 1497.660 ;
        RECT 2084.135 1497.460 2084.650 1497.600 ;
        RECT 2084.330 1497.400 2084.650 1497.460 ;
        RECT 2084.330 1400.700 2084.650 1400.760 ;
        RECT 2084.135 1400.560 2084.650 1400.700 ;
        RECT 2084.330 1400.500 2084.650 1400.560 ;
        RECT 2084.345 1352.760 2084.635 1352.805 ;
        RECT 2084.790 1352.760 2085.110 1352.820 ;
        RECT 2084.345 1352.620 2085.110 1352.760 ;
        RECT 2084.345 1352.575 2084.635 1352.620 ;
        RECT 2084.790 1352.560 2085.110 1352.620 ;
        RECT 2084.330 1304.140 2084.650 1304.200 ;
        RECT 2084.135 1304.000 2084.650 1304.140 ;
        RECT 2084.330 1303.940 2084.650 1304.000 ;
        RECT 2084.345 1256.200 2084.635 1256.245 ;
        RECT 2084.790 1256.200 2085.110 1256.260 ;
        RECT 2084.345 1256.060 2085.110 1256.200 ;
        RECT 2084.345 1256.015 2084.635 1256.060 ;
        RECT 2084.790 1256.000 2085.110 1256.060 ;
        RECT 2084.790 1159.300 2085.110 1159.360 ;
        RECT 2085.710 1159.300 2086.030 1159.360 ;
        RECT 2084.790 1159.160 2086.030 1159.300 ;
        RECT 2084.790 1159.100 2085.110 1159.160 ;
        RECT 2085.710 1159.100 2086.030 1159.160 ;
        RECT 2084.790 1062.740 2085.110 1062.800 ;
        RECT 2085.710 1062.740 2086.030 1062.800 ;
        RECT 2084.790 1062.600 2086.030 1062.740 ;
        RECT 2084.790 1062.540 2085.110 1062.600 ;
        RECT 2085.710 1062.540 2086.030 1062.600 ;
        RECT 2084.790 966.180 2085.110 966.240 ;
        RECT 2085.710 966.180 2086.030 966.240 ;
        RECT 2084.790 966.040 2086.030 966.180 ;
        RECT 2084.790 965.980 2085.110 966.040 ;
        RECT 2085.710 965.980 2086.030 966.040 ;
        RECT 2084.330 917.560 2084.650 917.620 ;
        RECT 2084.790 917.560 2085.110 917.620 ;
        RECT 2084.330 917.420 2085.110 917.560 ;
        RECT 2084.330 917.360 2084.650 917.420 ;
        RECT 2084.790 917.360 2085.110 917.420 ;
        RECT 2084.330 821.000 2084.650 821.060 ;
        RECT 2084.790 821.000 2085.110 821.060 ;
        RECT 2084.330 820.860 2085.110 821.000 ;
        RECT 2084.330 820.800 2084.650 820.860 ;
        RECT 2084.790 820.800 2085.110 820.860 ;
        RECT 2084.330 689.900 2084.650 690.160 ;
        RECT 2083.870 689.760 2084.190 689.820 ;
        RECT 2084.420 689.760 2084.560 689.900 ;
        RECT 2083.870 689.620 2084.560 689.760 ;
        RECT 2083.870 689.560 2084.190 689.620 ;
        RECT 2084.330 593.340 2084.650 593.600 ;
        RECT 2083.870 593.200 2084.190 593.260 ;
        RECT 2084.420 593.200 2084.560 593.340 ;
        RECT 2083.870 593.060 2084.560 593.200 ;
        RECT 2083.870 593.000 2084.190 593.060 ;
        RECT 2084.330 496.780 2084.650 497.040 ;
        RECT 2083.870 496.640 2084.190 496.700 ;
        RECT 2084.420 496.640 2084.560 496.780 ;
        RECT 2083.870 496.500 2084.560 496.640 ;
        RECT 2083.870 496.440 2084.190 496.500 ;
        RECT 2084.330 386.820 2084.650 386.880 ;
        RECT 2084.790 386.820 2085.110 386.880 ;
        RECT 2084.330 386.680 2085.110 386.820 ;
        RECT 2084.330 386.620 2084.650 386.680 ;
        RECT 2084.790 386.620 2085.110 386.680 ;
        RECT 2084.790 352.480 2085.110 352.540 ;
        RECT 2084.420 352.340 2085.110 352.480 ;
        RECT 2084.420 351.860 2084.560 352.340 ;
        RECT 2084.790 352.280 2085.110 352.340 ;
        RECT 2084.330 351.600 2084.650 351.860 ;
        RECT 2084.330 337.860 2084.650 337.920 ;
        RECT 2085.250 337.860 2085.570 337.920 ;
        RECT 2084.330 337.720 2085.570 337.860 ;
        RECT 2084.330 337.660 2084.650 337.720 ;
        RECT 2085.250 337.660 2085.570 337.720 ;
        RECT 2084.345 289.580 2084.635 289.625 ;
        RECT 2084.790 289.580 2085.110 289.640 ;
        RECT 2084.345 289.440 2085.110 289.580 ;
        RECT 2084.345 289.395 2084.635 289.440 ;
        RECT 2084.790 289.380 2085.110 289.440 ;
        RECT 2084.330 241.980 2084.650 242.040 ;
        RECT 2084.135 241.840 2084.650 241.980 ;
        RECT 2084.330 241.780 2084.650 241.840 ;
        RECT 2084.330 241.300 2084.650 241.360 ;
        RECT 2085.250 241.300 2085.570 241.360 ;
        RECT 2084.330 241.160 2085.570 241.300 ;
        RECT 2084.330 241.100 2084.650 241.160 ;
        RECT 2085.250 241.100 2085.570 241.160 ;
        RECT 2084.790 159.020 2085.110 159.080 ;
        RECT 2084.420 158.880 2085.110 159.020 ;
        RECT 2084.420 158.740 2084.560 158.880 ;
        RECT 2084.790 158.820 2085.110 158.880 ;
        RECT 2084.330 158.480 2084.650 158.740 ;
        RECT 2083.870 110.400 2084.190 110.460 ;
        RECT 2084.790 110.400 2085.110 110.460 ;
        RECT 2083.870 110.260 2085.110 110.400 ;
        RECT 2083.870 110.200 2084.190 110.260 ;
        RECT 2084.790 110.200 2085.110 110.260 ;
        RECT 2084.790 59.540 2085.110 59.800 ;
        RECT 2084.880 59.120 2085.020 59.540 ;
        RECT 2084.790 58.860 2085.110 59.120 ;
        RECT 1828.570 25.060 1828.890 25.120 ;
        RECT 2084.790 25.060 2085.110 25.120 ;
        RECT 1828.570 24.920 2085.110 25.060 ;
        RECT 1828.570 24.860 1828.890 24.920 ;
        RECT 2084.790 24.860 2085.110 24.920 ;
      LAYER via ;
        RECT 2083.900 1655.840 2084.160 1656.100 ;
        RECT 2084.820 1655.840 2085.080 1656.100 ;
        RECT 2084.820 1641.900 2085.080 1642.160 ;
        RECT 2084.360 1593.960 2084.620 1594.220 ;
        RECT 2083.900 1558.940 2084.160 1559.200 ;
        RECT 2084.820 1558.940 2085.080 1559.200 ;
        RECT 2084.820 1545.340 2085.080 1545.600 ;
        RECT 2084.360 1497.400 2084.620 1497.660 ;
        RECT 2084.360 1400.500 2084.620 1400.760 ;
        RECT 2084.820 1352.560 2085.080 1352.820 ;
        RECT 2084.360 1303.940 2084.620 1304.200 ;
        RECT 2084.820 1256.000 2085.080 1256.260 ;
        RECT 2084.820 1159.100 2085.080 1159.360 ;
        RECT 2085.740 1159.100 2086.000 1159.360 ;
        RECT 2084.820 1062.540 2085.080 1062.800 ;
        RECT 2085.740 1062.540 2086.000 1062.800 ;
        RECT 2084.820 965.980 2085.080 966.240 ;
        RECT 2085.740 965.980 2086.000 966.240 ;
        RECT 2084.360 917.360 2084.620 917.620 ;
        RECT 2084.820 917.360 2085.080 917.620 ;
        RECT 2084.360 820.800 2084.620 821.060 ;
        RECT 2084.820 820.800 2085.080 821.060 ;
        RECT 2084.360 689.900 2084.620 690.160 ;
        RECT 2083.900 689.560 2084.160 689.820 ;
        RECT 2084.360 593.340 2084.620 593.600 ;
        RECT 2083.900 593.000 2084.160 593.260 ;
        RECT 2084.360 496.780 2084.620 497.040 ;
        RECT 2083.900 496.440 2084.160 496.700 ;
        RECT 2084.360 386.620 2084.620 386.880 ;
        RECT 2084.820 386.620 2085.080 386.880 ;
        RECT 2084.820 352.280 2085.080 352.540 ;
        RECT 2084.360 351.600 2084.620 351.860 ;
        RECT 2084.360 337.660 2084.620 337.920 ;
        RECT 2085.280 337.660 2085.540 337.920 ;
        RECT 2084.820 289.380 2085.080 289.640 ;
        RECT 2084.360 241.780 2084.620 242.040 ;
        RECT 2084.360 241.100 2084.620 241.360 ;
        RECT 2085.280 241.100 2085.540 241.360 ;
        RECT 2084.820 158.820 2085.080 159.080 ;
        RECT 2084.360 158.480 2084.620 158.740 ;
        RECT 2083.900 110.200 2084.160 110.460 ;
        RECT 2084.820 110.200 2085.080 110.460 ;
        RECT 2084.820 59.540 2085.080 59.800 ;
        RECT 2084.820 58.860 2085.080 59.120 ;
        RECT 1828.600 24.860 1828.860 25.120 ;
        RECT 2084.820 24.860 2085.080 25.120 ;
      LAYER met2 ;
        RECT 2089.800 1700.410 2090.080 1704.000 ;
        RECT 2087.180 1700.270 2090.080 1700.410 ;
        RECT 2087.180 1677.970 2087.320 1700.270 ;
        RECT 2089.800 1700.000 2090.080 1700.270 ;
        RECT 2083.960 1677.830 2087.320 1677.970 ;
        RECT 2083.960 1656.130 2084.100 1677.830 ;
        RECT 2083.900 1655.810 2084.160 1656.130 ;
        RECT 2084.820 1655.810 2085.080 1656.130 ;
        RECT 2084.880 1642.190 2085.020 1655.810 ;
        RECT 2084.820 1641.870 2085.080 1642.190 ;
        RECT 2084.360 1593.930 2084.620 1594.250 ;
        RECT 2084.420 1559.650 2084.560 1593.930 ;
        RECT 2083.960 1559.510 2084.560 1559.650 ;
        RECT 2083.960 1559.230 2084.100 1559.510 ;
        RECT 2083.900 1558.910 2084.160 1559.230 ;
        RECT 2084.820 1558.910 2085.080 1559.230 ;
        RECT 2084.880 1545.630 2085.020 1558.910 ;
        RECT 2084.820 1545.310 2085.080 1545.630 ;
        RECT 2084.360 1497.370 2084.620 1497.690 ;
        RECT 2084.420 1473.290 2084.560 1497.370 ;
        RECT 2084.420 1473.150 2085.020 1473.290 ;
        RECT 2084.880 1414.130 2085.020 1473.150 ;
        RECT 2084.420 1413.990 2085.020 1414.130 ;
        RECT 2084.420 1400.790 2084.560 1413.990 ;
        RECT 2084.360 1400.470 2084.620 1400.790 ;
        RECT 2084.820 1352.530 2085.080 1352.850 ;
        RECT 2084.880 1317.570 2085.020 1352.530 ;
        RECT 2084.420 1317.430 2085.020 1317.570 ;
        RECT 2084.420 1304.230 2084.560 1317.430 ;
        RECT 2084.360 1303.910 2084.620 1304.230 ;
        RECT 2084.820 1255.970 2085.080 1256.290 ;
        RECT 2084.880 1221.010 2085.020 1255.970 ;
        RECT 2084.420 1220.870 2085.020 1221.010 ;
        RECT 2084.420 1207.525 2084.560 1220.870 ;
        RECT 2084.350 1207.155 2084.630 1207.525 ;
        RECT 2085.730 1207.155 2086.010 1207.525 ;
        RECT 2085.800 1159.390 2085.940 1207.155 ;
        RECT 2084.820 1159.070 2085.080 1159.390 ;
        RECT 2085.740 1159.070 2086.000 1159.390 ;
        RECT 2084.880 1124.450 2085.020 1159.070 ;
        RECT 2084.420 1124.310 2085.020 1124.450 ;
        RECT 2084.420 1110.965 2084.560 1124.310 ;
        RECT 2084.350 1110.595 2084.630 1110.965 ;
        RECT 2085.730 1110.595 2086.010 1110.965 ;
        RECT 2085.800 1062.830 2085.940 1110.595 ;
        RECT 2084.820 1062.510 2085.080 1062.830 ;
        RECT 2085.740 1062.510 2086.000 1062.830 ;
        RECT 2084.880 1027.890 2085.020 1062.510 ;
        RECT 2084.420 1027.750 2085.020 1027.890 ;
        RECT 2084.420 1014.405 2084.560 1027.750 ;
        RECT 2084.350 1014.035 2084.630 1014.405 ;
        RECT 2085.730 1014.035 2086.010 1014.405 ;
        RECT 2085.800 966.270 2085.940 1014.035 ;
        RECT 2084.820 965.950 2085.080 966.270 ;
        RECT 2085.740 965.950 2086.000 966.270 ;
        RECT 2084.880 931.330 2085.020 965.950 ;
        RECT 2084.420 931.190 2085.020 931.330 ;
        RECT 2084.420 917.650 2084.560 931.190 ;
        RECT 2084.360 917.330 2084.620 917.650 ;
        RECT 2084.820 917.330 2085.080 917.650 ;
        RECT 2084.880 834.770 2085.020 917.330 ;
        RECT 2084.420 834.630 2085.020 834.770 ;
        RECT 2084.420 821.090 2084.560 834.630 ;
        RECT 2084.360 820.770 2084.620 821.090 ;
        RECT 2084.820 820.770 2085.080 821.090 ;
        RECT 2084.880 738.210 2085.020 820.770 ;
        RECT 2084.420 738.070 2085.020 738.210 ;
        RECT 2084.420 690.190 2084.560 738.070 ;
        RECT 2084.360 689.870 2084.620 690.190 ;
        RECT 2083.900 689.530 2084.160 689.850 ;
        RECT 2083.960 676.445 2084.100 689.530 ;
        RECT 2083.890 676.075 2084.170 676.445 ;
        RECT 2084.810 676.075 2085.090 676.445 ;
        RECT 2084.880 641.650 2085.020 676.075 ;
        RECT 2084.420 641.510 2085.020 641.650 ;
        RECT 2084.420 593.630 2084.560 641.510 ;
        RECT 2084.360 593.310 2084.620 593.630 ;
        RECT 2083.900 592.970 2084.160 593.290 ;
        RECT 2083.960 579.885 2084.100 592.970 ;
        RECT 2083.890 579.515 2084.170 579.885 ;
        RECT 2084.810 579.515 2085.090 579.885 ;
        RECT 2084.880 545.090 2085.020 579.515 ;
        RECT 2084.420 544.950 2085.020 545.090 ;
        RECT 2084.420 497.070 2084.560 544.950 ;
        RECT 2084.360 496.750 2084.620 497.070 ;
        RECT 2083.900 496.410 2084.160 496.730 ;
        RECT 2083.960 483.325 2084.100 496.410 ;
        RECT 2083.890 482.955 2084.170 483.325 ;
        RECT 2084.810 482.955 2085.090 483.325 ;
        RECT 2084.880 448.530 2085.020 482.955 ;
        RECT 2084.420 448.390 2085.020 448.530 ;
        RECT 2084.420 386.910 2084.560 448.390 ;
        RECT 2084.360 386.590 2084.620 386.910 ;
        RECT 2084.820 386.590 2085.080 386.910 ;
        RECT 2084.880 352.570 2085.020 386.590 ;
        RECT 2084.820 352.250 2085.080 352.570 ;
        RECT 2084.360 351.570 2084.620 351.890 ;
        RECT 2084.420 337.950 2084.560 351.570 ;
        RECT 2084.360 337.630 2084.620 337.950 ;
        RECT 2085.280 337.630 2085.540 337.950 ;
        RECT 2085.340 290.090 2085.480 337.630 ;
        RECT 2084.880 289.950 2085.480 290.090 ;
        RECT 2084.880 289.670 2085.020 289.950 ;
        RECT 2084.820 289.350 2085.080 289.670 ;
        RECT 2084.360 241.750 2084.620 242.070 ;
        RECT 2084.420 241.390 2084.560 241.750 ;
        RECT 2084.360 241.070 2084.620 241.390 ;
        RECT 2085.280 241.070 2085.540 241.390 ;
        RECT 2085.340 193.530 2085.480 241.070 ;
        RECT 2084.880 193.390 2085.480 193.530 ;
        RECT 2084.880 159.110 2085.020 193.390 ;
        RECT 2084.820 158.790 2085.080 159.110 ;
        RECT 2084.360 158.450 2084.620 158.770 ;
        RECT 2084.420 110.570 2084.560 158.450 ;
        RECT 2083.960 110.490 2084.560 110.570 ;
        RECT 2083.900 110.430 2084.560 110.490 ;
        RECT 2083.900 110.170 2084.160 110.430 ;
        RECT 2084.820 110.170 2085.080 110.490 ;
        RECT 2084.880 59.830 2085.020 110.170 ;
        RECT 2084.820 59.510 2085.080 59.830 ;
        RECT 2084.820 58.830 2085.080 59.150 ;
        RECT 2084.880 25.150 2085.020 58.830 ;
        RECT 1828.600 24.830 1828.860 25.150 ;
        RECT 2084.820 24.830 2085.080 25.150 ;
        RECT 1828.660 2.400 1828.800 24.830 ;
        RECT 1828.450 -4.800 1829.010 2.400 ;
      LAYER via2 ;
        RECT 2084.350 1207.200 2084.630 1207.480 ;
        RECT 2085.730 1207.200 2086.010 1207.480 ;
        RECT 2084.350 1110.640 2084.630 1110.920 ;
        RECT 2085.730 1110.640 2086.010 1110.920 ;
        RECT 2084.350 1014.080 2084.630 1014.360 ;
        RECT 2085.730 1014.080 2086.010 1014.360 ;
        RECT 2083.890 676.120 2084.170 676.400 ;
        RECT 2084.810 676.120 2085.090 676.400 ;
        RECT 2083.890 579.560 2084.170 579.840 ;
        RECT 2084.810 579.560 2085.090 579.840 ;
        RECT 2083.890 483.000 2084.170 483.280 ;
        RECT 2084.810 483.000 2085.090 483.280 ;
      LAYER met3 ;
        RECT 2084.325 1207.490 2084.655 1207.505 ;
        RECT 2085.705 1207.490 2086.035 1207.505 ;
        RECT 2084.325 1207.190 2086.035 1207.490 ;
        RECT 2084.325 1207.175 2084.655 1207.190 ;
        RECT 2085.705 1207.175 2086.035 1207.190 ;
        RECT 2084.325 1110.930 2084.655 1110.945 ;
        RECT 2085.705 1110.930 2086.035 1110.945 ;
        RECT 2084.325 1110.630 2086.035 1110.930 ;
        RECT 2084.325 1110.615 2084.655 1110.630 ;
        RECT 2085.705 1110.615 2086.035 1110.630 ;
        RECT 2084.325 1014.370 2084.655 1014.385 ;
        RECT 2085.705 1014.370 2086.035 1014.385 ;
        RECT 2084.325 1014.070 2086.035 1014.370 ;
        RECT 2084.325 1014.055 2084.655 1014.070 ;
        RECT 2085.705 1014.055 2086.035 1014.070 ;
        RECT 2083.865 676.410 2084.195 676.425 ;
        RECT 2084.785 676.410 2085.115 676.425 ;
        RECT 2083.865 676.110 2085.115 676.410 ;
        RECT 2083.865 676.095 2084.195 676.110 ;
        RECT 2084.785 676.095 2085.115 676.110 ;
        RECT 2083.865 579.850 2084.195 579.865 ;
        RECT 2084.785 579.850 2085.115 579.865 ;
        RECT 2083.865 579.550 2085.115 579.850 ;
        RECT 2083.865 579.535 2084.195 579.550 ;
        RECT 2084.785 579.535 2085.115 579.550 ;
        RECT 2083.865 483.290 2084.195 483.305 ;
        RECT 2084.785 483.290 2085.115 483.305 ;
        RECT 2083.865 482.990 2085.115 483.290 ;
        RECT 2083.865 482.975 2084.195 482.990 ;
        RECT 2084.785 482.975 2085.115 482.990 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1846.050 29.140 1846.370 29.200 ;
        RECT 2098.130 29.140 2098.450 29.200 ;
        RECT 1846.050 29.000 2098.450 29.140 ;
        RECT 1846.050 28.940 1846.370 29.000 ;
        RECT 2098.130 28.940 2098.450 29.000 ;
      LAYER via ;
        RECT 1846.080 28.940 1846.340 29.200 ;
        RECT 2098.160 28.940 2098.420 29.200 ;
      LAYER met2 ;
        RECT 2099.000 1700.410 2099.280 1704.000 ;
        RECT 2098.220 1700.270 2099.280 1700.410 ;
        RECT 2098.220 29.230 2098.360 1700.270 ;
        RECT 2099.000 1700.000 2099.280 1700.270 ;
        RECT 1846.080 28.910 1846.340 29.230 ;
        RECT 2098.160 28.910 2098.420 29.230 ;
        RECT 1846.140 2.400 1846.280 28.910 ;
        RECT 1845.930 -4.800 1846.490 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1864.450 30.840 1864.770 30.900 ;
        RECT 2105.490 30.840 2105.810 30.900 ;
        RECT 1864.450 30.700 2105.810 30.840 ;
        RECT 1864.450 30.640 1864.770 30.700 ;
        RECT 2105.490 30.640 2105.810 30.700 ;
      LAYER via ;
        RECT 1864.480 30.640 1864.740 30.900 ;
        RECT 2105.520 30.640 2105.780 30.900 ;
      LAYER met2 ;
        RECT 2108.200 1700.410 2108.480 1704.000 ;
        RECT 2105.580 1700.270 2108.480 1700.410 ;
        RECT 2105.580 30.930 2105.720 1700.270 ;
        RECT 2108.200 1700.000 2108.480 1700.270 ;
        RECT 1864.480 30.610 1864.740 30.930 ;
        RECT 2105.520 30.610 2105.780 30.930 ;
        RECT 1864.540 22.170 1864.680 30.610 ;
        RECT 1864.080 22.030 1864.680 22.170 ;
        RECT 1864.080 2.400 1864.220 22.030 ;
        RECT 1863.870 -4.800 1864.430 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1525.965 1449.165 1526.135 1497.275 ;
        RECT 1525.965 1352.605 1526.135 1400.715 ;
        RECT 1525.965 1256.045 1526.135 1304.155 ;
        RECT 1525.505 669.545 1525.675 717.655 ;
        RECT 1524.585 620.925 1524.755 628.575 ;
        RECT 1525.505 531.505 1525.675 579.615 ;
        RECT 1525.965 386.325 1526.135 434.775 ;
        RECT 1525.965 338.045 1526.135 352.495 ;
        RECT 1525.505 67.065 1525.675 96.475 ;
      LAYER mcon ;
        RECT 1525.965 1497.105 1526.135 1497.275 ;
        RECT 1525.965 1400.545 1526.135 1400.715 ;
        RECT 1525.965 1303.985 1526.135 1304.155 ;
        RECT 1525.505 717.485 1525.675 717.655 ;
        RECT 1524.585 628.405 1524.755 628.575 ;
        RECT 1525.505 579.445 1525.675 579.615 ;
        RECT 1525.965 434.605 1526.135 434.775 ;
        RECT 1525.965 352.325 1526.135 352.495 ;
        RECT 1525.505 96.305 1525.675 96.475 ;
      LAYER met1 ;
        RECT 1525.890 1655.840 1526.210 1656.100 ;
        RECT 1525.980 1655.700 1526.120 1655.840 ;
        RECT 1526.350 1655.700 1526.670 1655.760 ;
        RECT 1525.980 1655.560 1526.670 1655.700 ;
        RECT 1526.350 1655.500 1526.670 1655.560 ;
        RECT 1525.890 1545.880 1526.210 1545.940 ;
        RECT 1526.350 1545.880 1526.670 1545.940 ;
        RECT 1525.890 1545.740 1526.670 1545.880 ;
        RECT 1525.890 1545.680 1526.210 1545.740 ;
        RECT 1526.350 1545.680 1526.670 1545.740 ;
        RECT 1525.890 1497.260 1526.210 1497.320 ;
        RECT 1525.695 1497.120 1526.210 1497.260 ;
        RECT 1525.890 1497.060 1526.210 1497.120 ;
        RECT 1525.890 1449.320 1526.210 1449.380 ;
        RECT 1525.695 1449.180 1526.210 1449.320 ;
        RECT 1525.890 1449.120 1526.210 1449.180 ;
        RECT 1525.890 1400.700 1526.210 1400.760 ;
        RECT 1525.695 1400.560 1526.210 1400.700 ;
        RECT 1525.890 1400.500 1526.210 1400.560 ;
        RECT 1525.890 1352.760 1526.210 1352.820 ;
        RECT 1525.695 1352.620 1526.210 1352.760 ;
        RECT 1525.890 1352.560 1526.210 1352.620 ;
        RECT 1525.890 1304.140 1526.210 1304.200 ;
        RECT 1525.695 1304.000 1526.210 1304.140 ;
        RECT 1525.890 1303.940 1526.210 1304.000 ;
        RECT 1525.890 1256.200 1526.210 1256.260 ;
        RECT 1525.695 1256.060 1526.210 1256.200 ;
        RECT 1525.890 1256.000 1526.210 1256.060 ;
        RECT 1525.890 1159.300 1526.210 1159.360 ;
        RECT 1526.810 1159.300 1527.130 1159.360 ;
        RECT 1525.890 1159.160 1527.130 1159.300 ;
        RECT 1525.890 1159.100 1526.210 1159.160 ;
        RECT 1526.810 1159.100 1527.130 1159.160 ;
        RECT 1525.890 1062.740 1526.210 1062.800 ;
        RECT 1526.810 1062.740 1527.130 1062.800 ;
        RECT 1525.890 1062.600 1527.130 1062.740 ;
        RECT 1525.890 1062.540 1526.210 1062.600 ;
        RECT 1526.810 1062.540 1527.130 1062.600 ;
        RECT 1525.890 966.180 1526.210 966.240 ;
        RECT 1526.810 966.180 1527.130 966.240 ;
        RECT 1525.890 966.040 1527.130 966.180 ;
        RECT 1525.890 965.980 1526.210 966.040 ;
        RECT 1526.810 965.980 1527.130 966.040 ;
        RECT 1525.430 717.640 1525.750 717.700 ;
        RECT 1525.235 717.500 1525.750 717.640 ;
        RECT 1525.430 717.440 1525.750 717.500 ;
        RECT 1525.430 669.700 1525.750 669.760 ;
        RECT 1525.235 669.560 1525.750 669.700 ;
        RECT 1525.430 669.500 1525.750 669.560 ;
        RECT 1524.525 628.560 1524.815 628.605 ;
        RECT 1525.430 628.560 1525.750 628.620 ;
        RECT 1524.525 628.420 1525.750 628.560 ;
        RECT 1524.525 628.375 1524.815 628.420 ;
        RECT 1525.430 628.360 1525.750 628.420 ;
        RECT 1524.510 621.080 1524.830 621.140 ;
        RECT 1524.315 620.940 1524.830 621.080 ;
        RECT 1524.510 620.880 1524.830 620.940 ;
        RECT 1525.430 579.600 1525.750 579.660 ;
        RECT 1525.235 579.460 1525.750 579.600 ;
        RECT 1525.430 579.400 1525.750 579.460 ;
        RECT 1525.445 531.660 1525.735 531.705 ;
        RECT 1525.890 531.660 1526.210 531.720 ;
        RECT 1525.445 531.520 1526.210 531.660 ;
        RECT 1525.445 531.475 1525.735 531.520 ;
        RECT 1525.890 531.460 1526.210 531.520 ;
        RECT 1525.890 434.760 1526.210 434.820 ;
        RECT 1525.695 434.620 1526.210 434.760 ;
        RECT 1525.890 434.560 1526.210 434.620 ;
        RECT 1525.890 386.480 1526.210 386.540 ;
        RECT 1525.695 386.340 1526.210 386.480 ;
        RECT 1525.890 386.280 1526.210 386.340 ;
        RECT 1525.890 352.480 1526.210 352.540 ;
        RECT 1525.695 352.340 1526.210 352.480 ;
        RECT 1525.890 352.280 1526.210 352.340 ;
        RECT 1525.890 338.200 1526.210 338.260 ;
        RECT 1525.695 338.060 1526.210 338.200 ;
        RECT 1525.890 338.000 1526.210 338.060 ;
        RECT 1525.890 255.920 1526.210 255.980 ;
        RECT 1525.520 255.780 1526.210 255.920 ;
        RECT 1525.520 255.300 1525.660 255.780 ;
        RECT 1525.890 255.720 1526.210 255.780 ;
        RECT 1525.430 255.040 1525.750 255.300 ;
        RECT 1525.430 96.460 1525.750 96.520 ;
        RECT 1525.235 96.320 1525.750 96.460 ;
        RECT 1525.430 96.260 1525.750 96.320 ;
        RECT 744.810 67.220 745.130 67.280 ;
        RECT 1525.445 67.220 1525.735 67.265 ;
        RECT 744.810 67.080 1525.735 67.220 ;
        RECT 744.810 67.020 745.130 67.080 ;
        RECT 1525.445 67.035 1525.735 67.080 ;
      LAYER via ;
        RECT 1525.920 1655.840 1526.180 1656.100 ;
        RECT 1526.380 1655.500 1526.640 1655.760 ;
        RECT 1525.920 1545.680 1526.180 1545.940 ;
        RECT 1526.380 1545.680 1526.640 1545.940 ;
        RECT 1525.920 1497.060 1526.180 1497.320 ;
        RECT 1525.920 1449.120 1526.180 1449.380 ;
        RECT 1525.920 1400.500 1526.180 1400.760 ;
        RECT 1525.920 1352.560 1526.180 1352.820 ;
        RECT 1525.920 1303.940 1526.180 1304.200 ;
        RECT 1525.920 1256.000 1526.180 1256.260 ;
        RECT 1525.920 1159.100 1526.180 1159.360 ;
        RECT 1526.840 1159.100 1527.100 1159.360 ;
        RECT 1525.920 1062.540 1526.180 1062.800 ;
        RECT 1526.840 1062.540 1527.100 1062.800 ;
        RECT 1525.920 965.980 1526.180 966.240 ;
        RECT 1526.840 965.980 1527.100 966.240 ;
        RECT 1525.460 717.440 1525.720 717.700 ;
        RECT 1525.460 669.500 1525.720 669.760 ;
        RECT 1525.460 628.360 1525.720 628.620 ;
        RECT 1524.540 620.880 1524.800 621.140 ;
        RECT 1525.460 579.400 1525.720 579.660 ;
        RECT 1525.920 531.460 1526.180 531.720 ;
        RECT 1525.920 434.560 1526.180 434.820 ;
        RECT 1525.920 386.280 1526.180 386.540 ;
        RECT 1525.920 352.280 1526.180 352.540 ;
        RECT 1525.920 338.000 1526.180 338.260 ;
        RECT 1525.920 255.720 1526.180 255.980 ;
        RECT 1525.460 255.040 1525.720 255.300 ;
        RECT 1525.460 96.260 1525.720 96.520 ;
        RECT 744.840 67.020 745.100 67.280 ;
      LAYER met2 ;
        RECT 1529.520 1700.410 1529.800 1704.000 ;
        RECT 1526.900 1700.270 1529.800 1700.410 ;
        RECT 1526.900 1677.970 1527.040 1700.270 ;
        RECT 1529.520 1700.000 1529.800 1700.270 ;
        RECT 1525.980 1677.830 1527.040 1677.970 ;
        RECT 1525.980 1656.130 1526.120 1677.830 ;
        RECT 1525.920 1655.810 1526.180 1656.130 ;
        RECT 1526.380 1655.470 1526.640 1655.790 ;
        RECT 1526.440 1545.970 1526.580 1655.470 ;
        RECT 1525.920 1545.650 1526.180 1545.970 ;
        RECT 1526.380 1545.650 1526.640 1545.970 ;
        RECT 1525.980 1497.350 1526.120 1545.650 ;
        RECT 1525.920 1497.030 1526.180 1497.350 ;
        RECT 1525.920 1449.090 1526.180 1449.410 ;
        RECT 1525.980 1400.790 1526.120 1449.090 ;
        RECT 1525.920 1400.470 1526.180 1400.790 ;
        RECT 1525.920 1352.530 1526.180 1352.850 ;
        RECT 1525.980 1304.230 1526.120 1352.530 ;
        RECT 1525.920 1303.910 1526.180 1304.230 ;
        RECT 1525.920 1255.970 1526.180 1256.290 ;
        RECT 1525.980 1207.525 1526.120 1255.970 ;
        RECT 1525.910 1207.155 1526.190 1207.525 ;
        RECT 1526.830 1207.155 1527.110 1207.525 ;
        RECT 1526.900 1159.390 1527.040 1207.155 ;
        RECT 1525.920 1159.070 1526.180 1159.390 ;
        RECT 1526.840 1159.070 1527.100 1159.390 ;
        RECT 1525.980 1110.965 1526.120 1159.070 ;
        RECT 1525.910 1110.595 1526.190 1110.965 ;
        RECT 1526.830 1110.595 1527.110 1110.965 ;
        RECT 1526.900 1062.830 1527.040 1110.595 ;
        RECT 1525.920 1062.510 1526.180 1062.830 ;
        RECT 1526.840 1062.510 1527.100 1062.830 ;
        RECT 1525.980 1014.405 1526.120 1062.510 ;
        RECT 1525.910 1014.035 1526.190 1014.405 ;
        RECT 1526.830 1014.035 1527.110 1014.405 ;
        RECT 1526.900 966.270 1527.040 1014.035 ;
        RECT 1525.920 965.950 1526.180 966.270 ;
        RECT 1526.840 965.950 1527.100 966.270 ;
        RECT 1525.980 835.450 1526.120 965.950 ;
        RECT 1525.520 835.310 1526.120 835.450 ;
        RECT 1525.520 834.770 1525.660 835.310 ;
        RECT 1525.520 834.630 1526.120 834.770 ;
        RECT 1525.980 773.685 1526.120 834.630 ;
        RECT 1525.910 773.315 1526.190 773.685 ;
        RECT 1525.910 772.635 1526.190 773.005 ;
        RECT 1525.980 738.890 1526.120 772.635 ;
        RECT 1525.980 738.750 1526.580 738.890 ;
        RECT 1526.440 725.405 1526.580 738.750 ;
        RECT 1526.370 725.035 1526.650 725.405 ;
        RECT 1525.450 724.355 1525.730 724.725 ;
        RECT 1525.520 717.730 1525.660 724.355 ;
        RECT 1525.460 717.410 1525.720 717.730 ;
        RECT 1525.460 669.470 1525.720 669.790 ;
        RECT 1525.520 628.650 1525.660 669.470 ;
        RECT 1525.460 628.330 1525.720 628.650 ;
        RECT 1524.540 620.850 1524.800 621.170 ;
        RECT 1524.600 579.885 1524.740 620.850 ;
        RECT 1524.530 579.515 1524.810 579.885 ;
        RECT 1525.450 579.515 1525.730 579.885 ;
        RECT 1525.460 579.370 1525.720 579.515 ;
        RECT 1525.920 531.435 1526.180 531.750 ;
        RECT 1525.910 531.065 1526.190 531.435 ;
        RECT 1526.370 529.875 1526.650 530.245 ;
        RECT 1526.440 496.130 1526.580 529.875 ;
        RECT 1525.980 495.990 1526.580 496.130 ;
        RECT 1525.980 434.850 1526.120 495.990 ;
        RECT 1525.920 434.530 1526.180 434.850 ;
        RECT 1525.920 386.250 1526.180 386.570 ;
        RECT 1525.980 352.570 1526.120 386.250 ;
        RECT 1525.920 352.250 1526.180 352.570 ;
        RECT 1525.920 337.970 1526.180 338.290 ;
        RECT 1525.980 256.010 1526.120 337.970 ;
        RECT 1525.920 255.690 1526.180 256.010 ;
        RECT 1525.460 255.010 1525.720 255.330 ;
        RECT 1525.520 96.550 1525.660 255.010 ;
        RECT 1525.460 96.230 1525.720 96.550 ;
        RECT 744.840 66.990 745.100 67.310 ;
        RECT 744.900 16.730 745.040 66.990 ;
        RECT 740.300 16.590 745.040 16.730 ;
        RECT 740.300 2.400 740.440 16.590 ;
        RECT 740.090 -4.800 740.650 2.400 ;
      LAYER via2 ;
        RECT 1525.910 1207.200 1526.190 1207.480 ;
        RECT 1526.830 1207.200 1527.110 1207.480 ;
        RECT 1525.910 1110.640 1526.190 1110.920 ;
        RECT 1526.830 1110.640 1527.110 1110.920 ;
        RECT 1525.910 1014.080 1526.190 1014.360 ;
        RECT 1526.830 1014.080 1527.110 1014.360 ;
        RECT 1525.910 773.360 1526.190 773.640 ;
        RECT 1525.910 772.680 1526.190 772.960 ;
        RECT 1526.370 725.080 1526.650 725.360 ;
        RECT 1525.450 724.400 1525.730 724.680 ;
        RECT 1524.530 579.560 1524.810 579.840 ;
        RECT 1525.450 579.560 1525.730 579.840 ;
        RECT 1525.910 531.110 1526.190 531.390 ;
        RECT 1526.370 529.920 1526.650 530.200 ;
      LAYER met3 ;
        RECT 1525.885 1207.490 1526.215 1207.505 ;
        RECT 1526.805 1207.490 1527.135 1207.505 ;
        RECT 1525.885 1207.190 1527.135 1207.490 ;
        RECT 1525.885 1207.175 1526.215 1207.190 ;
        RECT 1526.805 1207.175 1527.135 1207.190 ;
        RECT 1525.885 1110.930 1526.215 1110.945 ;
        RECT 1526.805 1110.930 1527.135 1110.945 ;
        RECT 1525.885 1110.630 1527.135 1110.930 ;
        RECT 1525.885 1110.615 1526.215 1110.630 ;
        RECT 1526.805 1110.615 1527.135 1110.630 ;
        RECT 1525.885 1014.370 1526.215 1014.385 ;
        RECT 1526.805 1014.370 1527.135 1014.385 ;
        RECT 1525.885 1014.070 1527.135 1014.370 ;
        RECT 1525.885 1014.055 1526.215 1014.070 ;
        RECT 1526.805 1014.055 1527.135 1014.070 ;
        RECT 1525.885 773.650 1526.215 773.665 ;
        RECT 1525.885 773.350 1526.890 773.650 ;
        RECT 1525.885 773.335 1526.215 773.350 ;
        RECT 1525.885 772.970 1526.215 772.985 ;
        RECT 1526.590 772.970 1526.890 773.350 ;
        RECT 1525.885 772.670 1526.890 772.970 ;
        RECT 1525.885 772.655 1526.215 772.670 ;
        RECT 1526.345 725.370 1526.675 725.385 ;
        RECT 1524.750 725.070 1526.675 725.370 ;
        RECT 1524.750 724.690 1525.050 725.070 ;
        RECT 1526.345 725.055 1526.675 725.070 ;
        RECT 1525.425 724.690 1525.755 724.705 ;
        RECT 1524.750 724.390 1525.755 724.690 ;
        RECT 1525.425 724.375 1525.755 724.390 ;
        RECT 1524.505 579.850 1524.835 579.865 ;
        RECT 1525.425 579.850 1525.755 579.865 ;
        RECT 1524.505 579.550 1525.755 579.850 ;
        RECT 1524.505 579.535 1524.835 579.550 ;
        RECT 1525.425 579.535 1525.755 579.550 ;
        RECT 1525.885 531.400 1526.215 531.415 ;
        RECT 1525.885 531.100 1526.890 531.400 ;
        RECT 1525.885 531.085 1526.215 531.100 ;
        RECT 1526.590 530.225 1526.890 531.100 ;
        RECT 1526.345 529.910 1526.890 530.225 ;
        RECT 1526.345 529.895 1526.675 529.910 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2112.005 1594.005 2112.175 1642.115 ;
        RECT 2112.465 1499.485 2112.635 1545.555 ;
        RECT 2112.005 786.505 2112.175 821.015 ;
        RECT 2112.005 689.605 2112.175 724.455 ;
        RECT 2112.005 496.485 2112.175 531.335 ;
        RECT 2112.005 386.325 2112.175 434.775 ;
      LAYER mcon ;
        RECT 2112.005 1641.945 2112.175 1642.115 ;
        RECT 2112.465 1545.385 2112.635 1545.555 ;
        RECT 2112.005 820.845 2112.175 821.015 ;
        RECT 2112.005 724.285 2112.175 724.455 ;
        RECT 2112.005 531.165 2112.175 531.335 ;
        RECT 2112.005 434.605 2112.175 434.775 ;
      LAYER met1 ;
        RECT 2111.470 1678.140 2111.790 1678.200 ;
        RECT 2116.070 1678.140 2116.390 1678.200 ;
        RECT 2111.470 1678.000 2116.390 1678.140 ;
        RECT 2111.470 1677.940 2111.790 1678.000 ;
        RECT 2116.070 1677.940 2116.390 1678.000 ;
        RECT 2111.470 1656.040 2111.790 1656.100 ;
        RECT 2112.390 1656.040 2112.710 1656.100 ;
        RECT 2111.470 1655.900 2112.710 1656.040 ;
        RECT 2111.470 1655.840 2111.790 1655.900 ;
        RECT 2112.390 1655.840 2112.710 1655.900 ;
        RECT 2111.945 1642.100 2112.235 1642.145 ;
        RECT 2112.390 1642.100 2112.710 1642.160 ;
        RECT 2111.945 1641.960 2112.710 1642.100 ;
        RECT 2111.945 1641.915 2112.235 1641.960 ;
        RECT 2112.390 1641.900 2112.710 1641.960 ;
        RECT 2111.930 1594.160 2112.250 1594.220 ;
        RECT 2111.735 1594.020 2112.250 1594.160 ;
        RECT 2111.930 1593.960 2112.250 1594.020 ;
        RECT 2111.470 1559.140 2111.790 1559.200 ;
        RECT 2112.390 1559.140 2112.710 1559.200 ;
        RECT 2111.470 1559.000 2112.710 1559.140 ;
        RECT 2111.470 1558.940 2111.790 1559.000 ;
        RECT 2112.390 1558.940 2112.710 1559.000 ;
        RECT 2112.390 1545.540 2112.710 1545.600 ;
        RECT 2112.195 1545.400 2112.710 1545.540 ;
        RECT 2112.390 1545.340 2112.710 1545.400 ;
        RECT 2112.390 1499.640 2112.710 1499.700 ;
        RECT 2112.195 1499.500 2112.710 1499.640 ;
        RECT 2112.390 1499.440 2112.710 1499.500 ;
        RECT 2111.470 1414.640 2111.790 1414.700 ;
        RECT 2112.390 1414.640 2112.710 1414.700 ;
        RECT 2111.470 1414.500 2112.710 1414.640 ;
        RECT 2111.470 1414.440 2111.790 1414.500 ;
        RECT 2112.390 1414.440 2112.710 1414.500 ;
        RECT 2111.470 1318.080 2111.790 1318.140 ;
        RECT 2112.390 1318.080 2112.710 1318.140 ;
        RECT 2111.470 1317.940 2112.710 1318.080 ;
        RECT 2111.470 1317.880 2111.790 1317.940 ;
        RECT 2112.390 1317.880 2112.710 1317.940 ;
        RECT 2111.470 1221.520 2111.790 1221.580 ;
        RECT 2112.390 1221.520 2112.710 1221.580 ;
        RECT 2111.470 1221.380 2112.710 1221.520 ;
        RECT 2111.470 1221.320 2111.790 1221.380 ;
        RECT 2112.390 1221.320 2112.710 1221.380 ;
        RECT 2111.470 1124.960 2111.790 1125.020 ;
        RECT 2112.390 1124.960 2112.710 1125.020 ;
        RECT 2111.470 1124.820 2112.710 1124.960 ;
        RECT 2111.470 1124.760 2111.790 1124.820 ;
        RECT 2112.390 1124.760 2112.710 1124.820 ;
        RECT 2111.470 1028.400 2111.790 1028.460 ;
        RECT 2112.390 1028.400 2112.710 1028.460 ;
        RECT 2111.470 1028.260 2112.710 1028.400 ;
        RECT 2111.470 1028.200 2111.790 1028.260 ;
        RECT 2112.390 1028.200 2112.710 1028.260 ;
        RECT 2111.470 931.840 2111.790 931.900 ;
        RECT 2112.390 931.840 2112.710 931.900 ;
        RECT 2111.470 931.700 2112.710 931.840 ;
        RECT 2111.470 931.640 2111.790 931.700 ;
        RECT 2112.390 931.640 2112.710 931.700 ;
        RECT 2112.390 869.620 2112.710 869.680 ;
        RECT 2113.310 869.620 2113.630 869.680 ;
        RECT 2112.390 869.480 2113.630 869.620 ;
        RECT 2112.390 869.420 2112.710 869.480 ;
        RECT 2113.310 869.420 2113.630 869.480 ;
        RECT 2111.470 835.280 2111.790 835.340 ;
        RECT 2112.390 835.280 2112.710 835.340 ;
        RECT 2111.470 835.140 2112.710 835.280 ;
        RECT 2111.470 835.080 2111.790 835.140 ;
        RECT 2112.390 835.080 2112.710 835.140 ;
        RECT 2111.930 821.000 2112.250 821.060 ;
        RECT 2111.735 820.860 2112.250 821.000 ;
        RECT 2111.930 820.800 2112.250 820.860 ;
        RECT 2111.930 786.660 2112.250 786.720 ;
        RECT 2111.735 786.520 2112.250 786.660 ;
        RECT 2111.930 786.460 2112.250 786.520 ;
        RECT 2111.470 738.380 2111.790 738.440 ;
        RECT 2112.390 738.380 2112.710 738.440 ;
        RECT 2111.470 738.240 2112.710 738.380 ;
        RECT 2111.470 738.180 2111.790 738.240 ;
        RECT 2112.390 738.180 2112.710 738.240 ;
        RECT 2111.930 724.440 2112.250 724.500 ;
        RECT 2111.735 724.300 2112.250 724.440 ;
        RECT 2111.930 724.240 2112.250 724.300 ;
        RECT 2111.930 689.760 2112.250 689.820 ;
        RECT 2111.735 689.620 2112.250 689.760 ;
        RECT 2111.930 689.560 2112.250 689.620 ;
        RECT 2111.470 641.820 2111.790 641.880 ;
        RECT 2112.390 641.820 2112.710 641.880 ;
        RECT 2111.470 641.680 2112.710 641.820 ;
        RECT 2111.470 641.620 2111.790 641.680 ;
        RECT 2112.390 641.620 2112.710 641.680 ;
        RECT 2111.930 593.340 2112.250 593.600 ;
        RECT 2112.020 593.200 2112.160 593.340 ;
        RECT 2112.390 593.200 2112.710 593.260 ;
        RECT 2112.020 593.060 2112.710 593.200 ;
        RECT 2112.390 593.000 2112.710 593.060 ;
        RECT 2111.470 545.260 2111.790 545.320 ;
        RECT 2112.390 545.260 2112.710 545.320 ;
        RECT 2111.470 545.120 2112.710 545.260 ;
        RECT 2111.470 545.060 2111.790 545.120 ;
        RECT 2112.390 545.060 2112.710 545.120 ;
        RECT 2111.930 531.320 2112.250 531.380 ;
        RECT 2111.735 531.180 2112.250 531.320 ;
        RECT 2111.930 531.120 2112.250 531.180 ;
        RECT 2111.930 496.640 2112.250 496.700 ;
        RECT 2111.735 496.500 2112.250 496.640 ;
        RECT 2111.930 496.440 2112.250 496.500 ;
        RECT 2111.470 448.700 2111.790 448.760 ;
        RECT 2112.390 448.700 2112.710 448.760 ;
        RECT 2111.470 448.560 2112.710 448.700 ;
        RECT 2111.470 448.500 2111.790 448.560 ;
        RECT 2112.390 448.500 2112.710 448.560 ;
        RECT 2111.930 434.760 2112.250 434.820 ;
        RECT 2111.735 434.620 2112.250 434.760 ;
        RECT 2111.930 434.560 2112.250 434.620 ;
        RECT 2111.945 386.480 2112.235 386.525 ;
        RECT 2112.390 386.480 2112.710 386.540 ;
        RECT 2111.945 386.340 2112.710 386.480 ;
        RECT 2111.945 386.295 2112.235 386.340 ;
        RECT 2112.390 386.280 2112.710 386.340 ;
        RECT 2111.930 338.200 2112.250 338.260 ;
        RECT 2112.390 338.200 2112.710 338.260 ;
        RECT 2111.930 338.060 2112.710 338.200 ;
        RECT 2111.930 338.000 2112.250 338.060 ;
        RECT 2112.390 338.000 2112.710 338.060 ;
        RECT 2111.930 241.640 2112.250 241.700 ;
        RECT 2112.390 241.640 2112.710 241.700 ;
        RECT 2111.930 241.500 2112.710 241.640 ;
        RECT 2111.930 241.440 2112.250 241.500 ;
        RECT 2112.390 241.440 2112.710 241.500 ;
        RECT 2111.930 138.280 2112.250 138.340 ;
        RECT 2112.390 138.280 2112.710 138.340 ;
        RECT 2111.930 138.140 2112.710 138.280 ;
        RECT 2111.930 138.080 2112.250 138.140 ;
        RECT 2112.390 138.080 2112.710 138.140 ;
        RECT 2110.550 112.780 2110.870 112.840 ;
        RECT 2111.930 112.780 2112.250 112.840 ;
        RECT 2110.550 112.640 2112.250 112.780 ;
        RECT 2110.550 112.580 2110.870 112.640 ;
        RECT 2111.930 112.580 2112.250 112.640 ;
        RECT 2110.550 48.520 2110.870 48.580 ;
        RECT 2111.930 48.520 2112.250 48.580 ;
        RECT 2110.550 48.380 2112.250 48.520 ;
        RECT 2110.550 48.320 2110.870 48.380 ;
        RECT 2111.930 48.320 2112.250 48.380 ;
        RECT 1881.930 25.400 1882.250 25.460 ;
        RECT 2111.930 25.400 2112.250 25.460 ;
        RECT 1881.930 25.260 2112.250 25.400 ;
        RECT 1881.930 25.200 1882.250 25.260 ;
        RECT 2111.930 25.200 2112.250 25.260 ;
      LAYER via ;
        RECT 2111.500 1677.940 2111.760 1678.200 ;
        RECT 2116.100 1677.940 2116.360 1678.200 ;
        RECT 2111.500 1655.840 2111.760 1656.100 ;
        RECT 2112.420 1655.840 2112.680 1656.100 ;
        RECT 2112.420 1641.900 2112.680 1642.160 ;
        RECT 2111.960 1593.960 2112.220 1594.220 ;
        RECT 2111.500 1558.940 2111.760 1559.200 ;
        RECT 2112.420 1558.940 2112.680 1559.200 ;
        RECT 2112.420 1545.340 2112.680 1545.600 ;
        RECT 2112.420 1499.440 2112.680 1499.700 ;
        RECT 2111.500 1414.440 2111.760 1414.700 ;
        RECT 2112.420 1414.440 2112.680 1414.700 ;
        RECT 2111.500 1317.880 2111.760 1318.140 ;
        RECT 2112.420 1317.880 2112.680 1318.140 ;
        RECT 2111.500 1221.320 2111.760 1221.580 ;
        RECT 2112.420 1221.320 2112.680 1221.580 ;
        RECT 2111.500 1124.760 2111.760 1125.020 ;
        RECT 2112.420 1124.760 2112.680 1125.020 ;
        RECT 2111.500 1028.200 2111.760 1028.460 ;
        RECT 2112.420 1028.200 2112.680 1028.460 ;
        RECT 2111.500 931.640 2111.760 931.900 ;
        RECT 2112.420 931.640 2112.680 931.900 ;
        RECT 2112.420 869.420 2112.680 869.680 ;
        RECT 2113.340 869.420 2113.600 869.680 ;
        RECT 2111.500 835.080 2111.760 835.340 ;
        RECT 2112.420 835.080 2112.680 835.340 ;
        RECT 2111.960 820.800 2112.220 821.060 ;
        RECT 2111.960 786.460 2112.220 786.720 ;
        RECT 2111.500 738.180 2111.760 738.440 ;
        RECT 2112.420 738.180 2112.680 738.440 ;
        RECT 2111.960 724.240 2112.220 724.500 ;
        RECT 2111.960 689.560 2112.220 689.820 ;
        RECT 2111.500 641.620 2111.760 641.880 ;
        RECT 2112.420 641.620 2112.680 641.880 ;
        RECT 2111.960 593.340 2112.220 593.600 ;
        RECT 2112.420 593.000 2112.680 593.260 ;
        RECT 2111.500 545.060 2111.760 545.320 ;
        RECT 2112.420 545.060 2112.680 545.320 ;
        RECT 2111.960 531.120 2112.220 531.380 ;
        RECT 2111.960 496.440 2112.220 496.700 ;
        RECT 2111.500 448.500 2111.760 448.760 ;
        RECT 2112.420 448.500 2112.680 448.760 ;
        RECT 2111.960 434.560 2112.220 434.820 ;
        RECT 2112.420 386.280 2112.680 386.540 ;
        RECT 2111.960 338.000 2112.220 338.260 ;
        RECT 2112.420 338.000 2112.680 338.260 ;
        RECT 2111.960 241.440 2112.220 241.700 ;
        RECT 2112.420 241.440 2112.680 241.700 ;
        RECT 2111.960 138.080 2112.220 138.340 ;
        RECT 2112.420 138.080 2112.680 138.340 ;
        RECT 2110.580 112.580 2110.840 112.840 ;
        RECT 2111.960 112.580 2112.220 112.840 ;
        RECT 2110.580 48.320 2110.840 48.580 ;
        RECT 2111.960 48.320 2112.220 48.580 ;
        RECT 1881.960 25.200 1882.220 25.460 ;
        RECT 2111.960 25.200 2112.220 25.460 ;
      LAYER met2 ;
        RECT 2117.400 1700.410 2117.680 1704.000 ;
        RECT 2116.160 1700.270 2117.680 1700.410 ;
        RECT 2116.160 1678.230 2116.300 1700.270 ;
        RECT 2117.400 1700.000 2117.680 1700.270 ;
        RECT 2111.500 1677.910 2111.760 1678.230 ;
        RECT 2116.100 1677.910 2116.360 1678.230 ;
        RECT 2111.560 1656.130 2111.700 1677.910 ;
        RECT 2111.500 1655.810 2111.760 1656.130 ;
        RECT 2112.420 1655.810 2112.680 1656.130 ;
        RECT 2112.480 1642.190 2112.620 1655.810 ;
        RECT 2112.420 1641.870 2112.680 1642.190 ;
        RECT 2111.960 1593.930 2112.220 1594.250 ;
        RECT 2112.020 1559.650 2112.160 1593.930 ;
        RECT 2111.560 1559.510 2112.160 1559.650 ;
        RECT 2111.560 1559.230 2111.700 1559.510 ;
        RECT 2111.500 1558.910 2111.760 1559.230 ;
        RECT 2112.420 1558.910 2112.680 1559.230 ;
        RECT 2112.480 1545.630 2112.620 1558.910 ;
        RECT 2112.420 1545.310 2112.680 1545.630 ;
        RECT 2112.420 1499.410 2112.680 1499.730 ;
        RECT 2112.480 1414.730 2112.620 1499.410 ;
        RECT 2111.500 1414.410 2111.760 1414.730 ;
        RECT 2112.420 1414.410 2112.680 1414.730 ;
        RECT 2111.560 1414.130 2111.700 1414.410 ;
        RECT 2111.560 1413.990 2112.160 1414.130 ;
        RECT 2112.020 1366.530 2112.160 1413.990 ;
        RECT 2112.020 1366.390 2112.620 1366.530 ;
        RECT 2112.480 1318.170 2112.620 1366.390 ;
        RECT 2111.500 1317.850 2111.760 1318.170 ;
        RECT 2112.420 1317.850 2112.680 1318.170 ;
        RECT 2111.560 1317.570 2111.700 1317.850 ;
        RECT 2111.560 1317.430 2112.160 1317.570 ;
        RECT 2112.020 1269.970 2112.160 1317.430 ;
        RECT 2112.020 1269.830 2112.620 1269.970 ;
        RECT 2112.480 1221.610 2112.620 1269.830 ;
        RECT 2111.500 1221.290 2111.760 1221.610 ;
        RECT 2112.420 1221.290 2112.680 1221.610 ;
        RECT 2111.560 1221.010 2111.700 1221.290 ;
        RECT 2111.560 1220.870 2112.160 1221.010 ;
        RECT 2112.020 1173.410 2112.160 1220.870 ;
        RECT 2112.020 1173.270 2112.620 1173.410 ;
        RECT 2112.480 1125.050 2112.620 1173.270 ;
        RECT 2111.500 1124.730 2111.760 1125.050 ;
        RECT 2112.420 1124.730 2112.680 1125.050 ;
        RECT 2111.560 1124.450 2111.700 1124.730 ;
        RECT 2111.560 1124.310 2112.160 1124.450 ;
        RECT 2112.020 1076.850 2112.160 1124.310 ;
        RECT 2112.020 1076.710 2112.620 1076.850 ;
        RECT 2112.480 1028.490 2112.620 1076.710 ;
        RECT 2111.500 1028.170 2111.760 1028.490 ;
        RECT 2112.420 1028.170 2112.680 1028.490 ;
        RECT 2111.560 1027.890 2111.700 1028.170 ;
        RECT 2111.560 1027.750 2112.160 1027.890 ;
        RECT 2112.020 980.290 2112.160 1027.750 ;
        RECT 2112.020 980.150 2112.620 980.290 ;
        RECT 2112.480 931.930 2112.620 980.150 ;
        RECT 2111.500 931.610 2111.760 931.930 ;
        RECT 2112.420 931.610 2112.680 931.930 ;
        RECT 2111.560 931.330 2111.700 931.610 ;
        RECT 2111.560 931.190 2112.160 931.330 ;
        RECT 2112.020 917.845 2112.160 931.190 ;
        RECT 2111.950 917.475 2112.230 917.845 ;
        RECT 2113.330 917.475 2113.610 917.845 ;
        RECT 2113.400 869.710 2113.540 917.475 ;
        RECT 2112.420 869.390 2112.680 869.710 ;
        RECT 2113.340 869.390 2113.600 869.710 ;
        RECT 2112.480 835.370 2112.620 869.390 ;
        RECT 2111.500 835.050 2111.760 835.370 ;
        RECT 2112.420 835.050 2112.680 835.370 ;
        RECT 2111.560 834.770 2111.700 835.050 ;
        RECT 2111.560 834.630 2112.160 834.770 ;
        RECT 2112.020 821.090 2112.160 834.630 ;
        RECT 2111.960 820.770 2112.220 821.090 ;
        RECT 2111.960 786.430 2112.220 786.750 ;
        RECT 2112.020 772.890 2112.160 786.430 ;
        RECT 2112.020 772.750 2112.620 772.890 ;
        RECT 2112.480 738.470 2112.620 772.750 ;
        RECT 2111.500 738.210 2111.760 738.470 ;
        RECT 2111.500 738.150 2112.160 738.210 ;
        RECT 2112.420 738.150 2112.680 738.470 ;
        RECT 2111.560 738.070 2112.160 738.150 ;
        RECT 2112.020 724.530 2112.160 738.070 ;
        RECT 2111.960 724.210 2112.220 724.530 ;
        RECT 2111.960 689.530 2112.220 689.850 ;
        RECT 2112.020 676.330 2112.160 689.530 ;
        RECT 2112.020 676.190 2112.620 676.330 ;
        RECT 2112.480 641.910 2112.620 676.190 ;
        RECT 2111.500 641.650 2111.760 641.910 ;
        RECT 2111.500 641.590 2112.160 641.650 ;
        RECT 2112.420 641.590 2112.680 641.910 ;
        RECT 2111.560 641.510 2112.160 641.590 ;
        RECT 2112.020 593.630 2112.160 641.510 ;
        RECT 2111.960 593.310 2112.220 593.630 ;
        RECT 2112.420 592.970 2112.680 593.290 ;
        RECT 2112.480 545.350 2112.620 592.970 ;
        RECT 2111.500 545.090 2111.760 545.350 ;
        RECT 2111.500 545.030 2112.160 545.090 ;
        RECT 2112.420 545.030 2112.680 545.350 ;
        RECT 2111.560 544.950 2112.160 545.030 ;
        RECT 2112.020 531.410 2112.160 544.950 ;
        RECT 2111.960 531.090 2112.220 531.410 ;
        RECT 2111.960 496.410 2112.220 496.730 ;
        RECT 2112.020 483.210 2112.160 496.410 ;
        RECT 2112.020 483.070 2112.620 483.210 ;
        RECT 2112.480 448.790 2112.620 483.070 ;
        RECT 2111.500 448.530 2111.760 448.790 ;
        RECT 2111.500 448.470 2112.160 448.530 ;
        RECT 2112.420 448.470 2112.680 448.790 ;
        RECT 2111.560 448.390 2112.160 448.470 ;
        RECT 2112.020 434.850 2112.160 448.390 ;
        RECT 2111.960 434.530 2112.220 434.850 ;
        RECT 2112.420 386.250 2112.680 386.570 ;
        RECT 2112.480 338.290 2112.620 386.250 ;
        RECT 2111.960 337.970 2112.220 338.290 ;
        RECT 2112.420 337.970 2112.680 338.290 ;
        RECT 2112.020 303.690 2112.160 337.970 ;
        RECT 2112.020 303.550 2112.620 303.690 ;
        RECT 2112.480 241.730 2112.620 303.550 ;
        RECT 2111.960 241.410 2112.220 241.730 ;
        RECT 2112.420 241.410 2112.680 241.730 ;
        RECT 2112.020 207.130 2112.160 241.410 ;
        RECT 2112.020 206.990 2112.620 207.130 ;
        RECT 2112.480 138.370 2112.620 206.990 ;
        RECT 2111.960 138.050 2112.220 138.370 ;
        RECT 2112.420 138.050 2112.680 138.370 ;
        RECT 2112.020 112.870 2112.160 138.050 ;
        RECT 2110.580 112.550 2110.840 112.870 ;
        RECT 2111.960 112.550 2112.220 112.870 ;
        RECT 2110.640 48.610 2110.780 112.550 ;
        RECT 2110.580 48.290 2110.840 48.610 ;
        RECT 2111.960 48.290 2112.220 48.610 ;
        RECT 2112.020 25.490 2112.160 48.290 ;
        RECT 1881.960 25.170 1882.220 25.490 ;
        RECT 2111.960 25.170 2112.220 25.490 ;
        RECT 1882.020 2.400 1882.160 25.170 ;
        RECT 1881.810 -4.800 1882.370 2.400 ;
      LAYER via2 ;
        RECT 2111.950 917.520 2112.230 917.800 ;
        RECT 2113.330 917.520 2113.610 917.800 ;
      LAYER met3 ;
        RECT 2111.925 917.810 2112.255 917.825 ;
        RECT 2113.305 917.810 2113.635 917.825 ;
        RECT 2111.925 917.510 2113.635 917.810 ;
        RECT 2111.925 917.495 2112.255 917.510 ;
        RECT 2113.305 917.495 2113.635 917.510 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1899.870 31.180 1900.190 31.240 ;
        RECT 2125.730 31.180 2126.050 31.240 ;
        RECT 1899.870 31.040 2126.050 31.180 ;
        RECT 1899.870 30.980 1900.190 31.040 ;
        RECT 2125.730 30.980 2126.050 31.040 ;
      LAYER via ;
        RECT 1899.900 30.980 1900.160 31.240 ;
        RECT 2125.760 30.980 2126.020 31.240 ;
      LAYER met2 ;
        RECT 2126.140 1700.410 2126.420 1704.000 ;
        RECT 2125.820 1700.270 2126.420 1700.410 ;
        RECT 2125.820 31.270 2125.960 1700.270 ;
        RECT 2126.140 1700.000 2126.420 1700.270 ;
        RECT 1899.900 30.950 1900.160 31.270 ;
        RECT 2125.760 30.950 2126.020 31.270 ;
        RECT 1899.960 2.400 1900.100 30.950 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1917.810 25.740 1918.130 25.800 ;
        RECT 2133.550 25.740 2133.870 25.800 ;
        RECT 1917.810 25.600 2133.870 25.740 ;
        RECT 1917.810 25.540 1918.130 25.600 ;
        RECT 2133.550 25.540 2133.870 25.600 ;
      LAYER via ;
        RECT 1917.840 25.540 1918.100 25.800 ;
        RECT 2133.580 25.540 2133.840 25.800 ;
      LAYER met2 ;
        RECT 2135.340 1700.410 2135.620 1704.000 ;
        RECT 2133.640 1700.270 2135.620 1700.410 ;
        RECT 2133.640 25.830 2133.780 1700.270 ;
        RECT 2135.340 1700.000 2135.620 1700.270 ;
        RECT 1917.840 25.510 1918.100 25.830 ;
        RECT 2133.580 25.510 2133.840 25.830 ;
        RECT 1917.900 2.400 1918.040 25.510 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2139.605 1594.005 2139.775 1642.115 ;
        RECT 2140.065 1497.445 2140.235 1545.555 ;
        RECT 2139.605 496.485 2139.775 531.335 ;
        RECT 2139.605 338.045 2139.775 381.735 ;
        RECT 2139.145 96.985 2139.315 144.755 ;
        RECT 2139.145 48.365 2139.315 96.475 ;
      LAYER mcon ;
        RECT 2139.605 1641.945 2139.775 1642.115 ;
        RECT 2140.065 1545.385 2140.235 1545.555 ;
        RECT 2139.605 531.165 2139.775 531.335 ;
        RECT 2139.605 381.565 2139.775 381.735 ;
        RECT 2139.145 144.585 2139.315 144.755 ;
        RECT 2139.145 96.305 2139.315 96.475 ;
      LAYER met1 ;
        RECT 2139.990 1671.680 2140.310 1671.740 ;
        RECT 2142.290 1671.680 2142.610 1671.740 ;
        RECT 2139.990 1671.540 2142.610 1671.680 ;
        RECT 2139.990 1671.480 2140.310 1671.540 ;
        RECT 2142.290 1671.480 2142.610 1671.540 ;
        RECT 2139.545 1642.100 2139.835 1642.145 ;
        RECT 2139.990 1642.100 2140.310 1642.160 ;
        RECT 2139.545 1641.960 2140.310 1642.100 ;
        RECT 2139.545 1641.915 2139.835 1641.960 ;
        RECT 2139.990 1641.900 2140.310 1641.960 ;
        RECT 2139.530 1594.160 2139.850 1594.220 ;
        RECT 2139.335 1594.020 2139.850 1594.160 ;
        RECT 2139.530 1593.960 2139.850 1594.020 ;
        RECT 2139.070 1559.140 2139.390 1559.200 ;
        RECT 2139.990 1559.140 2140.310 1559.200 ;
        RECT 2139.070 1559.000 2140.310 1559.140 ;
        RECT 2139.070 1558.940 2139.390 1559.000 ;
        RECT 2139.990 1558.940 2140.310 1559.000 ;
        RECT 2139.990 1545.540 2140.310 1545.600 ;
        RECT 2139.795 1545.400 2140.310 1545.540 ;
        RECT 2139.990 1545.340 2140.310 1545.400 ;
        RECT 2139.990 1497.600 2140.310 1497.660 ;
        RECT 2139.795 1497.460 2140.310 1497.600 ;
        RECT 2139.990 1497.400 2140.310 1497.460 ;
        RECT 2139.070 1414.640 2139.390 1414.700 ;
        RECT 2139.990 1414.640 2140.310 1414.700 ;
        RECT 2139.070 1414.500 2140.310 1414.640 ;
        RECT 2139.070 1414.440 2139.390 1414.500 ;
        RECT 2139.990 1414.440 2140.310 1414.500 ;
        RECT 2139.070 1318.080 2139.390 1318.140 ;
        RECT 2139.990 1318.080 2140.310 1318.140 ;
        RECT 2139.070 1317.940 2140.310 1318.080 ;
        RECT 2139.070 1317.880 2139.390 1317.940 ;
        RECT 2139.990 1317.880 2140.310 1317.940 ;
        RECT 2139.070 1221.520 2139.390 1221.580 ;
        RECT 2139.990 1221.520 2140.310 1221.580 ;
        RECT 2139.070 1221.380 2140.310 1221.520 ;
        RECT 2139.070 1221.320 2139.390 1221.380 ;
        RECT 2139.990 1221.320 2140.310 1221.380 ;
        RECT 2139.070 1124.960 2139.390 1125.020 ;
        RECT 2139.990 1124.960 2140.310 1125.020 ;
        RECT 2139.070 1124.820 2140.310 1124.960 ;
        RECT 2139.070 1124.760 2139.390 1124.820 ;
        RECT 2139.990 1124.760 2140.310 1124.820 ;
        RECT 2139.070 1028.400 2139.390 1028.460 ;
        RECT 2139.990 1028.400 2140.310 1028.460 ;
        RECT 2139.070 1028.260 2140.310 1028.400 ;
        RECT 2139.070 1028.200 2139.390 1028.260 ;
        RECT 2139.990 1028.200 2140.310 1028.260 ;
        RECT 2139.070 931.840 2139.390 931.900 ;
        RECT 2139.990 931.840 2140.310 931.900 ;
        RECT 2139.070 931.700 2140.310 931.840 ;
        RECT 2139.070 931.640 2139.390 931.700 ;
        RECT 2139.990 931.640 2140.310 931.700 ;
        RECT 2138.610 724.440 2138.930 724.500 ;
        RECT 2139.990 724.440 2140.310 724.500 ;
        RECT 2138.610 724.300 2140.310 724.440 ;
        RECT 2138.610 724.240 2138.930 724.300 ;
        RECT 2139.990 724.240 2140.310 724.300 ;
        RECT 2139.530 531.320 2139.850 531.380 ;
        RECT 2139.335 531.180 2139.850 531.320 ;
        RECT 2139.530 531.120 2139.850 531.180 ;
        RECT 2139.530 496.640 2139.850 496.700 ;
        RECT 2139.335 496.500 2139.850 496.640 ;
        RECT 2139.530 496.440 2139.850 496.500 ;
        RECT 2139.070 448.700 2139.390 448.760 ;
        RECT 2139.990 448.700 2140.310 448.760 ;
        RECT 2139.070 448.560 2140.310 448.700 ;
        RECT 2139.070 448.500 2139.390 448.560 ;
        RECT 2139.990 448.500 2140.310 448.560 ;
        RECT 2139.530 381.720 2139.850 381.780 ;
        RECT 2139.335 381.580 2139.850 381.720 ;
        RECT 2139.530 381.520 2139.850 381.580 ;
        RECT 2139.545 338.200 2139.835 338.245 ;
        RECT 2139.990 338.200 2140.310 338.260 ;
        RECT 2139.545 338.060 2140.310 338.200 ;
        RECT 2139.545 338.015 2139.835 338.060 ;
        RECT 2139.990 338.000 2140.310 338.060 ;
        RECT 2139.085 144.740 2139.375 144.785 ;
        RECT 2139.530 144.740 2139.850 144.800 ;
        RECT 2139.085 144.600 2139.850 144.740 ;
        RECT 2139.085 144.555 2139.375 144.600 ;
        RECT 2139.530 144.540 2139.850 144.600 ;
        RECT 2139.070 97.140 2139.390 97.200 ;
        RECT 2138.875 97.000 2139.390 97.140 ;
        RECT 2139.070 96.940 2139.390 97.000 ;
        RECT 2139.070 96.460 2139.390 96.520 ;
        RECT 2138.875 96.320 2139.390 96.460 ;
        RECT 2139.070 96.260 2139.390 96.320 ;
        RECT 2139.085 48.520 2139.375 48.565 ;
        RECT 2139.530 48.520 2139.850 48.580 ;
        RECT 2139.085 48.380 2139.850 48.520 ;
        RECT 2139.085 48.335 2139.375 48.380 ;
        RECT 2139.530 48.320 2139.850 48.380 ;
        RECT 1935.290 26.080 1935.610 26.140 ;
        RECT 2139.530 26.080 2139.850 26.140 ;
        RECT 1935.290 25.940 2139.850 26.080 ;
        RECT 1935.290 25.880 1935.610 25.940 ;
        RECT 2139.530 25.880 2139.850 25.940 ;
      LAYER via ;
        RECT 2140.020 1671.480 2140.280 1671.740 ;
        RECT 2142.320 1671.480 2142.580 1671.740 ;
        RECT 2140.020 1641.900 2140.280 1642.160 ;
        RECT 2139.560 1593.960 2139.820 1594.220 ;
        RECT 2139.100 1558.940 2139.360 1559.200 ;
        RECT 2140.020 1558.940 2140.280 1559.200 ;
        RECT 2140.020 1545.340 2140.280 1545.600 ;
        RECT 2140.020 1497.400 2140.280 1497.660 ;
        RECT 2139.100 1414.440 2139.360 1414.700 ;
        RECT 2140.020 1414.440 2140.280 1414.700 ;
        RECT 2139.100 1317.880 2139.360 1318.140 ;
        RECT 2140.020 1317.880 2140.280 1318.140 ;
        RECT 2139.100 1221.320 2139.360 1221.580 ;
        RECT 2140.020 1221.320 2140.280 1221.580 ;
        RECT 2139.100 1124.760 2139.360 1125.020 ;
        RECT 2140.020 1124.760 2140.280 1125.020 ;
        RECT 2139.100 1028.200 2139.360 1028.460 ;
        RECT 2140.020 1028.200 2140.280 1028.460 ;
        RECT 2139.100 931.640 2139.360 931.900 ;
        RECT 2140.020 931.640 2140.280 931.900 ;
        RECT 2138.640 724.240 2138.900 724.500 ;
        RECT 2140.020 724.240 2140.280 724.500 ;
        RECT 2139.560 531.120 2139.820 531.380 ;
        RECT 2139.560 496.440 2139.820 496.700 ;
        RECT 2139.100 448.500 2139.360 448.760 ;
        RECT 2140.020 448.500 2140.280 448.760 ;
        RECT 2139.560 381.520 2139.820 381.780 ;
        RECT 2140.020 338.000 2140.280 338.260 ;
        RECT 2139.560 144.540 2139.820 144.800 ;
        RECT 2139.100 96.940 2139.360 97.200 ;
        RECT 2139.100 96.260 2139.360 96.520 ;
        RECT 2139.560 48.320 2139.820 48.580 ;
        RECT 1935.320 25.880 1935.580 26.140 ;
        RECT 2139.560 25.880 2139.820 26.140 ;
      LAYER met2 ;
        RECT 2144.540 1700.410 2144.820 1704.000 ;
        RECT 2142.380 1700.270 2144.820 1700.410 ;
        RECT 2142.380 1671.770 2142.520 1700.270 ;
        RECT 2144.540 1700.000 2144.820 1700.270 ;
        RECT 2140.020 1671.450 2140.280 1671.770 ;
        RECT 2142.320 1671.450 2142.580 1671.770 ;
        RECT 2140.080 1642.190 2140.220 1671.450 ;
        RECT 2140.020 1641.870 2140.280 1642.190 ;
        RECT 2139.560 1593.930 2139.820 1594.250 ;
        RECT 2139.620 1559.650 2139.760 1593.930 ;
        RECT 2139.160 1559.510 2139.760 1559.650 ;
        RECT 2139.160 1559.230 2139.300 1559.510 ;
        RECT 2139.100 1558.910 2139.360 1559.230 ;
        RECT 2140.020 1558.910 2140.280 1559.230 ;
        RECT 2140.080 1545.630 2140.220 1558.910 ;
        RECT 2140.020 1545.310 2140.280 1545.630 ;
        RECT 2140.020 1497.370 2140.280 1497.690 ;
        RECT 2140.080 1414.730 2140.220 1497.370 ;
        RECT 2139.100 1414.410 2139.360 1414.730 ;
        RECT 2140.020 1414.410 2140.280 1414.730 ;
        RECT 2139.160 1414.130 2139.300 1414.410 ;
        RECT 2139.160 1413.990 2139.760 1414.130 ;
        RECT 2139.620 1366.530 2139.760 1413.990 ;
        RECT 2139.620 1366.390 2140.220 1366.530 ;
        RECT 2140.080 1318.170 2140.220 1366.390 ;
        RECT 2139.100 1317.850 2139.360 1318.170 ;
        RECT 2140.020 1317.850 2140.280 1318.170 ;
        RECT 2139.160 1317.570 2139.300 1317.850 ;
        RECT 2139.160 1317.430 2139.760 1317.570 ;
        RECT 2139.620 1269.970 2139.760 1317.430 ;
        RECT 2139.620 1269.830 2140.220 1269.970 ;
        RECT 2140.080 1221.610 2140.220 1269.830 ;
        RECT 2139.100 1221.290 2139.360 1221.610 ;
        RECT 2140.020 1221.290 2140.280 1221.610 ;
        RECT 2139.160 1221.010 2139.300 1221.290 ;
        RECT 2139.160 1220.870 2139.760 1221.010 ;
        RECT 2139.620 1173.410 2139.760 1220.870 ;
        RECT 2139.620 1173.270 2140.220 1173.410 ;
        RECT 2140.080 1125.050 2140.220 1173.270 ;
        RECT 2139.100 1124.730 2139.360 1125.050 ;
        RECT 2140.020 1124.730 2140.280 1125.050 ;
        RECT 2139.160 1124.450 2139.300 1124.730 ;
        RECT 2139.160 1124.310 2139.760 1124.450 ;
        RECT 2139.620 1076.850 2139.760 1124.310 ;
        RECT 2139.620 1076.710 2140.220 1076.850 ;
        RECT 2140.080 1028.490 2140.220 1076.710 ;
        RECT 2139.100 1028.170 2139.360 1028.490 ;
        RECT 2140.020 1028.170 2140.280 1028.490 ;
        RECT 2139.160 1027.890 2139.300 1028.170 ;
        RECT 2139.160 1027.750 2140.220 1027.890 ;
        RECT 2140.080 931.930 2140.220 1027.750 ;
        RECT 2139.100 931.610 2139.360 931.930 ;
        RECT 2140.020 931.610 2140.280 931.930 ;
        RECT 2139.160 931.330 2139.300 931.610 ;
        RECT 2139.160 931.190 2139.760 931.330 ;
        RECT 2139.620 835.450 2139.760 931.190 ;
        RECT 2139.160 835.310 2139.760 835.450 ;
        RECT 2139.160 834.770 2139.300 835.310 ;
        RECT 2139.160 834.630 2139.760 834.770 ;
        RECT 2139.620 738.890 2139.760 834.630 ;
        RECT 2139.160 738.750 2139.760 738.890 ;
        RECT 2139.160 738.210 2139.300 738.750 ;
        RECT 2139.160 738.070 2140.220 738.210 ;
        RECT 2140.080 724.530 2140.220 738.070 ;
        RECT 2138.640 724.210 2138.900 724.530 ;
        RECT 2140.020 724.210 2140.280 724.530 ;
        RECT 2138.700 676.445 2138.840 724.210 ;
        RECT 2138.630 676.075 2138.910 676.445 ;
        RECT 2139.550 676.075 2139.830 676.445 ;
        RECT 2139.620 642.330 2139.760 676.075 ;
        RECT 2139.160 642.190 2139.760 642.330 ;
        RECT 2139.160 641.650 2139.300 642.190 ;
        RECT 2139.160 641.510 2139.760 641.650 ;
        RECT 2139.620 545.770 2139.760 641.510 ;
        RECT 2139.160 545.630 2139.760 545.770 ;
        RECT 2139.160 545.090 2139.300 545.630 ;
        RECT 2139.160 544.950 2139.760 545.090 ;
        RECT 2139.620 531.410 2139.760 544.950 ;
        RECT 2139.560 531.090 2139.820 531.410 ;
        RECT 2139.560 496.410 2139.820 496.730 ;
        RECT 2139.620 483.210 2139.760 496.410 ;
        RECT 2139.620 483.070 2140.220 483.210 ;
        RECT 2140.080 448.790 2140.220 483.070 ;
        RECT 2139.100 448.530 2139.360 448.790 ;
        RECT 2139.100 448.470 2139.760 448.530 ;
        RECT 2140.020 448.470 2140.280 448.790 ;
        RECT 2139.160 448.390 2139.760 448.470 ;
        RECT 2139.620 381.810 2139.760 448.390 ;
        RECT 2139.560 381.490 2139.820 381.810 ;
        RECT 2140.020 337.970 2140.280 338.290 ;
        RECT 2140.080 255.410 2140.220 337.970 ;
        RECT 2139.160 255.270 2140.220 255.410 ;
        RECT 2139.160 254.730 2139.300 255.270 ;
        RECT 2139.160 254.590 2139.760 254.730 ;
        RECT 2139.620 159.530 2139.760 254.590 ;
        RECT 2139.620 159.390 2140.220 159.530 ;
        RECT 2140.080 145.250 2140.220 159.390 ;
        RECT 2139.620 145.110 2140.220 145.250 ;
        RECT 2139.620 144.830 2139.760 145.110 ;
        RECT 2139.560 144.510 2139.820 144.830 ;
        RECT 2139.100 96.910 2139.360 97.230 ;
        RECT 2139.160 96.550 2139.300 96.910 ;
        RECT 2139.100 96.230 2139.360 96.550 ;
        RECT 2139.560 48.290 2139.820 48.610 ;
        RECT 2139.620 26.170 2139.760 48.290 ;
        RECT 1935.320 25.850 1935.580 26.170 ;
        RECT 2139.560 25.850 2139.820 26.170 ;
        RECT 1935.380 2.400 1935.520 25.850 ;
        RECT 1935.170 -4.800 1935.730 2.400 ;
      LAYER via2 ;
        RECT 2138.630 676.120 2138.910 676.400 ;
        RECT 2139.550 676.120 2139.830 676.400 ;
      LAYER met3 ;
        RECT 2138.605 676.410 2138.935 676.425 ;
        RECT 2139.525 676.410 2139.855 676.425 ;
        RECT 2138.605 676.110 2139.855 676.410 ;
        RECT 2138.605 676.095 2138.935 676.110 ;
        RECT 2139.525 676.095 2139.855 676.110 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1953.230 26.420 1953.550 26.480 ;
        RECT 2153.330 26.420 2153.650 26.480 ;
        RECT 1953.230 26.280 2153.650 26.420 ;
        RECT 1953.230 26.220 1953.550 26.280 ;
        RECT 2153.330 26.220 2153.650 26.280 ;
      LAYER via ;
        RECT 1953.260 26.220 1953.520 26.480 ;
        RECT 2153.360 26.220 2153.620 26.480 ;
      LAYER met2 ;
        RECT 2153.740 1700.410 2154.020 1704.000 ;
        RECT 2153.420 1700.270 2154.020 1700.410 ;
        RECT 2153.420 26.510 2153.560 1700.270 ;
        RECT 2153.740 1700.000 2154.020 1700.270 ;
        RECT 1953.260 26.190 1953.520 26.510 ;
        RECT 2153.360 26.190 2153.620 26.510 ;
        RECT 1953.320 2.400 1953.460 26.190 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1971.170 26.760 1971.490 26.820 ;
        RECT 2160.690 26.760 2161.010 26.820 ;
        RECT 1971.170 26.620 2161.010 26.760 ;
        RECT 1971.170 26.560 1971.490 26.620 ;
        RECT 2160.690 26.560 2161.010 26.620 ;
      LAYER via ;
        RECT 1971.200 26.560 1971.460 26.820 ;
        RECT 2160.720 26.560 2160.980 26.820 ;
      LAYER met2 ;
        RECT 2162.940 1700.410 2163.220 1704.000 ;
        RECT 2160.780 1700.270 2163.220 1700.410 ;
        RECT 2160.780 26.850 2160.920 1700.270 ;
        RECT 2162.940 1700.000 2163.220 1700.270 ;
        RECT 1971.200 26.530 1971.460 26.850 ;
        RECT 2160.720 26.530 2160.980 26.850 ;
        RECT 1971.260 2.400 1971.400 26.530 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2168.585 1594.005 2168.755 1642.115 ;
        RECT 2167.205 1497.445 2167.375 1545.555 ;
        RECT 2168.125 1352.605 2168.295 1400.715 ;
        RECT 2168.125 1256.045 2168.295 1304.155 ;
        RECT 2168.585 966.025 2168.755 980.475 ;
        RECT 2168.125 579.785 2168.295 627.895 ;
        RECT 2168.125 496.485 2168.295 531.335 ;
        RECT 2168.125 386.325 2168.295 401.115 ;
        RECT 2168.125 241.485 2168.295 289.595 ;
      LAYER mcon ;
        RECT 2168.585 1641.945 2168.755 1642.115 ;
        RECT 2167.205 1545.385 2167.375 1545.555 ;
        RECT 2168.125 1400.545 2168.295 1400.715 ;
        RECT 2168.125 1303.985 2168.295 1304.155 ;
        RECT 2168.585 980.305 2168.755 980.475 ;
        RECT 2168.125 627.725 2168.295 627.895 ;
        RECT 2168.125 531.165 2168.295 531.335 ;
        RECT 2168.125 400.945 2168.295 401.115 ;
        RECT 2168.125 289.425 2168.295 289.595 ;
      LAYER met1 ;
        RECT 2168.510 1642.100 2168.830 1642.160 ;
        RECT 2168.315 1641.960 2168.830 1642.100 ;
        RECT 2168.510 1641.900 2168.830 1641.960 ;
        RECT 2168.525 1594.160 2168.815 1594.205 ;
        RECT 2168.970 1594.160 2169.290 1594.220 ;
        RECT 2168.525 1594.020 2169.290 1594.160 ;
        RECT 2168.525 1593.975 2168.815 1594.020 ;
        RECT 2168.970 1593.960 2169.290 1594.020 ;
        RECT 2167.130 1559.480 2167.450 1559.540 ;
        RECT 2168.970 1559.480 2169.290 1559.540 ;
        RECT 2167.130 1559.340 2169.290 1559.480 ;
        RECT 2167.130 1559.280 2167.450 1559.340 ;
        RECT 2168.970 1559.280 2169.290 1559.340 ;
        RECT 2167.130 1545.540 2167.450 1545.600 ;
        RECT 2166.935 1545.400 2167.450 1545.540 ;
        RECT 2167.130 1545.340 2167.450 1545.400 ;
        RECT 2167.145 1497.600 2167.435 1497.645 ;
        RECT 2168.510 1497.600 2168.830 1497.660 ;
        RECT 2167.145 1497.460 2168.830 1497.600 ;
        RECT 2167.145 1497.415 2167.435 1497.460 ;
        RECT 2168.510 1497.400 2168.830 1497.460 ;
        RECT 2168.050 1400.700 2168.370 1400.760 ;
        RECT 2167.855 1400.560 2168.370 1400.700 ;
        RECT 2168.050 1400.500 2168.370 1400.560 ;
        RECT 2168.065 1352.760 2168.355 1352.805 ;
        RECT 2168.510 1352.760 2168.830 1352.820 ;
        RECT 2168.065 1352.620 2168.830 1352.760 ;
        RECT 2168.065 1352.575 2168.355 1352.620 ;
        RECT 2168.510 1352.560 2168.830 1352.620 ;
        RECT 2168.050 1304.140 2168.370 1304.200 ;
        RECT 2167.855 1304.000 2168.370 1304.140 ;
        RECT 2168.050 1303.940 2168.370 1304.000 ;
        RECT 2168.065 1256.200 2168.355 1256.245 ;
        RECT 2168.510 1256.200 2168.830 1256.260 ;
        RECT 2168.065 1256.060 2168.830 1256.200 ;
        RECT 2168.065 1256.015 2168.355 1256.060 ;
        RECT 2168.510 1256.000 2168.830 1256.060 ;
        RECT 2167.130 1159.300 2167.450 1159.360 ;
        RECT 2168.510 1159.300 2168.830 1159.360 ;
        RECT 2167.130 1159.160 2168.830 1159.300 ;
        RECT 2167.130 1159.100 2167.450 1159.160 ;
        RECT 2168.510 1159.100 2168.830 1159.160 ;
        RECT 2167.130 1062.740 2167.450 1062.800 ;
        RECT 2168.510 1062.740 2168.830 1062.800 ;
        RECT 2167.130 1062.600 2168.830 1062.740 ;
        RECT 2167.130 1062.540 2167.450 1062.600 ;
        RECT 2168.510 1062.540 2168.830 1062.600 ;
        RECT 2168.510 980.460 2168.830 980.520 ;
        RECT 2168.315 980.320 2168.830 980.460 ;
        RECT 2168.510 980.260 2168.830 980.320 ;
        RECT 2168.510 966.180 2168.830 966.240 ;
        RECT 2168.315 966.040 2168.830 966.180 ;
        RECT 2168.510 965.980 2168.830 966.040 ;
        RECT 2168.050 869.620 2168.370 869.680 ;
        RECT 2168.510 869.620 2168.830 869.680 ;
        RECT 2168.050 869.480 2168.830 869.620 ;
        RECT 2168.050 869.420 2168.370 869.480 ;
        RECT 2168.510 869.420 2168.830 869.480 ;
        RECT 2168.050 738.520 2168.370 738.780 ;
        RECT 2168.140 738.100 2168.280 738.520 ;
        RECT 2168.050 737.840 2168.370 738.100 ;
        RECT 2168.050 627.880 2168.370 627.940 ;
        RECT 2167.855 627.740 2168.370 627.880 ;
        RECT 2168.050 627.680 2168.370 627.740 ;
        RECT 2168.050 579.940 2168.370 580.000 ;
        RECT 2167.855 579.800 2168.370 579.940 ;
        RECT 2168.050 579.740 2168.370 579.800 ;
        RECT 2168.050 531.320 2168.370 531.380 ;
        RECT 2167.855 531.180 2168.370 531.320 ;
        RECT 2168.050 531.120 2168.370 531.180 ;
        RECT 2168.050 496.640 2168.370 496.700 ;
        RECT 2167.855 496.500 2168.370 496.640 ;
        RECT 2168.050 496.440 2168.370 496.500 ;
        RECT 2168.065 401.100 2168.355 401.145 ;
        RECT 2168.510 401.100 2168.830 401.160 ;
        RECT 2168.065 400.960 2168.830 401.100 ;
        RECT 2168.065 400.915 2168.355 400.960 ;
        RECT 2168.510 400.900 2168.830 400.960 ;
        RECT 2168.050 386.480 2168.370 386.540 ;
        RECT 2167.855 386.340 2168.370 386.480 ;
        RECT 2168.050 386.280 2168.370 386.340 ;
        RECT 2167.590 303.520 2167.910 303.580 ;
        RECT 2168.510 303.520 2168.830 303.580 ;
        RECT 2167.590 303.380 2168.830 303.520 ;
        RECT 2167.590 303.320 2167.910 303.380 ;
        RECT 2168.510 303.320 2168.830 303.380 ;
        RECT 2168.065 289.580 2168.355 289.625 ;
        RECT 2168.510 289.580 2168.830 289.640 ;
        RECT 2168.065 289.440 2168.830 289.580 ;
        RECT 2168.065 289.395 2168.355 289.440 ;
        RECT 2168.510 289.380 2168.830 289.440 ;
        RECT 2168.050 241.640 2168.370 241.700 ;
        RECT 2167.855 241.500 2168.370 241.640 ;
        RECT 2168.050 241.440 2168.370 241.500 ;
        RECT 1989.110 27.100 1989.430 27.160 ;
        RECT 2168.050 27.100 2168.370 27.160 ;
        RECT 1989.110 26.960 2168.370 27.100 ;
        RECT 1989.110 26.900 1989.430 26.960 ;
        RECT 2168.050 26.900 2168.370 26.960 ;
      LAYER via ;
        RECT 2168.540 1641.900 2168.800 1642.160 ;
        RECT 2169.000 1593.960 2169.260 1594.220 ;
        RECT 2167.160 1559.280 2167.420 1559.540 ;
        RECT 2169.000 1559.280 2169.260 1559.540 ;
        RECT 2167.160 1545.340 2167.420 1545.600 ;
        RECT 2168.540 1497.400 2168.800 1497.660 ;
        RECT 2168.080 1400.500 2168.340 1400.760 ;
        RECT 2168.540 1352.560 2168.800 1352.820 ;
        RECT 2168.080 1303.940 2168.340 1304.200 ;
        RECT 2168.540 1256.000 2168.800 1256.260 ;
        RECT 2167.160 1159.100 2167.420 1159.360 ;
        RECT 2168.540 1159.100 2168.800 1159.360 ;
        RECT 2167.160 1062.540 2167.420 1062.800 ;
        RECT 2168.540 1062.540 2168.800 1062.800 ;
        RECT 2168.540 980.260 2168.800 980.520 ;
        RECT 2168.540 965.980 2168.800 966.240 ;
        RECT 2168.080 869.420 2168.340 869.680 ;
        RECT 2168.540 869.420 2168.800 869.680 ;
        RECT 2168.080 738.520 2168.340 738.780 ;
        RECT 2168.080 737.840 2168.340 738.100 ;
        RECT 2168.080 627.680 2168.340 627.940 ;
        RECT 2168.080 579.740 2168.340 580.000 ;
        RECT 2168.080 531.120 2168.340 531.380 ;
        RECT 2168.080 496.440 2168.340 496.700 ;
        RECT 2168.540 400.900 2168.800 401.160 ;
        RECT 2168.080 386.280 2168.340 386.540 ;
        RECT 2167.620 303.320 2167.880 303.580 ;
        RECT 2168.540 303.320 2168.800 303.580 ;
        RECT 2168.540 289.380 2168.800 289.640 ;
        RECT 2168.080 241.440 2168.340 241.700 ;
        RECT 1989.140 26.900 1989.400 27.160 ;
        RECT 2168.080 26.900 2168.340 27.160 ;
      LAYER met2 ;
        RECT 2172.140 1700.410 2172.420 1704.000 ;
        RECT 2170.900 1700.270 2172.420 1700.410 ;
        RECT 2170.900 1643.405 2171.040 1700.270 ;
        RECT 2172.140 1700.000 2172.420 1700.270 ;
        RECT 2170.830 1643.035 2171.110 1643.405 ;
        RECT 2168.530 1642.355 2168.810 1642.725 ;
        RECT 2168.600 1642.190 2168.740 1642.355 ;
        RECT 2168.540 1641.870 2168.800 1642.190 ;
        RECT 2169.000 1593.930 2169.260 1594.250 ;
        RECT 2169.060 1559.570 2169.200 1593.930 ;
        RECT 2167.160 1559.250 2167.420 1559.570 ;
        RECT 2169.000 1559.250 2169.260 1559.570 ;
        RECT 2167.220 1545.630 2167.360 1559.250 ;
        RECT 2167.160 1545.310 2167.420 1545.630 ;
        RECT 2168.540 1497.370 2168.800 1497.690 ;
        RECT 2168.600 1425.010 2168.740 1497.370 ;
        RECT 2168.140 1424.870 2168.740 1425.010 ;
        RECT 2168.140 1400.790 2168.280 1424.870 ;
        RECT 2168.080 1400.470 2168.340 1400.790 ;
        RECT 2168.540 1352.530 2168.800 1352.850 ;
        RECT 2168.600 1317.570 2168.740 1352.530 ;
        RECT 2168.140 1317.430 2168.740 1317.570 ;
        RECT 2168.140 1304.230 2168.280 1317.430 ;
        RECT 2168.080 1303.910 2168.340 1304.230 ;
        RECT 2168.540 1255.970 2168.800 1256.290 ;
        RECT 2168.600 1221.010 2168.740 1255.970 ;
        RECT 2168.140 1220.870 2168.740 1221.010 ;
        RECT 2168.140 1207.525 2168.280 1220.870 ;
        RECT 2167.150 1207.155 2167.430 1207.525 ;
        RECT 2168.070 1207.155 2168.350 1207.525 ;
        RECT 2167.220 1159.390 2167.360 1207.155 ;
        RECT 2167.160 1159.070 2167.420 1159.390 ;
        RECT 2168.540 1159.070 2168.800 1159.390 ;
        RECT 2168.600 1124.450 2168.740 1159.070 ;
        RECT 2168.140 1124.310 2168.740 1124.450 ;
        RECT 2168.140 1110.965 2168.280 1124.310 ;
        RECT 2167.150 1110.595 2167.430 1110.965 ;
        RECT 2168.070 1110.595 2168.350 1110.965 ;
        RECT 2167.220 1062.830 2167.360 1110.595 ;
        RECT 2167.160 1062.510 2167.420 1062.830 ;
        RECT 2168.540 1062.510 2168.800 1062.830 ;
        RECT 2168.600 980.550 2168.740 1062.510 ;
        RECT 2168.540 980.230 2168.800 980.550 ;
        RECT 2168.540 965.950 2168.800 966.270 ;
        RECT 2168.600 869.710 2168.740 965.950 ;
        RECT 2168.080 869.390 2168.340 869.710 ;
        RECT 2168.540 869.390 2168.800 869.710 ;
        RECT 2168.140 787.170 2168.280 869.390 ;
        RECT 2167.680 787.030 2168.280 787.170 ;
        RECT 2167.680 786.490 2167.820 787.030 ;
        RECT 2167.680 786.350 2168.280 786.490 ;
        RECT 2168.140 738.810 2168.280 786.350 ;
        RECT 2168.080 738.490 2168.340 738.810 ;
        RECT 2168.080 737.810 2168.340 738.130 ;
        RECT 2168.140 627.970 2168.280 737.810 ;
        RECT 2168.080 627.650 2168.340 627.970 ;
        RECT 2168.080 579.710 2168.340 580.030 ;
        RECT 2168.140 531.410 2168.280 579.710 ;
        RECT 2168.080 531.090 2168.340 531.410 ;
        RECT 2168.080 496.410 2168.340 496.730 ;
        RECT 2168.140 483.210 2168.280 496.410 ;
        RECT 2168.140 483.070 2168.740 483.210 ;
        RECT 2168.600 401.190 2168.740 483.070 ;
        RECT 2168.540 400.870 2168.800 401.190 ;
        RECT 2168.080 386.250 2168.340 386.570 ;
        RECT 2168.140 303.690 2168.280 386.250 ;
        RECT 2167.680 303.610 2168.280 303.690 ;
        RECT 2167.620 303.550 2168.280 303.610 ;
        RECT 2167.620 303.290 2167.880 303.550 ;
        RECT 2168.540 303.290 2168.800 303.610 ;
        RECT 2168.600 289.670 2168.740 303.290 ;
        RECT 2168.540 289.350 2168.800 289.670 ;
        RECT 2168.080 241.410 2168.340 241.730 ;
        RECT 2168.140 207.130 2168.280 241.410 ;
        RECT 2167.680 206.990 2168.280 207.130 ;
        RECT 2167.680 206.450 2167.820 206.990 ;
        RECT 2167.680 206.310 2168.280 206.450 ;
        RECT 2168.140 110.570 2168.280 206.310 ;
        RECT 2167.680 110.430 2168.280 110.570 ;
        RECT 2167.680 109.890 2167.820 110.430 ;
        RECT 2167.680 109.750 2168.280 109.890 ;
        RECT 2168.140 27.190 2168.280 109.750 ;
        RECT 1989.140 26.870 1989.400 27.190 ;
        RECT 2168.080 26.870 2168.340 27.190 ;
        RECT 1989.200 2.400 1989.340 26.870 ;
        RECT 1988.990 -4.800 1989.550 2.400 ;
      LAYER via2 ;
        RECT 2170.830 1643.080 2171.110 1643.360 ;
        RECT 2168.530 1642.400 2168.810 1642.680 ;
        RECT 2167.150 1207.200 2167.430 1207.480 ;
        RECT 2168.070 1207.200 2168.350 1207.480 ;
        RECT 2167.150 1110.640 2167.430 1110.920 ;
        RECT 2168.070 1110.640 2168.350 1110.920 ;
      LAYER met3 ;
        RECT 2170.805 1643.370 2171.135 1643.385 ;
        RECT 2167.830 1643.070 2171.135 1643.370 ;
        RECT 2167.830 1642.690 2168.130 1643.070 ;
        RECT 2170.805 1643.055 2171.135 1643.070 ;
        RECT 2168.505 1642.690 2168.835 1642.705 ;
        RECT 2167.830 1642.390 2168.835 1642.690 ;
        RECT 2168.505 1642.375 2168.835 1642.390 ;
        RECT 2167.125 1207.490 2167.455 1207.505 ;
        RECT 2168.045 1207.490 2168.375 1207.505 ;
        RECT 2167.125 1207.190 2168.375 1207.490 ;
        RECT 2167.125 1207.175 2167.455 1207.190 ;
        RECT 2168.045 1207.175 2168.375 1207.190 ;
        RECT 2167.125 1110.930 2167.455 1110.945 ;
        RECT 2168.045 1110.930 2168.375 1110.945 ;
        RECT 2167.125 1110.630 2168.375 1110.930 ;
        RECT 2167.125 1110.615 2167.455 1110.630 ;
        RECT 2168.045 1110.615 2168.375 1110.630 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2006.590 27.440 2006.910 27.500 ;
        RECT 2180.930 27.440 2181.250 27.500 ;
        RECT 2006.590 27.300 2181.250 27.440 ;
        RECT 2006.590 27.240 2006.910 27.300 ;
        RECT 2180.930 27.240 2181.250 27.300 ;
      LAYER via ;
        RECT 2006.620 27.240 2006.880 27.500 ;
        RECT 2180.960 27.240 2181.220 27.500 ;
      LAYER met2 ;
        RECT 2181.340 1700.410 2181.620 1704.000 ;
        RECT 2181.020 1700.270 2181.620 1700.410 ;
        RECT 2181.020 27.530 2181.160 1700.270 ;
        RECT 2181.340 1700.000 2181.620 1700.270 ;
        RECT 2006.620 27.210 2006.880 27.530 ;
        RECT 2180.960 27.210 2181.220 27.530 ;
        RECT 2006.680 2.400 2006.820 27.210 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2024.530 23.700 2024.850 23.760 ;
        RECT 2188.750 23.700 2189.070 23.760 ;
        RECT 2024.530 23.560 2189.070 23.700 ;
        RECT 2024.530 23.500 2024.850 23.560 ;
        RECT 2188.750 23.500 2189.070 23.560 ;
      LAYER via ;
        RECT 2024.560 23.500 2024.820 23.760 ;
        RECT 2188.780 23.500 2189.040 23.760 ;
      LAYER met2 ;
        RECT 2190.540 1700.410 2190.820 1704.000 ;
        RECT 2188.840 1700.270 2190.820 1700.410 ;
        RECT 2188.840 23.790 2188.980 1700.270 ;
        RECT 2190.540 1700.000 2190.820 1700.270 ;
        RECT 2024.560 23.470 2024.820 23.790 ;
        RECT 2188.780 23.470 2189.040 23.790 ;
        RECT 2024.620 2.400 2024.760 23.470 ;
        RECT 2024.410 -4.800 2024.970 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2163.065 1688.865 2163.235 1689.715 ;
      LAYER mcon ;
        RECT 2163.065 1689.545 2163.235 1689.715 ;
      LAYER met1 ;
        RECT 2163.005 1689.700 2163.295 1689.745 ;
        RECT 2199.790 1689.700 2200.110 1689.760 ;
        RECT 2163.005 1689.560 2200.110 1689.700 ;
        RECT 2163.005 1689.515 2163.295 1689.560 ;
        RECT 2199.790 1689.500 2200.110 1689.560 ;
        RECT 2048.910 1689.020 2049.230 1689.080 ;
        RECT 2163.005 1689.020 2163.295 1689.065 ;
        RECT 2048.910 1688.880 2163.295 1689.020 ;
        RECT 2048.910 1688.820 2049.230 1688.880 ;
        RECT 2163.005 1688.835 2163.295 1688.880 ;
        RECT 2042.470 17.240 2042.790 17.300 ;
        RECT 2048.910 17.240 2049.230 17.300 ;
        RECT 2042.470 17.100 2049.230 17.240 ;
        RECT 2042.470 17.040 2042.790 17.100 ;
        RECT 2048.910 17.040 2049.230 17.100 ;
      LAYER via ;
        RECT 2199.820 1689.500 2200.080 1689.760 ;
        RECT 2048.940 1688.820 2049.200 1689.080 ;
        RECT 2042.500 17.040 2042.760 17.300 ;
        RECT 2048.940 17.040 2049.200 17.300 ;
      LAYER met2 ;
        RECT 2199.740 1700.000 2200.020 1704.000 ;
        RECT 2199.880 1689.790 2200.020 1700.000 ;
        RECT 2199.820 1689.470 2200.080 1689.790 ;
        RECT 2048.940 1688.790 2049.200 1689.110 ;
        RECT 2049.000 17.330 2049.140 1688.790 ;
        RECT 2042.500 17.010 2042.760 17.330 ;
        RECT 2048.940 17.010 2049.200 17.330 ;
        RECT 2042.560 2.400 2042.700 17.010 ;
        RECT 2042.350 -4.800 2042.910 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 758.610 66.880 758.930 66.940 ;
        RECT 1539.690 66.880 1540.010 66.940 ;
        RECT 758.610 66.740 1540.010 66.880 ;
        RECT 758.610 66.680 758.930 66.740 ;
        RECT 1539.690 66.680 1540.010 66.740 ;
      LAYER via ;
        RECT 758.640 66.680 758.900 66.940 ;
        RECT 1539.720 66.680 1539.980 66.940 ;
      LAYER met2 ;
        RECT 1538.720 1700.410 1539.000 1704.000 ;
        RECT 1538.720 1700.270 1539.920 1700.410 ;
        RECT 1538.720 1700.000 1539.000 1700.270 ;
        RECT 1539.780 66.970 1539.920 1700.270 ;
        RECT 758.640 66.650 758.900 66.970 ;
        RECT 1539.720 66.650 1539.980 66.970 ;
        RECT 758.700 17.410 758.840 66.650 ;
        RECT 757.780 17.270 758.840 17.410 ;
        RECT 757.780 2.400 757.920 17.270 ;
        RECT 757.570 -4.800 758.130 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2062.710 1688.680 2063.030 1688.740 ;
        RECT 2208.990 1688.680 2209.310 1688.740 ;
        RECT 2062.710 1688.540 2209.310 1688.680 ;
        RECT 2062.710 1688.480 2063.030 1688.540 ;
        RECT 2208.990 1688.480 2209.310 1688.540 ;
        RECT 2060.410 20.640 2060.730 20.700 ;
        RECT 2062.710 20.640 2063.030 20.700 ;
        RECT 2060.410 20.500 2063.030 20.640 ;
        RECT 2060.410 20.440 2060.730 20.500 ;
        RECT 2062.710 20.440 2063.030 20.500 ;
      LAYER via ;
        RECT 2062.740 1688.480 2063.000 1688.740 ;
        RECT 2209.020 1688.480 2209.280 1688.740 ;
        RECT 2060.440 20.440 2060.700 20.700 ;
        RECT 2062.740 20.440 2063.000 20.700 ;
      LAYER met2 ;
        RECT 2208.940 1700.000 2209.220 1704.000 ;
        RECT 2209.080 1688.770 2209.220 1700.000 ;
        RECT 2062.740 1688.450 2063.000 1688.770 ;
        RECT 2209.020 1688.450 2209.280 1688.770 ;
        RECT 2062.800 20.730 2062.940 1688.450 ;
        RECT 2060.440 20.410 2060.700 20.730 ;
        RECT 2062.740 20.410 2063.000 20.730 ;
        RECT 2060.500 2.400 2060.640 20.410 ;
        RECT 2060.290 -4.800 2060.850 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2083.410 1690.040 2083.730 1690.100 ;
        RECT 2218.190 1690.040 2218.510 1690.100 ;
        RECT 2083.410 1689.900 2218.510 1690.040 ;
        RECT 2083.410 1689.840 2083.730 1689.900 ;
        RECT 2218.190 1689.840 2218.510 1689.900 ;
        RECT 2078.350 20.640 2078.670 20.700 ;
        RECT 2083.410 20.640 2083.730 20.700 ;
        RECT 2078.350 20.500 2083.730 20.640 ;
        RECT 2078.350 20.440 2078.670 20.500 ;
        RECT 2083.410 20.440 2083.730 20.500 ;
      LAYER via ;
        RECT 2083.440 1689.840 2083.700 1690.100 ;
        RECT 2218.220 1689.840 2218.480 1690.100 ;
        RECT 2078.380 20.440 2078.640 20.700 ;
        RECT 2083.440 20.440 2083.700 20.700 ;
      LAYER met2 ;
        RECT 2218.140 1700.000 2218.420 1704.000 ;
        RECT 2218.280 1690.130 2218.420 1700.000 ;
        RECT 2083.440 1689.810 2083.700 1690.130 ;
        RECT 2218.220 1689.810 2218.480 1690.130 ;
        RECT 2083.500 20.730 2083.640 1689.810 ;
        RECT 2078.380 20.410 2078.640 20.730 ;
        RECT 2083.440 20.410 2083.700 20.730 ;
        RECT 2078.440 2.400 2078.580 20.410 ;
        RECT 2078.230 -4.800 2078.790 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2101.350 1690.380 2101.670 1690.440 ;
        RECT 2227.390 1690.380 2227.710 1690.440 ;
        RECT 2101.350 1690.240 2227.710 1690.380 ;
        RECT 2101.350 1690.180 2101.670 1690.240 ;
        RECT 2227.390 1690.180 2227.710 1690.240 ;
        RECT 2095.830 20.640 2096.150 20.700 ;
        RECT 2101.350 20.640 2101.670 20.700 ;
        RECT 2095.830 20.500 2101.670 20.640 ;
        RECT 2095.830 20.440 2096.150 20.500 ;
        RECT 2101.350 20.440 2101.670 20.500 ;
      LAYER via ;
        RECT 2101.380 1690.180 2101.640 1690.440 ;
        RECT 2227.420 1690.180 2227.680 1690.440 ;
        RECT 2095.860 20.440 2096.120 20.700 ;
        RECT 2101.380 20.440 2101.640 20.700 ;
      LAYER met2 ;
        RECT 2227.340 1700.000 2227.620 1704.000 ;
        RECT 2227.480 1690.470 2227.620 1700.000 ;
        RECT 2101.380 1690.150 2101.640 1690.470 ;
        RECT 2227.420 1690.150 2227.680 1690.470 ;
        RECT 2101.440 20.730 2101.580 1690.150 ;
        RECT 2095.860 20.410 2096.120 20.730 ;
        RECT 2101.380 20.410 2101.640 20.730 ;
        RECT 2095.920 2.400 2096.060 20.410 ;
        RECT 2095.710 -4.800 2096.270 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2163.065 1685.465 2163.235 1686.995 ;
      LAYER mcon ;
        RECT 2163.065 1686.825 2163.235 1686.995 ;
      LAYER met1 ;
        RECT 2163.005 1686.980 2163.295 1687.025 ;
        RECT 2236.590 1686.980 2236.910 1687.040 ;
        RECT 2163.005 1686.840 2236.910 1686.980 ;
        RECT 2163.005 1686.795 2163.295 1686.840 ;
        RECT 2236.590 1686.780 2236.910 1686.840 ;
        RECT 2117.910 1685.620 2118.230 1685.680 ;
        RECT 2163.005 1685.620 2163.295 1685.665 ;
        RECT 2117.910 1685.480 2163.295 1685.620 ;
        RECT 2117.910 1685.420 2118.230 1685.480 ;
        RECT 2163.005 1685.435 2163.295 1685.480 ;
        RECT 2113.770 20.640 2114.090 20.700 ;
        RECT 2117.910 20.640 2118.230 20.700 ;
        RECT 2113.770 20.500 2118.230 20.640 ;
        RECT 2113.770 20.440 2114.090 20.500 ;
        RECT 2117.910 20.440 2118.230 20.500 ;
      LAYER via ;
        RECT 2236.620 1686.780 2236.880 1687.040 ;
        RECT 2117.940 1685.420 2118.200 1685.680 ;
        RECT 2113.800 20.440 2114.060 20.700 ;
        RECT 2117.940 20.440 2118.200 20.700 ;
      LAYER met2 ;
        RECT 2236.540 1700.000 2236.820 1704.000 ;
        RECT 2236.680 1687.070 2236.820 1700.000 ;
        RECT 2236.620 1686.750 2236.880 1687.070 ;
        RECT 2117.940 1685.390 2118.200 1685.710 ;
        RECT 2118.000 20.730 2118.140 1685.390 ;
        RECT 2113.800 20.410 2114.060 20.730 ;
        RECT 2117.940 20.410 2118.200 20.730 ;
        RECT 2113.860 2.400 2114.000 20.410 ;
        RECT 2113.650 -4.800 2114.210 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2166.745 1685.805 2166.915 1686.655 ;
      LAYER mcon ;
        RECT 2166.745 1686.485 2166.915 1686.655 ;
      LAYER met1 ;
        RECT 2142.750 1686.640 2143.070 1686.700 ;
        RECT 2166.685 1686.640 2166.975 1686.685 ;
        RECT 2142.750 1686.500 2166.975 1686.640 ;
        RECT 2142.750 1686.440 2143.070 1686.500 ;
        RECT 2166.685 1686.455 2166.975 1686.500 ;
        RECT 2166.685 1685.960 2166.975 1686.005 ;
        RECT 2245.790 1685.960 2246.110 1686.020 ;
        RECT 2166.685 1685.820 2246.110 1685.960 ;
        RECT 2166.685 1685.775 2166.975 1685.820 ;
        RECT 2245.790 1685.760 2246.110 1685.820 ;
        RECT 2131.710 17.580 2132.030 17.640 ;
        RECT 2142.290 17.580 2142.610 17.640 ;
        RECT 2131.710 17.440 2142.610 17.580 ;
        RECT 2131.710 17.380 2132.030 17.440 ;
        RECT 2142.290 17.380 2142.610 17.440 ;
      LAYER via ;
        RECT 2142.780 1686.440 2143.040 1686.700 ;
        RECT 2245.820 1685.760 2246.080 1686.020 ;
        RECT 2131.740 17.380 2132.000 17.640 ;
        RECT 2142.320 17.380 2142.580 17.640 ;
      LAYER met2 ;
        RECT 2245.740 1700.000 2246.020 1704.000 ;
        RECT 2142.780 1686.410 2143.040 1686.730 ;
        RECT 2142.840 1671.170 2142.980 1686.410 ;
        RECT 2245.880 1686.050 2246.020 1700.000 ;
        RECT 2245.820 1685.730 2246.080 1686.050 ;
        RECT 2142.380 1671.030 2142.980 1671.170 ;
        RECT 2142.380 17.670 2142.520 1671.030 ;
        RECT 2131.740 17.350 2132.000 17.670 ;
        RECT 2142.320 17.350 2142.580 17.670 ;
        RECT 2131.800 2.400 2131.940 17.350 ;
        RECT 2131.590 -4.800 2132.150 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2179.165 1685.125 2179.335 1687.675 ;
        RECT 2162.605 1684.785 2164.155 1684.955 ;
        RECT 2162.605 1683.765 2162.775 1684.785 ;
      LAYER mcon ;
        RECT 2179.165 1687.505 2179.335 1687.675 ;
        RECT 2163.985 1684.785 2164.155 1684.955 ;
      LAYER met1 ;
        RECT 2179.105 1687.660 2179.395 1687.705 ;
        RECT 2254.990 1687.660 2255.310 1687.720 ;
        RECT 2179.105 1687.520 2255.310 1687.660 ;
        RECT 2179.105 1687.475 2179.395 1687.520 ;
        RECT 2254.990 1687.460 2255.310 1687.520 ;
        RECT 2179.105 1685.280 2179.395 1685.325 ;
        RECT 2164.460 1685.140 2179.395 1685.280 ;
        RECT 2163.925 1684.940 2164.215 1684.985 ;
        RECT 2164.460 1684.940 2164.600 1685.140 ;
        RECT 2179.105 1685.095 2179.395 1685.140 ;
        RECT 2163.925 1684.800 2164.600 1684.940 ;
        RECT 2163.925 1684.755 2164.215 1684.800 ;
        RECT 2152.410 1683.920 2152.730 1683.980 ;
        RECT 2162.545 1683.920 2162.835 1683.965 ;
        RECT 2152.410 1683.780 2162.835 1683.920 ;
        RECT 2152.410 1683.720 2152.730 1683.780 ;
        RECT 2162.545 1683.735 2162.835 1683.780 ;
        RECT 2149.650 20.640 2149.970 20.700 ;
        RECT 2152.410 20.640 2152.730 20.700 ;
        RECT 2149.650 20.500 2152.730 20.640 ;
        RECT 2149.650 20.440 2149.970 20.500 ;
        RECT 2152.410 20.440 2152.730 20.500 ;
      LAYER via ;
        RECT 2255.020 1687.460 2255.280 1687.720 ;
        RECT 2152.440 1683.720 2152.700 1683.980 ;
        RECT 2149.680 20.440 2149.940 20.700 ;
        RECT 2152.440 20.440 2152.700 20.700 ;
      LAYER met2 ;
        RECT 2254.940 1700.000 2255.220 1704.000 ;
        RECT 2255.080 1687.750 2255.220 1700.000 ;
        RECT 2255.020 1687.430 2255.280 1687.750 ;
        RECT 2152.440 1683.690 2152.700 1684.010 ;
        RECT 2152.500 20.730 2152.640 1683.690 ;
        RECT 2149.680 20.410 2149.940 20.730 ;
        RECT 2152.440 20.410 2152.700 20.730 ;
        RECT 2149.740 2.400 2149.880 20.410 ;
        RECT 2149.530 -4.800 2150.090 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2206.765 1684.785 2206.935 1688.015 ;
      LAYER mcon ;
        RECT 2206.765 1687.845 2206.935 1688.015 ;
      LAYER met1 ;
        RECT 2206.705 1688.000 2206.995 1688.045 ;
        RECT 2264.190 1688.000 2264.510 1688.060 ;
        RECT 2206.705 1687.860 2264.510 1688.000 ;
        RECT 2206.705 1687.815 2206.995 1687.860 ;
        RECT 2264.190 1687.800 2264.510 1687.860 ;
        RECT 2173.110 1684.940 2173.430 1685.000 ;
        RECT 2206.705 1684.940 2206.995 1684.985 ;
        RECT 2173.110 1684.800 2206.995 1684.940 ;
        RECT 2173.110 1684.740 2173.430 1684.800 ;
        RECT 2206.705 1684.755 2206.995 1684.800 ;
        RECT 2167.590 20.640 2167.910 20.700 ;
        RECT 2173.110 20.640 2173.430 20.700 ;
        RECT 2167.590 20.500 2173.430 20.640 ;
        RECT 2167.590 20.440 2167.910 20.500 ;
        RECT 2173.110 20.440 2173.430 20.500 ;
      LAYER via ;
        RECT 2264.220 1687.800 2264.480 1688.060 ;
        RECT 2173.140 1684.740 2173.400 1685.000 ;
        RECT 2167.620 20.440 2167.880 20.700 ;
        RECT 2173.140 20.440 2173.400 20.700 ;
      LAYER met2 ;
        RECT 2264.140 1700.000 2264.420 1704.000 ;
        RECT 2264.280 1688.090 2264.420 1700.000 ;
        RECT 2264.220 1687.770 2264.480 1688.090 ;
        RECT 2173.140 1684.710 2173.400 1685.030 ;
        RECT 2173.200 20.730 2173.340 1684.710 ;
        RECT 2167.620 20.410 2167.880 20.730 ;
        RECT 2173.140 20.410 2173.400 20.730 ;
        RECT 2167.680 2.400 2167.820 20.410 ;
        RECT 2167.470 -4.800 2168.030 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2211.750 1688.680 2212.070 1688.740 ;
        RECT 2273.390 1688.680 2273.710 1688.740 ;
        RECT 2211.750 1688.540 2273.710 1688.680 ;
        RECT 2211.750 1688.480 2212.070 1688.540 ;
        RECT 2273.390 1688.480 2273.710 1688.540 ;
        RECT 2185.070 20.640 2185.390 20.700 ;
        RECT 2211.750 20.640 2212.070 20.700 ;
        RECT 2185.070 20.500 2212.070 20.640 ;
        RECT 2185.070 20.440 2185.390 20.500 ;
        RECT 2211.750 20.440 2212.070 20.500 ;
      LAYER via ;
        RECT 2211.780 1688.480 2212.040 1688.740 ;
        RECT 2273.420 1688.480 2273.680 1688.740 ;
        RECT 2185.100 20.440 2185.360 20.700 ;
        RECT 2211.780 20.440 2212.040 20.700 ;
      LAYER met2 ;
        RECT 2273.340 1700.000 2273.620 1704.000 ;
        RECT 2273.480 1688.770 2273.620 1700.000 ;
        RECT 2211.780 1688.450 2212.040 1688.770 ;
        RECT 2273.420 1688.450 2273.680 1688.770 ;
        RECT 2211.840 20.730 2211.980 1688.450 ;
        RECT 2185.100 20.410 2185.360 20.730 ;
        RECT 2211.780 20.410 2212.040 20.730 ;
        RECT 2185.160 2.400 2185.300 20.410 ;
        RECT 2184.950 -4.800 2185.510 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2225.090 1689.020 2225.410 1689.080 ;
        RECT 2282.590 1689.020 2282.910 1689.080 ;
        RECT 2225.090 1688.880 2282.910 1689.020 ;
        RECT 2225.090 1688.820 2225.410 1688.880 ;
        RECT 2282.590 1688.820 2282.910 1688.880 ;
        RECT 2203.010 20.300 2203.330 20.360 ;
        RECT 2225.090 20.300 2225.410 20.360 ;
        RECT 2203.010 20.160 2225.410 20.300 ;
        RECT 2203.010 20.100 2203.330 20.160 ;
        RECT 2225.090 20.100 2225.410 20.160 ;
      LAYER via ;
        RECT 2225.120 1688.820 2225.380 1689.080 ;
        RECT 2282.620 1688.820 2282.880 1689.080 ;
        RECT 2203.040 20.100 2203.300 20.360 ;
        RECT 2225.120 20.100 2225.380 20.360 ;
      LAYER met2 ;
        RECT 2282.540 1700.000 2282.820 1704.000 ;
        RECT 2282.680 1689.110 2282.820 1700.000 ;
        RECT 2225.120 1688.790 2225.380 1689.110 ;
        RECT 2282.620 1688.790 2282.880 1689.110 ;
        RECT 2225.180 20.390 2225.320 1688.790 ;
        RECT 2203.040 20.070 2203.300 20.390 ;
        RECT 2225.120 20.070 2225.380 20.390 ;
        RECT 2203.100 2.400 2203.240 20.070 ;
        RECT 2202.890 -4.800 2203.450 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2232.450 1687.320 2232.770 1687.380 ;
        RECT 2291.790 1687.320 2292.110 1687.380 ;
        RECT 2232.450 1687.180 2292.110 1687.320 ;
        RECT 2232.450 1687.120 2232.770 1687.180 ;
        RECT 2291.790 1687.120 2292.110 1687.180 ;
        RECT 2220.950 15.540 2221.270 15.600 ;
        RECT 2232.450 15.540 2232.770 15.600 ;
        RECT 2220.950 15.400 2232.770 15.540 ;
        RECT 2220.950 15.340 2221.270 15.400 ;
        RECT 2232.450 15.340 2232.770 15.400 ;
      LAYER via ;
        RECT 2232.480 1687.120 2232.740 1687.380 ;
        RECT 2291.820 1687.120 2292.080 1687.380 ;
        RECT 2220.980 15.340 2221.240 15.600 ;
        RECT 2232.480 15.340 2232.740 15.600 ;
      LAYER met2 ;
        RECT 2291.740 1700.000 2292.020 1704.000 ;
        RECT 2291.880 1687.410 2292.020 1700.000 ;
        RECT 2232.480 1687.090 2232.740 1687.410 ;
        RECT 2291.820 1687.090 2292.080 1687.410 ;
        RECT 2232.540 15.630 2232.680 1687.090 ;
        RECT 2220.980 15.310 2221.240 15.630 ;
        RECT 2232.480 15.310 2232.740 15.630 ;
        RECT 2221.040 2.400 2221.180 15.310 ;
        RECT 2220.830 -4.800 2221.390 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 779.310 68.240 779.630 68.300 ;
        RECT 1545.670 68.240 1545.990 68.300 ;
        RECT 779.310 68.100 1545.990 68.240 ;
        RECT 779.310 68.040 779.630 68.100 ;
        RECT 1545.670 68.040 1545.990 68.100 ;
      LAYER via ;
        RECT 779.340 68.040 779.600 68.300 ;
        RECT 1545.700 68.040 1545.960 68.300 ;
      LAYER met2 ;
        RECT 1547.920 1700.410 1548.200 1704.000 ;
        RECT 1545.760 1700.270 1548.200 1700.410 ;
        RECT 1545.760 68.330 1545.900 1700.270 ;
        RECT 1547.920 1700.000 1548.200 1700.270 ;
        RECT 779.340 68.010 779.600 68.330 ;
        RECT 1545.700 68.010 1545.960 68.330 ;
        RECT 779.400 16.730 779.540 68.010 ;
        RECT 775.720 16.590 779.540 16.730 ;
        RECT 775.720 2.400 775.860 16.590 ;
        RECT 775.510 -4.800 776.070 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2242.110 1686.300 2242.430 1686.360 ;
        RECT 2300.990 1686.300 2301.310 1686.360 ;
        RECT 2242.110 1686.160 2301.310 1686.300 ;
        RECT 2242.110 1686.100 2242.430 1686.160 ;
        RECT 2300.990 1686.100 2301.310 1686.160 ;
        RECT 2238.890 16.560 2239.210 16.620 ;
        RECT 2242.110 16.560 2242.430 16.620 ;
        RECT 2238.890 16.420 2242.430 16.560 ;
        RECT 2238.890 16.360 2239.210 16.420 ;
        RECT 2242.110 16.360 2242.430 16.420 ;
      LAYER via ;
        RECT 2242.140 1686.100 2242.400 1686.360 ;
        RECT 2301.020 1686.100 2301.280 1686.360 ;
        RECT 2238.920 16.360 2239.180 16.620 ;
        RECT 2242.140 16.360 2242.400 16.620 ;
      LAYER met2 ;
        RECT 2300.940 1700.000 2301.220 1704.000 ;
        RECT 2301.080 1686.390 2301.220 1700.000 ;
        RECT 2242.140 1686.070 2242.400 1686.390 ;
        RECT 2301.020 1686.070 2301.280 1686.390 ;
        RECT 2242.200 16.650 2242.340 1686.070 ;
        RECT 2238.920 16.330 2239.180 16.650 ;
        RECT 2242.140 16.330 2242.400 16.650 ;
        RECT 2238.980 2.400 2239.120 16.330 ;
        RECT 2238.770 -4.800 2239.330 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2266.950 1689.700 2267.270 1689.760 ;
        RECT 2310.190 1689.700 2310.510 1689.760 ;
        RECT 2266.950 1689.560 2310.510 1689.700 ;
        RECT 2266.950 1689.500 2267.270 1689.560 ;
        RECT 2310.190 1689.500 2310.510 1689.560 ;
        RECT 2256.370 20.640 2256.690 20.700 ;
        RECT 2266.950 20.640 2267.270 20.700 ;
        RECT 2256.370 20.500 2267.270 20.640 ;
        RECT 2256.370 20.440 2256.690 20.500 ;
        RECT 2266.950 20.440 2267.270 20.500 ;
      LAYER via ;
        RECT 2266.980 1689.500 2267.240 1689.760 ;
        RECT 2310.220 1689.500 2310.480 1689.760 ;
        RECT 2256.400 20.440 2256.660 20.700 ;
        RECT 2266.980 20.440 2267.240 20.700 ;
      LAYER met2 ;
        RECT 2310.140 1700.000 2310.420 1704.000 ;
        RECT 2310.280 1689.790 2310.420 1700.000 ;
        RECT 2266.980 1689.470 2267.240 1689.790 ;
        RECT 2310.220 1689.470 2310.480 1689.790 ;
        RECT 2267.040 20.730 2267.180 1689.470 ;
        RECT 2256.400 20.410 2256.660 20.730 ;
        RECT 2266.980 20.410 2267.240 20.730 ;
        RECT 2256.460 2.400 2256.600 20.410 ;
        RECT 2256.250 -4.800 2256.810 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2280.290 1688.340 2280.610 1688.400 ;
        RECT 2319.390 1688.340 2319.710 1688.400 ;
        RECT 2280.290 1688.200 2319.710 1688.340 ;
        RECT 2280.290 1688.140 2280.610 1688.200 ;
        RECT 2319.390 1688.140 2319.710 1688.200 ;
        RECT 2274.310 20.300 2274.630 20.360 ;
        RECT 2280.290 20.300 2280.610 20.360 ;
        RECT 2274.310 20.160 2280.610 20.300 ;
        RECT 2274.310 20.100 2274.630 20.160 ;
        RECT 2280.290 20.100 2280.610 20.160 ;
      LAYER via ;
        RECT 2280.320 1688.140 2280.580 1688.400 ;
        RECT 2319.420 1688.140 2319.680 1688.400 ;
        RECT 2274.340 20.100 2274.600 20.360 ;
        RECT 2280.320 20.100 2280.580 20.360 ;
      LAYER met2 ;
        RECT 2319.340 1700.000 2319.620 1704.000 ;
        RECT 2319.480 1688.430 2319.620 1700.000 ;
        RECT 2280.320 1688.110 2280.580 1688.430 ;
        RECT 2319.420 1688.110 2319.680 1688.430 ;
        RECT 2280.380 20.390 2280.520 1688.110 ;
        RECT 2274.340 20.070 2274.600 20.390 ;
        RECT 2280.320 20.070 2280.580 20.390 ;
        RECT 2274.400 2.400 2274.540 20.070 ;
        RECT 2274.190 -4.800 2274.750 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2322.150 1683.920 2322.470 1683.980 ;
        RECT 2328.590 1683.920 2328.910 1683.980 ;
        RECT 2322.150 1683.780 2328.910 1683.920 ;
        RECT 2322.150 1683.720 2322.470 1683.780 ;
        RECT 2328.590 1683.720 2328.910 1683.780 ;
        RECT 2292.250 18.260 2292.570 18.320 ;
        RECT 2322.150 18.260 2322.470 18.320 ;
        RECT 2292.250 18.120 2322.470 18.260 ;
        RECT 2292.250 18.060 2292.570 18.120 ;
        RECT 2322.150 18.060 2322.470 18.120 ;
      LAYER via ;
        RECT 2322.180 1683.720 2322.440 1683.980 ;
        RECT 2328.620 1683.720 2328.880 1683.980 ;
        RECT 2292.280 18.060 2292.540 18.320 ;
        RECT 2322.180 18.060 2322.440 18.320 ;
      LAYER met2 ;
        RECT 2328.540 1700.000 2328.820 1704.000 ;
        RECT 2328.680 1684.010 2328.820 1700.000 ;
        RECT 2322.180 1683.690 2322.440 1684.010 ;
        RECT 2328.620 1683.690 2328.880 1684.010 ;
        RECT 2322.240 18.350 2322.380 1683.690 ;
        RECT 2292.280 18.030 2292.540 18.350 ;
        RECT 2322.180 18.030 2322.440 18.350 ;
        RECT 2292.340 2.400 2292.480 18.030 ;
        RECT 2292.130 -4.800 2292.690 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2332.805 1594.005 2332.975 1608.115 ;
        RECT 2332.805 1497.445 2332.975 1545.555 ;
        RECT 2332.805 1352.605 2332.975 1400.715 ;
        RECT 2332.805 1256.045 2332.975 1304.155 ;
        RECT 2332.805 786.505 2332.975 821.015 ;
        RECT 2332.805 689.605 2332.975 724.455 ;
        RECT 2333.265 572.645 2333.435 620.755 ;
        RECT 2332.345 385.645 2332.515 427.635 ;
        RECT 2332.805 241.485 2332.975 289.595 ;
      LAYER mcon ;
        RECT 2332.805 1607.945 2332.975 1608.115 ;
        RECT 2332.805 1545.385 2332.975 1545.555 ;
        RECT 2332.805 1400.545 2332.975 1400.715 ;
        RECT 2332.805 1303.985 2332.975 1304.155 ;
        RECT 2332.805 820.845 2332.975 821.015 ;
        RECT 2332.805 724.285 2332.975 724.455 ;
        RECT 2333.265 620.585 2333.435 620.755 ;
        RECT 2332.345 427.465 2332.515 427.635 ;
        RECT 2332.805 289.425 2332.975 289.595 ;
      LAYER met1 ;
        RECT 2332.730 1666.580 2333.050 1666.640 ;
        RECT 2335.490 1666.580 2335.810 1666.640 ;
        RECT 2332.730 1666.440 2335.810 1666.580 ;
        RECT 2332.730 1666.380 2333.050 1666.440 ;
        RECT 2335.490 1666.380 2335.810 1666.440 ;
        RECT 2332.730 1608.100 2333.050 1608.160 ;
        RECT 2332.535 1607.960 2333.050 1608.100 ;
        RECT 2332.730 1607.900 2333.050 1607.960 ;
        RECT 2332.730 1594.160 2333.050 1594.220 ;
        RECT 2332.535 1594.020 2333.050 1594.160 ;
        RECT 2332.730 1593.960 2333.050 1594.020 ;
        RECT 2332.270 1559.140 2332.590 1559.200 ;
        RECT 2333.190 1559.140 2333.510 1559.200 ;
        RECT 2332.270 1559.000 2333.510 1559.140 ;
        RECT 2332.270 1558.940 2332.590 1559.000 ;
        RECT 2333.190 1558.940 2333.510 1559.000 ;
        RECT 2332.745 1545.540 2333.035 1545.585 ;
        RECT 2333.190 1545.540 2333.510 1545.600 ;
        RECT 2332.745 1545.400 2333.510 1545.540 ;
        RECT 2332.745 1545.355 2333.035 1545.400 ;
        RECT 2333.190 1545.340 2333.510 1545.400 ;
        RECT 2332.730 1497.600 2333.050 1497.660 ;
        RECT 2332.535 1497.460 2333.050 1497.600 ;
        RECT 2332.730 1497.400 2333.050 1497.460 ;
        RECT 2332.270 1462.580 2332.590 1462.640 ;
        RECT 2333.190 1462.580 2333.510 1462.640 ;
        RECT 2332.270 1462.440 2333.510 1462.580 ;
        RECT 2332.270 1462.380 2332.590 1462.440 ;
        RECT 2333.190 1462.380 2333.510 1462.440 ;
        RECT 2332.730 1400.700 2333.050 1400.760 ;
        RECT 2332.535 1400.560 2333.050 1400.700 ;
        RECT 2332.730 1400.500 2333.050 1400.560 ;
        RECT 2332.745 1352.760 2333.035 1352.805 ;
        RECT 2333.190 1352.760 2333.510 1352.820 ;
        RECT 2332.745 1352.620 2333.510 1352.760 ;
        RECT 2332.745 1352.575 2333.035 1352.620 ;
        RECT 2333.190 1352.560 2333.510 1352.620 ;
        RECT 2332.730 1304.140 2333.050 1304.200 ;
        RECT 2332.535 1304.000 2333.050 1304.140 ;
        RECT 2332.730 1303.940 2333.050 1304.000 ;
        RECT 2332.745 1256.200 2333.035 1256.245 ;
        RECT 2333.190 1256.200 2333.510 1256.260 ;
        RECT 2332.745 1256.060 2333.510 1256.200 ;
        RECT 2332.745 1256.015 2333.035 1256.060 ;
        RECT 2333.190 1256.000 2333.510 1256.060 ;
        RECT 2332.730 1207.240 2333.050 1207.300 ;
        RECT 2333.190 1207.240 2333.510 1207.300 ;
        RECT 2332.730 1207.100 2333.510 1207.240 ;
        RECT 2332.730 1207.040 2333.050 1207.100 ;
        RECT 2333.190 1207.040 2333.510 1207.100 ;
        RECT 2332.730 1110.680 2333.050 1110.740 ;
        RECT 2333.190 1110.680 2333.510 1110.740 ;
        RECT 2332.730 1110.540 2333.510 1110.680 ;
        RECT 2332.730 1110.480 2333.050 1110.540 ;
        RECT 2333.190 1110.480 2333.510 1110.540 ;
        RECT 2332.270 835.280 2332.590 835.340 ;
        RECT 2333.190 835.280 2333.510 835.340 ;
        RECT 2332.270 835.140 2333.510 835.280 ;
        RECT 2332.270 835.080 2332.590 835.140 ;
        RECT 2333.190 835.080 2333.510 835.140 ;
        RECT 2332.730 821.000 2333.050 821.060 ;
        RECT 2332.535 820.860 2333.050 821.000 ;
        RECT 2332.730 820.800 2333.050 820.860 ;
        RECT 2332.730 786.660 2333.050 786.720 ;
        RECT 2332.535 786.520 2333.050 786.660 ;
        RECT 2332.730 786.460 2333.050 786.520 ;
        RECT 2332.270 738.380 2332.590 738.440 ;
        RECT 2333.190 738.380 2333.510 738.440 ;
        RECT 2332.270 738.240 2333.510 738.380 ;
        RECT 2332.270 738.180 2332.590 738.240 ;
        RECT 2333.190 738.180 2333.510 738.240 ;
        RECT 2332.730 724.440 2333.050 724.500 ;
        RECT 2332.535 724.300 2333.050 724.440 ;
        RECT 2332.730 724.240 2333.050 724.300 ;
        RECT 2332.730 689.760 2333.050 689.820 ;
        RECT 2332.535 689.620 2333.050 689.760 ;
        RECT 2332.730 689.560 2333.050 689.620 ;
        RECT 2333.190 620.740 2333.510 620.800 ;
        RECT 2332.995 620.600 2333.510 620.740 ;
        RECT 2333.190 620.540 2333.510 620.600 ;
        RECT 2333.205 572.800 2333.495 572.845 ;
        RECT 2334.110 572.800 2334.430 572.860 ;
        RECT 2333.205 572.660 2334.430 572.800 ;
        RECT 2333.205 572.615 2333.495 572.660 ;
        RECT 2334.110 572.600 2334.430 572.660 ;
        RECT 2332.730 476.240 2333.050 476.300 ;
        RECT 2334.110 476.240 2334.430 476.300 ;
        RECT 2332.730 476.100 2334.430 476.240 ;
        RECT 2332.730 476.040 2333.050 476.100 ;
        RECT 2334.110 476.040 2334.430 476.100 ;
        RECT 2332.730 435.100 2333.050 435.160 ;
        RECT 2333.190 435.100 2333.510 435.160 ;
        RECT 2332.730 434.960 2333.510 435.100 ;
        RECT 2332.730 434.900 2333.050 434.960 ;
        RECT 2333.190 434.900 2333.510 434.960 ;
        RECT 2332.270 427.620 2332.590 427.680 ;
        RECT 2332.075 427.480 2332.590 427.620 ;
        RECT 2332.270 427.420 2332.590 427.480 ;
        RECT 2332.285 385.800 2332.575 385.845 ;
        RECT 2332.730 385.800 2333.050 385.860 ;
        RECT 2332.285 385.660 2333.050 385.800 ;
        RECT 2332.285 385.615 2332.575 385.660 ;
        RECT 2332.730 385.600 2333.050 385.660 ;
        RECT 2332.745 289.580 2333.035 289.625 ;
        RECT 2333.190 289.580 2333.510 289.640 ;
        RECT 2332.745 289.440 2333.510 289.580 ;
        RECT 2332.745 289.395 2333.035 289.440 ;
        RECT 2333.190 289.380 2333.510 289.440 ;
        RECT 2332.730 241.640 2333.050 241.700 ;
        RECT 2332.535 241.500 2333.050 241.640 ;
        RECT 2332.730 241.440 2333.050 241.500 ;
        RECT 2310.190 14.520 2310.510 14.580 ;
        RECT 2333.650 14.520 2333.970 14.580 ;
        RECT 2310.190 14.380 2333.970 14.520 ;
        RECT 2310.190 14.320 2310.510 14.380 ;
        RECT 2333.650 14.320 2333.970 14.380 ;
      LAYER via ;
        RECT 2332.760 1666.380 2333.020 1666.640 ;
        RECT 2335.520 1666.380 2335.780 1666.640 ;
        RECT 2332.760 1607.900 2333.020 1608.160 ;
        RECT 2332.760 1593.960 2333.020 1594.220 ;
        RECT 2332.300 1558.940 2332.560 1559.200 ;
        RECT 2333.220 1558.940 2333.480 1559.200 ;
        RECT 2333.220 1545.340 2333.480 1545.600 ;
        RECT 2332.760 1497.400 2333.020 1497.660 ;
        RECT 2332.300 1462.380 2332.560 1462.640 ;
        RECT 2333.220 1462.380 2333.480 1462.640 ;
        RECT 2332.760 1400.500 2333.020 1400.760 ;
        RECT 2333.220 1352.560 2333.480 1352.820 ;
        RECT 2332.760 1303.940 2333.020 1304.200 ;
        RECT 2333.220 1256.000 2333.480 1256.260 ;
        RECT 2332.760 1207.040 2333.020 1207.300 ;
        RECT 2333.220 1207.040 2333.480 1207.300 ;
        RECT 2332.760 1110.480 2333.020 1110.740 ;
        RECT 2333.220 1110.480 2333.480 1110.740 ;
        RECT 2332.300 835.080 2332.560 835.340 ;
        RECT 2333.220 835.080 2333.480 835.340 ;
        RECT 2332.760 820.800 2333.020 821.060 ;
        RECT 2332.760 786.460 2333.020 786.720 ;
        RECT 2332.300 738.180 2332.560 738.440 ;
        RECT 2333.220 738.180 2333.480 738.440 ;
        RECT 2332.760 724.240 2333.020 724.500 ;
        RECT 2332.760 689.560 2333.020 689.820 ;
        RECT 2333.220 620.540 2333.480 620.800 ;
        RECT 2334.140 572.600 2334.400 572.860 ;
        RECT 2332.760 476.040 2333.020 476.300 ;
        RECT 2334.140 476.040 2334.400 476.300 ;
        RECT 2332.760 434.900 2333.020 435.160 ;
        RECT 2333.220 434.900 2333.480 435.160 ;
        RECT 2332.300 427.420 2332.560 427.680 ;
        RECT 2332.760 385.600 2333.020 385.860 ;
        RECT 2333.220 289.380 2333.480 289.640 ;
        RECT 2332.760 241.440 2333.020 241.700 ;
        RECT 2310.220 14.320 2310.480 14.580 ;
        RECT 2333.680 14.320 2333.940 14.580 ;
      LAYER met2 ;
        RECT 2337.740 1700.410 2338.020 1704.000 ;
        RECT 2335.580 1700.270 2338.020 1700.410 ;
        RECT 2335.580 1666.670 2335.720 1700.270 ;
        RECT 2337.740 1700.000 2338.020 1700.270 ;
        RECT 2332.760 1666.350 2333.020 1666.670 ;
        RECT 2335.520 1666.350 2335.780 1666.670 ;
        RECT 2332.820 1608.190 2332.960 1666.350 ;
        RECT 2332.760 1607.870 2333.020 1608.190 ;
        RECT 2332.760 1593.930 2333.020 1594.250 ;
        RECT 2332.820 1559.650 2332.960 1593.930 ;
        RECT 2332.360 1559.510 2332.960 1559.650 ;
        RECT 2332.360 1559.230 2332.500 1559.510 ;
        RECT 2332.300 1558.910 2332.560 1559.230 ;
        RECT 2333.220 1558.910 2333.480 1559.230 ;
        RECT 2333.280 1545.630 2333.420 1558.910 ;
        RECT 2333.220 1545.310 2333.480 1545.630 ;
        RECT 2332.760 1497.370 2333.020 1497.690 ;
        RECT 2332.820 1463.090 2332.960 1497.370 ;
        RECT 2332.360 1462.950 2332.960 1463.090 ;
        RECT 2332.360 1462.670 2332.500 1462.950 ;
        RECT 2332.300 1462.350 2332.560 1462.670 ;
        RECT 2333.220 1462.350 2333.480 1462.670 ;
        RECT 2333.280 1401.210 2333.420 1462.350 ;
        RECT 2332.820 1401.070 2333.420 1401.210 ;
        RECT 2332.820 1400.790 2332.960 1401.070 ;
        RECT 2332.760 1400.470 2333.020 1400.790 ;
        RECT 2333.220 1352.530 2333.480 1352.850 ;
        RECT 2333.280 1317.570 2333.420 1352.530 ;
        RECT 2332.820 1317.430 2333.420 1317.570 ;
        RECT 2332.820 1304.230 2332.960 1317.430 ;
        RECT 2332.760 1303.910 2333.020 1304.230 ;
        RECT 2333.220 1255.970 2333.480 1256.290 ;
        RECT 2333.280 1221.010 2333.420 1255.970 ;
        RECT 2332.820 1220.870 2333.420 1221.010 ;
        RECT 2332.820 1207.330 2332.960 1220.870 ;
        RECT 2332.760 1207.010 2333.020 1207.330 ;
        RECT 2333.220 1207.010 2333.480 1207.330 ;
        RECT 2333.280 1124.450 2333.420 1207.010 ;
        RECT 2332.820 1124.310 2333.420 1124.450 ;
        RECT 2332.820 1110.770 2332.960 1124.310 ;
        RECT 2332.760 1110.450 2333.020 1110.770 ;
        RECT 2333.220 1110.450 2333.480 1110.770 ;
        RECT 2333.280 1027.890 2333.420 1110.450 ;
        RECT 2332.820 1027.750 2333.420 1027.890 ;
        RECT 2332.820 980.290 2332.960 1027.750 ;
        RECT 2332.360 980.150 2332.960 980.290 ;
        RECT 2332.360 979.610 2332.500 980.150 ;
        RECT 2332.360 979.470 2332.960 979.610 ;
        RECT 2332.820 932.010 2332.960 979.470 ;
        RECT 2332.820 931.870 2333.420 932.010 ;
        RECT 2333.280 835.370 2333.420 931.870 ;
        RECT 2332.300 835.050 2332.560 835.370 ;
        RECT 2333.220 835.050 2333.480 835.370 ;
        RECT 2332.360 834.770 2332.500 835.050 ;
        RECT 2332.360 834.630 2332.960 834.770 ;
        RECT 2332.820 821.090 2332.960 834.630 ;
        RECT 2332.760 820.770 2333.020 821.090 ;
        RECT 2332.760 786.430 2333.020 786.750 ;
        RECT 2332.820 772.890 2332.960 786.430 ;
        RECT 2332.820 772.750 2333.420 772.890 ;
        RECT 2333.280 738.470 2333.420 772.750 ;
        RECT 2332.300 738.210 2332.560 738.470 ;
        RECT 2332.300 738.150 2332.960 738.210 ;
        RECT 2333.220 738.150 2333.480 738.470 ;
        RECT 2332.360 738.070 2332.960 738.150 ;
        RECT 2332.820 724.530 2332.960 738.070 ;
        RECT 2332.760 724.210 2333.020 724.530 ;
        RECT 2332.760 689.530 2333.020 689.850 ;
        RECT 2332.820 676.330 2332.960 689.530 ;
        RECT 2332.820 676.190 2333.420 676.330 ;
        RECT 2333.280 620.830 2333.420 676.190 ;
        RECT 2333.220 620.510 2333.480 620.830 ;
        RECT 2334.140 572.570 2334.400 572.890 ;
        RECT 2334.200 476.330 2334.340 572.570 ;
        RECT 2332.760 476.010 2333.020 476.330 ;
        RECT 2334.140 476.010 2334.400 476.330 ;
        RECT 2332.820 449.210 2332.960 476.010 ;
        RECT 2332.820 449.070 2333.420 449.210 ;
        RECT 2333.280 435.190 2333.420 449.070 ;
        RECT 2332.760 434.930 2333.020 435.190 ;
        RECT 2332.360 434.870 2333.020 434.930 ;
        RECT 2333.220 434.870 2333.480 435.190 ;
        RECT 2332.360 434.790 2332.960 434.870 ;
        RECT 2332.360 427.710 2332.500 434.790 ;
        RECT 2332.300 427.390 2332.560 427.710 ;
        RECT 2332.760 385.570 2333.020 385.890 ;
        RECT 2332.820 303.690 2332.960 385.570 ;
        RECT 2332.820 303.550 2333.420 303.690 ;
        RECT 2333.280 289.670 2333.420 303.550 ;
        RECT 2333.220 289.350 2333.480 289.670 ;
        RECT 2332.760 241.410 2333.020 241.730 ;
        RECT 2332.820 207.130 2332.960 241.410 ;
        RECT 2332.820 206.990 2333.420 207.130 ;
        RECT 2333.280 62.290 2333.420 206.990 ;
        RECT 2333.280 62.150 2333.880 62.290 ;
        RECT 2333.740 14.610 2333.880 62.150 ;
        RECT 2310.220 14.290 2310.480 14.610 ;
        RECT 2333.680 14.290 2333.940 14.610 ;
        RECT 2310.280 2.400 2310.420 14.290 ;
        RECT 2310.070 -4.800 2310.630 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2331.810 1688.340 2332.130 1688.400 ;
        RECT 2346.990 1688.340 2347.310 1688.400 ;
        RECT 2331.810 1688.200 2347.310 1688.340 ;
        RECT 2331.810 1688.140 2332.130 1688.200 ;
        RECT 2346.990 1688.140 2347.310 1688.200 ;
        RECT 2328.130 17.580 2328.450 17.640 ;
        RECT 2331.810 17.580 2332.130 17.640 ;
        RECT 2328.130 17.440 2332.130 17.580 ;
        RECT 2328.130 17.380 2328.450 17.440 ;
        RECT 2331.810 17.380 2332.130 17.440 ;
      LAYER via ;
        RECT 2331.840 1688.140 2332.100 1688.400 ;
        RECT 2347.020 1688.140 2347.280 1688.400 ;
        RECT 2328.160 17.380 2328.420 17.640 ;
        RECT 2331.840 17.380 2332.100 17.640 ;
      LAYER met2 ;
        RECT 2346.940 1700.000 2347.220 1704.000 ;
        RECT 2347.080 1688.430 2347.220 1700.000 ;
        RECT 2331.840 1688.110 2332.100 1688.430 ;
        RECT 2347.020 1688.110 2347.280 1688.430 ;
        RECT 2331.900 17.670 2332.040 1688.110 ;
        RECT 2328.160 17.350 2328.420 17.670 ;
        RECT 2331.840 17.350 2332.100 17.670 ;
        RECT 2328.220 2.400 2328.360 17.350 ;
        RECT 2328.010 -4.800 2328.570 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2349.290 1683.920 2349.610 1683.980 ;
        RECT 2356.190 1683.920 2356.510 1683.980 ;
        RECT 2349.290 1683.780 2356.510 1683.920 ;
        RECT 2349.290 1683.720 2349.610 1683.780 ;
        RECT 2356.190 1683.720 2356.510 1683.780 ;
        RECT 2345.610 20.640 2345.930 20.700 ;
        RECT 2349.290 20.640 2349.610 20.700 ;
        RECT 2345.610 20.500 2349.610 20.640 ;
        RECT 2345.610 20.440 2345.930 20.500 ;
        RECT 2349.290 20.440 2349.610 20.500 ;
      LAYER via ;
        RECT 2349.320 1683.720 2349.580 1683.980 ;
        RECT 2356.220 1683.720 2356.480 1683.980 ;
        RECT 2345.640 20.440 2345.900 20.700 ;
        RECT 2349.320 20.440 2349.580 20.700 ;
      LAYER met2 ;
        RECT 2356.140 1700.000 2356.420 1704.000 ;
        RECT 2356.280 1684.010 2356.420 1700.000 ;
        RECT 2349.320 1683.690 2349.580 1684.010 ;
        RECT 2356.220 1683.690 2356.480 1684.010 ;
        RECT 2349.380 20.730 2349.520 1683.690 ;
        RECT 2345.640 20.410 2345.900 20.730 ;
        RECT 2349.320 20.410 2349.580 20.730 ;
        RECT 2345.700 2.400 2345.840 20.410 ;
        RECT 2345.490 -4.800 2346.050 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2360.405 1594.005 2360.575 1642.115 ;
        RECT 2360.405 1497.445 2360.575 1545.555 ;
        RECT 2360.405 1352.605 2360.575 1400.715 ;
        RECT 2360.405 1256.045 2360.575 1304.155 ;
        RECT 2360.405 338.045 2360.575 427.635 ;
        RECT 2360.405 241.485 2360.575 289.595 ;
        RECT 2360.865 155.805 2361.035 193.035 ;
        RECT 2360.865 96.645 2361.035 111.435 ;
      LAYER mcon ;
        RECT 2360.405 1641.945 2360.575 1642.115 ;
        RECT 2360.405 1545.385 2360.575 1545.555 ;
        RECT 2360.405 1400.545 2360.575 1400.715 ;
        RECT 2360.405 1303.985 2360.575 1304.155 ;
        RECT 2360.405 427.465 2360.575 427.635 ;
        RECT 2360.405 289.425 2360.575 289.595 ;
        RECT 2360.865 192.865 2361.035 193.035 ;
        RECT 2360.865 111.265 2361.035 111.435 ;
      LAYER met1 ;
        RECT 2360.345 1642.100 2360.635 1642.145 ;
        RECT 2360.790 1642.100 2361.110 1642.160 ;
        RECT 2360.345 1641.960 2361.110 1642.100 ;
        RECT 2360.345 1641.915 2360.635 1641.960 ;
        RECT 2360.790 1641.900 2361.110 1641.960 ;
        RECT 2360.330 1594.160 2360.650 1594.220 ;
        RECT 2360.135 1594.020 2360.650 1594.160 ;
        RECT 2360.330 1593.960 2360.650 1594.020 ;
        RECT 2359.870 1559.140 2360.190 1559.200 ;
        RECT 2360.790 1559.140 2361.110 1559.200 ;
        RECT 2359.870 1559.000 2361.110 1559.140 ;
        RECT 2359.870 1558.940 2360.190 1559.000 ;
        RECT 2360.790 1558.940 2361.110 1559.000 ;
        RECT 2360.345 1545.540 2360.635 1545.585 ;
        RECT 2360.790 1545.540 2361.110 1545.600 ;
        RECT 2360.345 1545.400 2361.110 1545.540 ;
        RECT 2360.345 1545.355 2360.635 1545.400 ;
        RECT 2360.790 1545.340 2361.110 1545.400 ;
        RECT 2360.330 1497.600 2360.650 1497.660 ;
        RECT 2360.135 1497.460 2360.650 1497.600 ;
        RECT 2360.330 1497.400 2360.650 1497.460 ;
        RECT 2359.870 1462.580 2360.190 1462.640 ;
        RECT 2360.790 1462.580 2361.110 1462.640 ;
        RECT 2359.870 1462.440 2361.110 1462.580 ;
        RECT 2359.870 1462.380 2360.190 1462.440 ;
        RECT 2360.790 1462.380 2361.110 1462.440 ;
        RECT 2360.330 1400.700 2360.650 1400.760 ;
        RECT 2360.135 1400.560 2360.650 1400.700 ;
        RECT 2360.330 1400.500 2360.650 1400.560 ;
        RECT 2360.345 1352.760 2360.635 1352.805 ;
        RECT 2360.790 1352.760 2361.110 1352.820 ;
        RECT 2360.345 1352.620 2361.110 1352.760 ;
        RECT 2360.345 1352.575 2360.635 1352.620 ;
        RECT 2360.790 1352.560 2361.110 1352.620 ;
        RECT 2360.330 1304.140 2360.650 1304.200 ;
        RECT 2360.135 1304.000 2360.650 1304.140 ;
        RECT 2360.330 1303.940 2360.650 1304.000 ;
        RECT 2360.345 1256.200 2360.635 1256.245 ;
        RECT 2360.790 1256.200 2361.110 1256.260 ;
        RECT 2360.345 1256.060 2361.110 1256.200 ;
        RECT 2360.345 1256.015 2360.635 1256.060 ;
        RECT 2360.790 1256.000 2361.110 1256.060 ;
        RECT 2360.790 1159.300 2361.110 1159.360 ;
        RECT 2361.710 1159.300 2362.030 1159.360 ;
        RECT 2360.790 1159.160 2362.030 1159.300 ;
        RECT 2360.790 1159.100 2361.110 1159.160 ;
        RECT 2361.710 1159.100 2362.030 1159.160 ;
        RECT 2360.790 1062.740 2361.110 1062.800 ;
        RECT 2361.710 1062.740 2362.030 1062.800 ;
        RECT 2360.790 1062.600 2362.030 1062.740 ;
        RECT 2360.790 1062.540 2361.110 1062.600 ;
        RECT 2361.710 1062.540 2362.030 1062.600 ;
        RECT 2360.790 966.180 2361.110 966.240 ;
        RECT 2361.710 966.180 2362.030 966.240 ;
        RECT 2360.790 966.040 2362.030 966.180 ;
        RECT 2360.790 965.980 2361.110 966.040 ;
        RECT 2361.710 965.980 2362.030 966.040 ;
        RECT 2360.790 869.620 2361.110 869.680 ;
        RECT 2361.710 869.620 2362.030 869.680 ;
        RECT 2360.790 869.480 2362.030 869.620 ;
        RECT 2360.790 869.420 2361.110 869.480 ;
        RECT 2361.710 869.420 2362.030 869.480 ;
        RECT 2360.330 821.000 2360.650 821.060 ;
        RECT 2361.710 821.000 2362.030 821.060 ;
        RECT 2360.330 820.860 2362.030 821.000 ;
        RECT 2360.330 820.800 2360.650 820.860 ;
        RECT 2361.710 820.800 2362.030 820.860 ;
        RECT 2360.330 689.900 2360.650 690.160 ;
        RECT 2359.870 689.760 2360.190 689.820 ;
        RECT 2360.420 689.760 2360.560 689.900 ;
        RECT 2359.870 689.620 2360.560 689.760 ;
        RECT 2359.870 689.560 2360.190 689.620 ;
        RECT 2360.330 593.340 2360.650 593.600 ;
        RECT 2359.870 593.200 2360.190 593.260 ;
        RECT 2360.420 593.200 2360.560 593.340 ;
        RECT 2359.870 593.060 2360.560 593.200 ;
        RECT 2359.870 593.000 2360.190 593.060 ;
        RECT 2360.330 496.780 2360.650 497.040 ;
        RECT 2359.870 496.640 2360.190 496.700 ;
        RECT 2360.420 496.640 2360.560 496.780 ;
        RECT 2359.870 496.500 2360.560 496.640 ;
        RECT 2359.870 496.440 2360.190 496.500 ;
        RECT 2360.330 427.620 2360.650 427.680 ;
        RECT 2360.135 427.480 2360.650 427.620 ;
        RECT 2360.330 427.420 2360.650 427.480 ;
        RECT 2360.330 338.200 2360.650 338.260 ;
        RECT 2360.135 338.060 2360.650 338.200 ;
        RECT 2360.330 338.000 2360.650 338.060 ;
        RECT 2359.870 303.520 2360.190 303.580 ;
        RECT 2360.790 303.520 2361.110 303.580 ;
        RECT 2359.870 303.380 2361.110 303.520 ;
        RECT 2359.870 303.320 2360.190 303.380 ;
        RECT 2360.790 303.320 2361.110 303.380 ;
        RECT 2360.345 289.580 2360.635 289.625 ;
        RECT 2360.790 289.580 2361.110 289.640 ;
        RECT 2360.345 289.440 2361.110 289.580 ;
        RECT 2360.345 289.395 2360.635 289.440 ;
        RECT 2360.790 289.380 2361.110 289.440 ;
        RECT 2360.330 241.640 2360.650 241.700 ;
        RECT 2360.135 241.500 2360.650 241.640 ;
        RECT 2360.330 241.440 2360.650 241.500 ;
        RECT 2359.870 206.960 2360.190 207.020 ;
        RECT 2360.790 206.960 2361.110 207.020 ;
        RECT 2359.870 206.820 2361.110 206.960 ;
        RECT 2359.870 206.760 2360.190 206.820 ;
        RECT 2360.790 206.760 2361.110 206.820 ;
        RECT 2360.790 193.020 2361.110 193.080 ;
        RECT 2360.595 192.880 2361.110 193.020 ;
        RECT 2360.790 192.820 2361.110 192.880 ;
        RECT 2360.790 155.960 2361.110 156.020 ;
        RECT 2360.595 155.820 2361.110 155.960 ;
        RECT 2360.790 155.760 2361.110 155.820 ;
        RECT 2360.790 111.420 2361.110 111.480 ;
        RECT 2360.595 111.280 2361.110 111.420 ;
        RECT 2360.790 111.220 2361.110 111.280 ;
        RECT 2360.790 96.800 2361.110 96.860 ;
        RECT 2360.595 96.660 2361.110 96.800 ;
        RECT 2360.790 96.600 2361.110 96.660 ;
        RECT 2360.790 20.640 2361.110 20.700 ;
        RECT 2363.550 20.640 2363.870 20.700 ;
        RECT 2360.790 20.500 2363.870 20.640 ;
        RECT 2360.790 20.440 2361.110 20.500 ;
        RECT 2363.550 20.440 2363.870 20.500 ;
      LAYER via ;
        RECT 2360.820 1641.900 2361.080 1642.160 ;
        RECT 2360.360 1593.960 2360.620 1594.220 ;
        RECT 2359.900 1558.940 2360.160 1559.200 ;
        RECT 2360.820 1558.940 2361.080 1559.200 ;
        RECT 2360.820 1545.340 2361.080 1545.600 ;
        RECT 2360.360 1497.400 2360.620 1497.660 ;
        RECT 2359.900 1462.380 2360.160 1462.640 ;
        RECT 2360.820 1462.380 2361.080 1462.640 ;
        RECT 2360.360 1400.500 2360.620 1400.760 ;
        RECT 2360.820 1352.560 2361.080 1352.820 ;
        RECT 2360.360 1303.940 2360.620 1304.200 ;
        RECT 2360.820 1256.000 2361.080 1256.260 ;
        RECT 2360.820 1159.100 2361.080 1159.360 ;
        RECT 2361.740 1159.100 2362.000 1159.360 ;
        RECT 2360.820 1062.540 2361.080 1062.800 ;
        RECT 2361.740 1062.540 2362.000 1062.800 ;
        RECT 2360.820 965.980 2361.080 966.240 ;
        RECT 2361.740 965.980 2362.000 966.240 ;
        RECT 2360.820 869.420 2361.080 869.680 ;
        RECT 2361.740 869.420 2362.000 869.680 ;
        RECT 2360.360 820.800 2360.620 821.060 ;
        RECT 2361.740 820.800 2362.000 821.060 ;
        RECT 2360.360 689.900 2360.620 690.160 ;
        RECT 2359.900 689.560 2360.160 689.820 ;
        RECT 2360.360 593.340 2360.620 593.600 ;
        RECT 2359.900 593.000 2360.160 593.260 ;
        RECT 2360.360 496.780 2360.620 497.040 ;
        RECT 2359.900 496.440 2360.160 496.700 ;
        RECT 2360.360 427.420 2360.620 427.680 ;
        RECT 2360.360 338.000 2360.620 338.260 ;
        RECT 2359.900 303.320 2360.160 303.580 ;
        RECT 2360.820 303.320 2361.080 303.580 ;
        RECT 2360.820 289.380 2361.080 289.640 ;
        RECT 2360.360 241.440 2360.620 241.700 ;
        RECT 2359.900 206.760 2360.160 207.020 ;
        RECT 2360.820 206.760 2361.080 207.020 ;
        RECT 2360.820 192.820 2361.080 193.080 ;
        RECT 2360.820 155.760 2361.080 156.020 ;
        RECT 2360.820 111.220 2361.080 111.480 ;
        RECT 2360.820 96.600 2361.080 96.860 ;
        RECT 2360.820 20.440 2361.080 20.700 ;
        RECT 2363.580 20.440 2363.840 20.700 ;
      LAYER met2 ;
        RECT 2365.340 1700.410 2365.620 1704.000 ;
        RECT 2362.720 1700.270 2365.620 1700.410 ;
        RECT 2362.720 1666.410 2362.860 1700.270 ;
        RECT 2365.340 1700.000 2365.620 1700.270 ;
        RECT 2360.880 1666.270 2362.860 1666.410 ;
        RECT 2360.880 1642.190 2361.020 1666.270 ;
        RECT 2360.820 1641.870 2361.080 1642.190 ;
        RECT 2360.360 1593.930 2360.620 1594.250 ;
        RECT 2360.420 1559.650 2360.560 1593.930 ;
        RECT 2359.960 1559.510 2360.560 1559.650 ;
        RECT 2359.960 1559.230 2360.100 1559.510 ;
        RECT 2359.900 1558.910 2360.160 1559.230 ;
        RECT 2360.820 1558.910 2361.080 1559.230 ;
        RECT 2360.880 1545.630 2361.020 1558.910 ;
        RECT 2360.820 1545.310 2361.080 1545.630 ;
        RECT 2360.360 1497.370 2360.620 1497.690 ;
        RECT 2360.420 1463.090 2360.560 1497.370 ;
        RECT 2359.960 1462.950 2360.560 1463.090 ;
        RECT 2359.960 1462.670 2360.100 1462.950 ;
        RECT 2359.900 1462.350 2360.160 1462.670 ;
        RECT 2360.820 1462.350 2361.080 1462.670 ;
        RECT 2360.880 1401.210 2361.020 1462.350 ;
        RECT 2360.420 1401.070 2361.020 1401.210 ;
        RECT 2360.420 1400.790 2360.560 1401.070 ;
        RECT 2360.360 1400.470 2360.620 1400.790 ;
        RECT 2360.820 1352.530 2361.080 1352.850 ;
        RECT 2360.880 1317.570 2361.020 1352.530 ;
        RECT 2360.420 1317.430 2361.020 1317.570 ;
        RECT 2360.420 1304.230 2360.560 1317.430 ;
        RECT 2360.360 1303.910 2360.620 1304.230 ;
        RECT 2360.820 1255.970 2361.080 1256.290 ;
        RECT 2360.880 1221.010 2361.020 1255.970 ;
        RECT 2360.420 1220.870 2361.020 1221.010 ;
        RECT 2360.420 1207.525 2360.560 1220.870 ;
        RECT 2360.350 1207.155 2360.630 1207.525 ;
        RECT 2361.730 1207.155 2362.010 1207.525 ;
        RECT 2361.800 1159.390 2361.940 1207.155 ;
        RECT 2360.820 1159.070 2361.080 1159.390 ;
        RECT 2361.740 1159.070 2362.000 1159.390 ;
        RECT 2360.880 1124.450 2361.020 1159.070 ;
        RECT 2360.420 1124.310 2361.020 1124.450 ;
        RECT 2360.420 1110.965 2360.560 1124.310 ;
        RECT 2360.350 1110.595 2360.630 1110.965 ;
        RECT 2361.730 1110.595 2362.010 1110.965 ;
        RECT 2361.800 1062.830 2361.940 1110.595 ;
        RECT 2360.820 1062.510 2361.080 1062.830 ;
        RECT 2361.740 1062.510 2362.000 1062.830 ;
        RECT 2360.880 1027.890 2361.020 1062.510 ;
        RECT 2360.420 1027.750 2361.020 1027.890 ;
        RECT 2360.420 1014.405 2360.560 1027.750 ;
        RECT 2360.350 1014.035 2360.630 1014.405 ;
        RECT 2361.730 1014.035 2362.010 1014.405 ;
        RECT 2361.800 966.270 2361.940 1014.035 ;
        RECT 2360.820 965.950 2361.080 966.270 ;
        RECT 2361.740 965.950 2362.000 966.270 ;
        RECT 2360.880 931.330 2361.020 965.950 ;
        RECT 2360.420 931.190 2361.020 931.330 ;
        RECT 2360.420 917.845 2360.560 931.190 ;
        RECT 2360.350 917.475 2360.630 917.845 ;
        RECT 2361.730 917.475 2362.010 917.845 ;
        RECT 2361.800 869.710 2361.940 917.475 ;
        RECT 2360.820 869.390 2361.080 869.710 ;
        RECT 2361.740 869.390 2362.000 869.710 ;
        RECT 2360.880 834.770 2361.020 869.390 ;
        RECT 2360.420 834.630 2361.020 834.770 ;
        RECT 2360.420 821.090 2360.560 834.630 ;
        RECT 2360.360 820.770 2360.620 821.090 ;
        RECT 2361.740 820.770 2362.000 821.090 ;
        RECT 2361.800 773.005 2361.940 820.770 ;
        RECT 2360.810 772.635 2361.090 773.005 ;
        RECT 2361.730 772.635 2362.010 773.005 ;
        RECT 2360.880 738.210 2361.020 772.635 ;
        RECT 2360.420 738.070 2361.020 738.210 ;
        RECT 2360.420 690.190 2360.560 738.070 ;
        RECT 2360.360 689.870 2360.620 690.190 ;
        RECT 2359.900 689.530 2360.160 689.850 ;
        RECT 2359.960 676.445 2360.100 689.530 ;
        RECT 2359.890 676.075 2360.170 676.445 ;
        RECT 2360.810 676.075 2361.090 676.445 ;
        RECT 2360.880 641.650 2361.020 676.075 ;
        RECT 2360.420 641.510 2361.020 641.650 ;
        RECT 2360.420 593.630 2360.560 641.510 ;
        RECT 2360.360 593.310 2360.620 593.630 ;
        RECT 2359.900 592.970 2360.160 593.290 ;
        RECT 2359.960 579.885 2360.100 592.970 ;
        RECT 2359.890 579.515 2360.170 579.885 ;
        RECT 2360.810 579.515 2361.090 579.885 ;
        RECT 2360.880 545.090 2361.020 579.515 ;
        RECT 2360.420 544.950 2361.020 545.090 ;
        RECT 2360.420 497.070 2360.560 544.950 ;
        RECT 2360.360 496.750 2360.620 497.070 ;
        RECT 2359.900 496.410 2360.160 496.730 ;
        RECT 2359.960 483.325 2360.100 496.410 ;
        RECT 2359.890 482.955 2360.170 483.325 ;
        RECT 2360.810 482.955 2361.090 483.325 ;
        RECT 2360.880 448.530 2361.020 482.955 ;
        RECT 2360.420 448.390 2361.020 448.530 ;
        RECT 2360.420 427.710 2360.560 448.390 ;
        RECT 2360.360 427.390 2360.620 427.710 ;
        RECT 2360.360 337.970 2360.620 338.290 ;
        RECT 2360.420 303.690 2360.560 337.970 ;
        RECT 2359.960 303.610 2360.560 303.690 ;
        RECT 2359.900 303.550 2360.560 303.610 ;
        RECT 2359.900 303.290 2360.160 303.550 ;
        RECT 2360.820 303.290 2361.080 303.610 ;
        RECT 2360.880 289.670 2361.020 303.290 ;
        RECT 2360.820 289.350 2361.080 289.670 ;
        RECT 2360.360 241.410 2360.620 241.730 ;
        RECT 2360.420 207.130 2360.560 241.410 ;
        RECT 2359.960 207.050 2360.560 207.130 ;
        RECT 2359.900 206.990 2360.560 207.050 ;
        RECT 2359.900 206.730 2360.160 206.990 ;
        RECT 2360.820 206.730 2361.080 207.050 ;
        RECT 2360.880 193.110 2361.020 206.730 ;
        RECT 2360.820 192.790 2361.080 193.110 ;
        RECT 2360.820 155.730 2361.080 156.050 ;
        RECT 2360.880 111.510 2361.020 155.730 ;
        RECT 2360.820 111.190 2361.080 111.510 ;
        RECT 2360.820 96.570 2361.080 96.890 ;
        RECT 2360.880 20.730 2361.020 96.570 ;
        RECT 2360.820 20.410 2361.080 20.730 ;
        RECT 2363.580 20.410 2363.840 20.730 ;
        RECT 2363.640 2.400 2363.780 20.410 ;
        RECT 2363.430 -4.800 2363.990 2.400 ;
      LAYER via2 ;
        RECT 2360.350 1207.200 2360.630 1207.480 ;
        RECT 2361.730 1207.200 2362.010 1207.480 ;
        RECT 2360.350 1110.640 2360.630 1110.920 ;
        RECT 2361.730 1110.640 2362.010 1110.920 ;
        RECT 2360.350 1014.080 2360.630 1014.360 ;
        RECT 2361.730 1014.080 2362.010 1014.360 ;
        RECT 2360.350 917.520 2360.630 917.800 ;
        RECT 2361.730 917.520 2362.010 917.800 ;
        RECT 2360.810 772.680 2361.090 772.960 ;
        RECT 2361.730 772.680 2362.010 772.960 ;
        RECT 2359.890 676.120 2360.170 676.400 ;
        RECT 2360.810 676.120 2361.090 676.400 ;
        RECT 2359.890 579.560 2360.170 579.840 ;
        RECT 2360.810 579.560 2361.090 579.840 ;
        RECT 2359.890 483.000 2360.170 483.280 ;
        RECT 2360.810 483.000 2361.090 483.280 ;
      LAYER met3 ;
        RECT 2360.325 1207.490 2360.655 1207.505 ;
        RECT 2361.705 1207.490 2362.035 1207.505 ;
        RECT 2360.325 1207.190 2362.035 1207.490 ;
        RECT 2360.325 1207.175 2360.655 1207.190 ;
        RECT 2361.705 1207.175 2362.035 1207.190 ;
        RECT 2360.325 1110.930 2360.655 1110.945 ;
        RECT 2361.705 1110.930 2362.035 1110.945 ;
        RECT 2360.325 1110.630 2362.035 1110.930 ;
        RECT 2360.325 1110.615 2360.655 1110.630 ;
        RECT 2361.705 1110.615 2362.035 1110.630 ;
        RECT 2360.325 1014.370 2360.655 1014.385 ;
        RECT 2361.705 1014.370 2362.035 1014.385 ;
        RECT 2360.325 1014.070 2362.035 1014.370 ;
        RECT 2360.325 1014.055 2360.655 1014.070 ;
        RECT 2361.705 1014.055 2362.035 1014.070 ;
        RECT 2360.325 917.810 2360.655 917.825 ;
        RECT 2361.705 917.810 2362.035 917.825 ;
        RECT 2360.325 917.510 2362.035 917.810 ;
        RECT 2360.325 917.495 2360.655 917.510 ;
        RECT 2361.705 917.495 2362.035 917.510 ;
        RECT 2360.785 772.970 2361.115 772.985 ;
        RECT 2361.705 772.970 2362.035 772.985 ;
        RECT 2360.785 772.670 2362.035 772.970 ;
        RECT 2360.785 772.655 2361.115 772.670 ;
        RECT 2361.705 772.655 2362.035 772.670 ;
        RECT 2359.865 676.410 2360.195 676.425 ;
        RECT 2360.785 676.410 2361.115 676.425 ;
        RECT 2359.865 676.110 2361.115 676.410 ;
        RECT 2359.865 676.095 2360.195 676.110 ;
        RECT 2360.785 676.095 2361.115 676.110 ;
        RECT 2359.865 579.850 2360.195 579.865 ;
        RECT 2360.785 579.850 2361.115 579.865 ;
        RECT 2359.865 579.550 2361.115 579.850 ;
        RECT 2359.865 579.535 2360.195 579.550 ;
        RECT 2360.785 579.535 2361.115 579.550 ;
        RECT 2359.865 483.290 2360.195 483.305 ;
        RECT 2360.785 483.290 2361.115 483.305 ;
        RECT 2359.865 482.990 2361.115 483.290 ;
        RECT 2359.865 482.975 2360.195 482.990 ;
        RECT 2360.785 482.975 2361.115 482.990 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2374.590 1683.920 2374.910 1683.980 ;
        RECT 2380.110 1683.920 2380.430 1683.980 ;
        RECT 2374.590 1683.780 2380.430 1683.920 ;
        RECT 2374.590 1683.720 2374.910 1683.780 ;
        RECT 2380.110 1683.720 2380.430 1683.780 ;
      LAYER via ;
        RECT 2374.620 1683.720 2374.880 1683.980 ;
        RECT 2380.140 1683.720 2380.400 1683.980 ;
      LAYER met2 ;
        RECT 2374.540 1700.000 2374.820 1704.000 ;
        RECT 2374.680 1684.010 2374.820 1700.000 ;
        RECT 2374.620 1683.690 2374.880 1684.010 ;
        RECT 2380.140 1683.690 2380.400 1684.010 ;
        RECT 2380.200 18.090 2380.340 1683.690 ;
        RECT 2380.200 17.950 2381.720 18.090 ;
        RECT 2381.580 2.400 2381.720 17.950 ;
        RECT 2381.370 -4.800 2381.930 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2383.790 1684.600 2384.110 1684.660 ;
        RECT 2387.010 1684.600 2387.330 1684.660 ;
        RECT 2383.790 1684.460 2387.330 1684.600 ;
        RECT 2383.790 1684.400 2384.110 1684.460 ;
        RECT 2387.010 1684.400 2387.330 1684.460 ;
        RECT 2387.010 20.300 2387.330 20.360 ;
        RECT 2399.430 20.300 2399.750 20.360 ;
        RECT 2387.010 20.160 2399.750 20.300 ;
        RECT 2387.010 20.100 2387.330 20.160 ;
        RECT 2399.430 20.100 2399.750 20.160 ;
      LAYER via ;
        RECT 2383.820 1684.400 2384.080 1684.660 ;
        RECT 2387.040 1684.400 2387.300 1684.660 ;
        RECT 2387.040 20.100 2387.300 20.360 ;
        RECT 2399.460 20.100 2399.720 20.360 ;
      LAYER met2 ;
        RECT 2383.740 1700.000 2384.020 1704.000 ;
        RECT 2383.880 1684.690 2384.020 1700.000 ;
        RECT 2383.820 1684.370 2384.080 1684.690 ;
        RECT 2387.040 1684.370 2387.300 1684.690 ;
        RECT 2387.100 20.390 2387.240 1684.370 ;
        RECT 2387.040 20.070 2387.300 20.390 ;
        RECT 2399.460 20.070 2399.720 20.390 ;
        RECT 2399.520 2.400 2399.660 20.070 ;
        RECT 2399.310 -4.800 2399.870 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1553.565 1449.165 1553.735 1497.275 ;
        RECT 1553.565 1352.605 1553.735 1400.715 ;
        RECT 1553.565 1256.045 1553.735 1304.155 ;
        RECT 1553.565 593.045 1553.735 627.895 ;
        RECT 1553.565 483.225 1553.735 496.995 ;
        RECT 1553.565 386.325 1553.735 434.775 ;
        RECT 1553.105 276.165 1553.275 324.275 ;
      LAYER mcon ;
        RECT 1553.565 1497.105 1553.735 1497.275 ;
        RECT 1553.565 1400.545 1553.735 1400.715 ;
        RECT 1553.565 1303.985 1553.735 1304.155 ;
        RECT 1553.565 627.725 1553.735 627.895 ;
        RECT 1553.565 496.825 1553.735 496.995 ;
        RECT 1553.565 434.605 1553.735 434.775 ;
        RECT 1553.105 324.105 1553.275 324.275 ;
      LAYER met1 ;
        RECT 1553.490 1678.140 1553.810 1678.200 ;
        RECT 1555.790 1678.140 1556.110 1678.200 ;
        RECT 1553.490 1678.000 1556.110 1678.140 ;
        RECT 1553.490 1677.940 1553.810 1678.000 ;
        RECT 1555.790 1677.940 1556.110 1678.000 ;
        RECT 1553.490 1497.260 1553.810 1497.320 ;
        RECT 1553.295 1497.120 1553.810 1497.260 ;
        RECT 1553.490 1497.060 1553.810 1497.120 ;
        RECT 1553.490 1449.320 1553.810 1449.380 ;
        RECT 1553.295 1449.180 1553.810 1449.320 ;
        RECT 1553.490 1449.120 1553.810 1449.180 ;
        RECT 1553.490 1400.700 1553.810 1400.760 ;
        RECT 1553.295 1400.560 1553.810 1400.700 ;
        RECT 1553.490 1400.500 1553.810 1400.560 ;
        RECT 1553.490 1352.760 1553.810 1352.820 ;
        RECT 1553.295 1352.620 1553.810 1352.760 ;
        RECT 1553.490 1352.560 1553.810 1352.620 ;
        RECT 1553.490 1304.140 1553.810 1304.200 ;
        RECT 1553.295 1304.000 1553.810 1304.140 ;
        RECT 1553.490 1303.940 1553.810 1304.000 ;
        RECT 1553.490 1256.200 1553.810 1256.260 ;
        RECT 1553.295 1256.060 1553.810 1256.200 ;
        RECT 1553.490 1256.000 1553.810 1256.060 ;
        RECT 1553.490 1159.300 1553.810 1159.360 ;
        RECT 1554.410 1159.300 1554.730 1159.360 ;
        RECT 1553.490 1159.160 1554.730 1159.300 ;
        RECT 1553.490 1159.100 1553.810 1159.160 ;
        RECT 1554.410 1159.100 1554.730 1159.160 ;
        RECT 1553.490 1062.740 1553.810 1062.800 ;
        RECT 1554.410 1062.740 1554.730 1062.800 ;
        RECT 1553.490 1062.600 1554.730 1062.740 ;
        RECT 1553.490 1062.540 1553.810 1062.600 ;
        RECT 1554.410 1062.540 1554.730 1062.600 ;
        RECT 1553.490 869.620 1553.810 869.680 ;
        RECT 1554.410 869.620 1554.730 869.680 ;
        RECT 1553.490 869.480 1554.730 869.620 ;
        RECT 1553.490 869.420 1553.810 869.480 ;
        RECT 1554.410 869.420 1554.730 869.480 ;
        RECT 1553.490 821.000 1553.810 821.060 ;
        RECT 1554.410 821.000 1554.730 821.060 ;
        RECT 1553.490 820.860 1554.730 821.000 ;
        RECT 1553.490 820.800 1553.810 820.860 ;
        RECT 1554.410 820.800 1554.730 820.860 ;
        RECT 1553.490 627.880 1553.810 627.940 ;
        RECT 1553.295 627.740 1553.810 627.880 ;
        RECT 1553.490 627.680 1553.810 627.740 ;
        RECT 1553.490 593.200 1553.810 593.260 ;
        RECT 1553.295 593.060 1553.810 593.200 ;
        RECT 1553.490 593.000 1553.810 593.060 ;
        RECT 1553.490 496.980 1553.810 497.040 ;
        RECT 1553.295 496.840 1553.810 496.980 ;
        RECT 1553.490 496.780 1553.810 496.840 ;
        RECT 1553.490 483.380 1553.810 483.440 ;
        RECT 1553.295 483.240 1553.810 483.380 ;
        RECT 1553.490 483.180 1553.810 483.240 ;
        RECT 1553.490 434.760 1553.810 434.820 ;
        RECT 1553.295 434.620 1553.810 434.760 ;
        RECT 1553.490 434.560 1553.810 434.620 ;
        RECT 1553.490 386.480 1553.810 386.540 ;
        RECT 1553.295 386.340 1553.810 386.480 ;
        RECT 1553.490 386.280 1553.810 386.340 ;
        RECT 1553.030 338.200 1553.350 338.260 ;
        RECT 1553.490 338.200 1553.810 338.260 ;
        RECT 1553.030 338.060 1553.810 338.200 ;
        RECT 1553.030 338.000 1553.350 338.060 ;
        RECT 1553.490 338.000 1553.810 338.060 ;
        RECT 1553.030 324.260 1553.350 324.320 ;
        RECT 1552.835 324.120 1553.350 324.260 ;
        RECT 1553.030 324.060 1553.350 324.120 ;
        RECT 1553.045 276.320 1553.335 276.365 ;
        RECT 1554.410 276.320 1554.730 276.380 ;
        RECT 1553.045 276.180 1554.730 276.320 ;
        RECT 1553.045 276.135 1553.335 276.180 ;
        RECT 1554.410 276.120 1554.730 276.180 ;
        RECT 1553.030 186.560 1553.350 186.620 ;
        RECT 1553.950 186.560 1554.270 186.620 ;
        RECT 1553.030 186.420 1554.270 186.560 ;
        RECT 1553.030 186.360 1553.350 186.420 ;
        RECT 1553.950 186.360 1554.270 186.420 ;
        RECT 799.550 68.580 799.870 68.640 ;
        RECT 1553.490 68.580 1553.810 68.640 ;
        RECT 799.550 68.440 1553.810 68.580 ;
        RECT 799.550 68.380 799.870 68.440 ;
        RECT 1553.490 68.380 1553.810 68.440 ;
        RECT 793.570 20.980 793.890 21.040 ;
        RECT 799.550 20.980 799.870 21.040 ;
        RECT 793.570 20.840 799.870 20.980 ;
        RECT 793.570 20.780 793.890 20.840 ;
        RECT 799.550 20.780 799.870 20.840 ;
      LAYER via ;
        RECT 1553.520 1677.940 1553.780 1678.200 ;
        RECT 1555.820 1677.940 1556.080 1678.200 ;
        RECT 1553.520 1497.060 1553.780 1497.320 ;
        RECT 1553.520 1449.120 1553.780 1449.380 ;
        RECT 1553.520 1400.500 1553.780 1400.760 ;
        RECT 1553.520 1352.560 1553.780 1352.820 ;
        RECT 1553.520 1303.940 1553.780 1304.200 ;
        RECT 1553.520 1256.000 1553.780 1256.260 ;
        RECT 1553.520 1159.100 1553.780 1159.360 ;
        RECT 1554.440 1159.100 1554.700 1159.360 ;
        RECT 1553.520 1062.540 1553.780 1062.800 ;
        RECT 1554.440 1062.540 1554.700 1062.800 ;
        RECT 1553.520 869.420 1553.780 869.680 ;
        RECT 1554.440 869.420 1554.700 869.680 ;
        RECT 1553.520 820.800 1553.780 821.060 ;
        RECT 1554.440 820.800 1554.700 821.060 ;
        RECT 1553.520 627.680 1553.780 627.940 ;
        RECT 1553.520 593.000 1553.780 593.260 ;
        RECT 1553.520 496.780 1553.780 497.040 ;
        RECT 1553.520 483.180 1553.780 483.440 ;
        RECT 1553.520 434.560 1553.780 434.820 ;
        RECT 1553.520 386.280 1553.780 386.540 ;
        RECT 1553.060 338.000 1553.320 338.260 ;
        RECT 1553.520 338.000 1553.780 338.260 ;
        RECT 1553.060 324.060 1553.320 324.320 ;
        RECT 1554.440 276.120 1554.700 276.380 ;
        RECT 1553.060 186.360 1553.320 186.620 ;
        RECT 1553.980 186.360 1554.240 186.620 ;
        RECT 799.580 68.380 799.840 68.640 ;
        RECT 1553.520 68.380 1553.780 68.640 ;
        RECT 793.600 20.780 793.860 21.040 ;
        RECT 799.580 20.780 799.840 21.040 ;
      LAYER met2 ;
        RECT 1557.120 1700.410 1557.400 1704.000 ;
        RECT 1555.880 1700.270 1557.400 1700.410 ;
        RECT 1555.880 1678.230 1556.020 1700.270 ;
        RECT 1557.120 1700.000 1557.400 1700.270 ;
        RECT 1553.520 1677.910 1553.780 1678.230 ;
        RECT 1555.820 1677.910 1556.080 1678.230 ;
        RECT 1553.580 1559.650 1553.720 1677.910 ;
        RECT 1553.120 1559.510 1553.720 1559.650 ;
        RECT 1553.120 1558.970 1553.260 1559.510 ;
        RECT 1553.120 1558.830 1553.720 1558.970 ;
        RECT 1553.580 1497.350 1553.720 1558.830 ;
        RECT 1553.520 1497.030 1553.780 1497.350 ;
        RECT 1553.520 1449.090 1553.780 1449.410 ;
        RECT 1553.580 1400.790 1553.720 1449.090 ;
        RECT 1553.520 1400.470 1553.780 1400.790 ;
        RECT 1553.520 1352.530 1553.780 1352.850 ;
        RECT 1553.580 1304.230 1553.720 1352.530 ;
        RECT 1553.520 1303.910 1553.780 1304.230 ;
        RECT 1553.520 1255.970 1553.780 1256.290 ;
        RECT 1553.580 1207.525 1553.720 1255.970 ;
        RECT 1553.510 1207.155 1553.790 1207.525 ;
        RECT 1554.430 1207.155 1554.710 1207.525 ;
        RECT 1554.500 1159.390 1554.640 1207.155 ;
        RECT 1553.520 1159.070 1553.780 1159.390 ;
        RECT 1554.440 1159.070 1554.700 1159.390 ;
        RECT 1553.580 1110.965 1553.720 1159.070 ;
        RECT 1553.510 1110.595 1553.790 1110.965 ;
        RECT 1554.430 1110.595 1554.710 1110.965 ;
        RECT 1554.500 1062.830 1554.640 1110.595 ;
        RECT 1553.520 1062.510 1553.780 1062.830 ;
        RECT 1554.440 1062.510 1554.700 1062.830 ;
        RECT 1553.580 980.290 1553.720 1062.510 ;
        RECT 1553.120 980.150 1553.720 980.290 ;
        RECT 1553.120 979.610 1553.260 980.150 ;
        RECT 1553.120 979.470 1553.720 979.610 ;
        RECT 1553.580 917.845 1553.720 979.470 ;
        RECT 1553.510 917.475 1553.790 917.845 ;
        RECT 1554.430 917.475 1554.710 917.845 ;
        RECT 1554.500 869.710 1554.640 917.475 ;
        RECT 1553.520 869.390 1553.780 869.710 ;
        RECT 1554.440 869.390 1554.700 869.710 ;
        RECT 1553.580 821.090 1553.720 869.390 ;
        RECT 1553.520 820.770 1553.780 821.090 ;
        RECT 1554.440 820.770 1554.700 821.090 ;
        RECT 1554.500 773.005 1554.640 820.770 ;
        RECT 1553.510 772.635 1553.790 773.005 ;
        RECT 1554.430 772.635 1554.710 773.005 ;
        RECT 1553.580 690.610 1553.720 772.635 ;
        RECT 1553.120 690.470 1553.720 690.610 ;
        RECT 1553.120 689.930 1553.260 690.470 ;
        RECT 1553.120 689.790 1553.720 689.930 ;
        RECT 1553.580 627.970 1553.720 689.790 ;
        RECT 1553.520 627.650 1553.780 627.970 ;
        RECT 1553.520 592.970 1553.780 593.290 ;
        RECT 1553.580 497.070 1553.720 592.970 ;
        RECT 1553.520 496.750 1553.780 497.070 ;
        RECT 1553.520 483.150 1553.780 483.470 ;
        RECT 1553.580 434.850 1553.720 483.150 ;
        RECT 1553.520 434.530 1553.780 434.850 ;
        RECT 1553.520 386.250 1553.780 386.570 ;
        RECT 1553.580 338.290 1553.720 386.250 ;
        RECT 1553.060 337.970 1553.320 338.290 ;
        RECT 1553.520 337.970 1553.780 338.290 ;
        RECT 1553.120 324.350 1553.260 337.970 ;
        RECT 1553.060 324.030 1553.320 324.350 ;
        RECT 1554.440 276.090 1554.700 276.410 ;
        RECT 1554.500 235.125 1554.640 276.090 ;
        RECT 1554.430 234.755 1554.710 235.125 ;
        RECT 1553.970 233.395 1554.250 233.765 ;
        RECT 1554.040 186.650 1554.180 233.395 ;
        RECT 1553.060 186.330 1553.320 186.650 ;
        RECT 1553.980 186.330 1554.240 186.650 ;
        RECT 1553.120 113.970 1553.260 186.330 ;
        RECT 1553.120 113.830 1553.720 113.970 ;
        RECT 1553.580 68.670 1553.720 113.830 ;
        RECT 799.580 68.350 799.840 68.670 ;
        RECT 1553.520 68.350 1553.780 68.670 ;
        RECT 799.640 21.070 799.780 68.350 ;
        RECT 793.600 20.750 793.860 21.070 ;
        RECT 799.580 20.750 799.840 21.070 ;
        RECT 793.660 2.400 793.800 20.750 ;
        RECT 793.450 -4.800 794.010 2.400 ;
      LAYER via2 ;
        RECT 1553.510 1207.200 1553.790 1207.480 ;
        RECT 1554.430 1207.200 1554.710 1207.480 ;
        RECT 1553.510 1110.640 1553.790 1110.920 ;
        RECT 1554.430 1110.640 1554.710 1110.920 ;
        RECT 1553.510 917.520 1553.790 917.800 ;
        RECT 1554.430 917.520 1554.710 917.800 ;
        RECT 1553.510 772.680 1553.790 772.960 ;
        RECT 1554.430 772.680 1554.710 772.960 ;
        RECT 1554.430 234.800 1554.710 235.080 ;
        RECT 1553.970 233.440 1554.250 233.720 ;
      LAYER met3 ;
        RECT 1553.485 1207.490 1553.815 1207.505 ;
        RECT 1554.405 1207.490 1554.735 1207.505 ;
        RECT 1553.485 1207.190 1554.735 1207.490 ;
        RECT 1553.485 1207.175 1553.815 1207.190 ;
        RECT 1554.405 1207.175 1554.735 1207.190 ;
        RECT 1553.485 1110.930 1553.815 1110.945 ;
        RECT 1554.405 1110.930 1554.735 1110.945 ;
        RECT 1553.485 1110.630 1554.735 1110.930 ;
        RECT 1553.485 1110.615 1553.815 1110.630 ;
        RECT 1554.405 1110.615 1554.735 1110.630 ;
        RECT 1553.485 917.810 1553.815 917.825 ;
        RECT 1554.405 917.810 1554.735 917.825 ;
        RECT 1553.485 917.510 1554.735 917.810 ;
        RECT 1553.485 917.495 1553.815 917.510 ;
        RECT 1554.405 917.495 1554.735 917.510 ;
        RECT 1553.485 772.970 1553.815 772.985 ;
        RECT 1554.405 772.970 1554.735 772.985 ;
        RECT 1553.485 772.670 1554.735 772.970 ;
        RECT 1553.485 772.655 1553.815 772.670 ;
        RECT 1554.405 772.655 1554.735 772.670 ;
        RECT 1554.405 235.090 1554.735 235.105 ;
        RECT 1553.270 234.790 1554.735 235.090 ;
        RECT 1553.270 233.730 1553.570 234.790 ;
        RECT 1554.405 234.775 1554.735 234.790 ;
        RECT 1553.945 233.730 1554.275 233.745 ;
        RECT 1553.270 233.430 1554.275 233.730 ;
        RECT 1553.945 233.415 1554.275 233.430 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 641.310 59.060 641.630 59.120 ;
        RECT 1476.670 59.060 1476.990 59.120 ;
        RECT 641.310 58.920 1476.990 59.060 ;
        RECT 641.310 58.860 641.630 58.920 ;
        RECT 1476.670 58.860 1476.990 58.920 ;
      LAYER via ;
        RECT 641.340 58.860 641.600 59.120 ;
        RECT 1476.700 58.860 1476.960 59.120 ;
      LAYER met2 ;
        RECT 1477.540 1700.410 1477.820 1704.000 ;
        RECT 1476.760 1700.270 1477.820 1700.410 ;
        RECT 1476.760 59.150 1476.900 1700.270 ;
        RECT 1477.540 1700.000 1477.820 1700.270 ;
        RECT 641.340 58.830 641.600 59.150 ;
        RECT 1476.700 58.830 1476.960 59.150 ;
        RECT 641.400 17.410 641.540 58.830 ;
        RECT 639.100 17.270 641.540 17.410 ;
        RECT 639.100 2.400 639.240 17.270 ;
        RECT 638.890 -4.800 639.450 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2395.750 1684.940 2396.070 1685.000 ;
        RECT 2422.890 1684.940 2423.210 1685.000 ;
        RECT 2395.750 1684.800 2423.210 1684.940 ;
        RECT 2395.750 1684.740 2396.070 1684.800 ;
        RECT 2422.890 1684.740 2423.210 1684.800 ;
      LAYER via ;
        RECT 2395.780 1684.740 2396.040 1685.000 ;
        RECT 2422.920 1684.740 2423.180 1685.000 ;
      LAYER met2 ;
        RECT 2395.700 1700.000 2395.980 1704.000 ;
        RECT 2395.840 1685.030 2395.980 1700.000 ;
        RECT 2395.780 1684.710 2396.040 1685.030 ;
        RECT 2422.920 1684.710 2423.180 1685.030 ;
        RECT 2422.980 2.400 2423.120 1684.710 ;
        RECT 2422.770 -4.800 2423.330 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2404.950 1684.260 2405.270 1684.320 ;
        RECT 2425.190 1684.260 2425.510 1684.320 ;
        RECT 2404.950 1684.120 2425.510 1684.260 ;
        RECT 2404.950 1684.060 2405.270 1684.120 ;
        RECT 2425.190 1684.060 2425.510 1684.120 ;
        RECT 2425.190 16.220 2425.510 16.280 ;
        RECT 2440.830 16.220 2441.150 16.280 ;
        RECT 2425.190 16.080 2441.150 16.220 ;
        RECT 2425.190 16.020 2425.510 16.080 ;
        RECT 2440.830 16.020 2441.150 16.080 ;
      LAYER via ;
        RECT 2404.980 1684.060 2405.240 1684.320 ;
        RECT 2425.220 1684.060 2425.480 1684.320 ;
        RECT 2425.220 16.020 2425.480 16.280 ;
        RECT 2440.860 16.020 2441.120 16.280 ;
      LAYER met2 ;
        RECT 2404.900 1700.000 2405.180 1704.000 ;
        RECT 2405.040 1684.350 2405.180 1700.000 ;
        RECT 2404.980 1684.030 2405.240 1684.350 ;
        RECT 2425.220 1684.030 2425.480 1684.350 ;
        RECT 2425.280 16.310 2425.420 1684.030 ;
        RECT 2425.220 15.990 2425.480 16.310 ;
        RECT 2440.860 15.990 2441.120 16.310 ;
        RECT 2440.920 2.400 2441.060 15.990 ;
        RECT 2440.710 -4.800 2441.270 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2414.150 1686.980 2414.470 1687.040 ;
        RECT 2457.390 1686.980 2457.710 1687.040 ;
        RECT 2414.150 1686.840 2457.710 1686.980 ;
        RECT 2414.150 1686.780 2414.470 1686.840 ;
        RECT 2457.390 1686.780 2457.710 1686.840 ;
      LAYER via ;
        RECT 2414.180 1686.780 2414.440 1687.040 ;
        RECT 2457.420 1686.780 2457.680 1687.040 ;
      LAYER met2 ;
        RECT 2414.100 1700.000 2414.380 1704.000 ;
        RECT 2414.240 1687.070 2414.380 1700.000 ;
        RECT 2414.180 1686.750 2414.440 1687.070 ;
        RECT 2457.420 1686.750 2457.680 1687.070 ;
        RECT 2457.480 3.130 2457.620 1686.750 ;
        RECT 2457.480 2.990 2458.540 3.130 ;
        RECT 2458.400 2.960 2458.540 2.990 ;
        RECT 2458.400 2.820 2459.000 2.960 ;
        RECT 2458.860 2.400 2459.000 2.820 ;
        RECT 2458.650 -4.800 2459.210 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2423.350 1683.920 2423.670 1683.980 ;
        RECT 2428.410 1683.920 2428.730 1683.980 ;
        RECT 2423.350 1683.780 2428.730 1683.920 ;
        RECT 2423.350 1683.720 2423.670 1683.780 ;
        RECT 2428.410 1683.720 2428.730 1683.780 ;
        RECT 2428.410 18.600 2428.730 18.660 ;
        RECT 2476.710 18.600 2477.030 18.660 ;
        RECT 2428.410 18.460 2477.030 18.600 ;
        RECT 2428.410 18.400 2428.730 18.460 ;
        RECT 2476.710 18.400 2477.030 18.460 ;
      LAYER via ;
        RECT 2423.380 1683.720 2423.640 1683.980 ;
        RECT 2428.440 1683.720 2428.700 1683.980 ;
        RECT 2428.440 18.400 2428.700 18.660 ;
        RECT 2476.740 18.400 2477.000 18.660 ;
      LAYER met2 ;
        RECT 2423.300 1700.000 2423.580 1704.000 ;
        RECT 2423.440 1684.010 2423.580 1700.000 ;
        RECT 2423.380 1683.690 2423.640 1684.010 ;
        RECT 2428.440 1683.690 2428.700 1684.010 ;
        RECT 2428.500 18.690 2428.640 1683.690 ;
        RECT 2428.440 18.370 2428.700 18.690 ;
        RECT 2476.740 18.370 2477.000 18.690 ;
        RECT 2476.800 2.400 2476.940 18.370 ;
        RECT 2476.590 -4.800 2477.150 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2435.310 17.580 2435.630 17.640 ;
        RECT 2494.650 17.580 2494.970 17.640 ;
        RECT 2435.310 17.440 2494.970 17.580 ;
        RECT 2435.310 17.380 2435.630 17.440 ;
        RECT 2494.650 17.380 2494.970 17.440 ;
      LAYER via ;
        RECT 2435.340 17.380 2435.600 17.640 ;
        RECT 2494.680 17.380 2494.940 17.640 ;
      LAYER met2 ;
        RECT 2432.500 1700.410 2432.780 1704.000 ;
        RECT 2432.500 1700.270 2435.540 1700.410 ;
        RECT 2432.500 1700.000 2432.780 1700.270 ;
        RECT 2435.400 17.670 2435.540 1700.270 ;
        RECT 2435.340 17.350 2435.600 17.670 ;
        RECT 2494.680 17.350 2494.940 17.670 ;
        RECT 2494.740 2.400 2494.880 17.350 ;
        RECT 2494.530 -4.800 2495.090 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2442.210 16.560 2442.530 16.620 ;
        RECT 2512.130 16.560 2512.450 16.620 ;
        RECT 2442.210 16.420 2512.450 16.560 ;
        RECT 2442.210 16.360 2442.530 16.420 ;
        RECT 2512.130 16.360 2512.450 16.420 ;
      LAYER via ;
        RECT 2442.240 16.360 2442.500 16.620 ;
        RECT 2512.160 16.360 2512.420 16.620 ;
      LAYER met2 ;
        RECT 2441.700 1700.410 2441.980 1704.000 ;
        RECT 2441.700 1700.270 2442.440 1700.410 ;
        RECT 2441.700 1700.000 2441.980 1700.270 ;
        RECT 2442.300 16.650 2442.440 1700.270 ;
        RECT 2442.240 16.330 2442.500 16.650 ;
        RECT 2512.160 16.330 2512.420 16.650 ;
        RECT 2512.220 2.400 2512.360 16.330 ;
        RECT 2512.010 -4.800 2512.570 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2450.950 1689.700 2451.270 1689.760 ;
        RECT 2507.990 1689.700 2508.310 1689.760 ;
        RECT 2450.950 1689.560 2508.310 1689.700 ;
        RECT 2450.950 1689.500 2451.270 1689.560 ;
        RECT 2507.990 1689.500 2508.310 1689.560 ;
        RECT 2507.990 15.540 2508.310 15.600 ;
        RECT 2530.070 15.540 2530.390 15.600 ;
        RECT 2507.990 15.400 2530.390 15.540 ;
        RECT 2507.990 15.340 2508.310 15.400 ;
        RECT 2530.070 15.340 2530.390 15.400 ;
      LAYER via ;
        RECT 2450.980 1689.500 2451.240 1689.760 ;
        RECT 2508.020 1689.500 2508.280 1689.760 ;
        RECT 2508.020 15.340 2508.280 15.600 ;
        RECT 2530.100 15.340 2530.360 15.600 ;
      LAYER met2 ;
        RECT 2450.900 1700.000 2451.180 1704.000 ;
        RECT 2451.040 1689.790 2451.180 1700.000 ;
        RECT 2450.980 1689.470 2451.240 1689.790 ;
        RECT 2508.020 1689.470 2508.280 1689.790 ;
        RECT 2508.080 15.630 2508.220 1689.470 ;
        RECT 2508.020 15.310 2508.280 15.630 ;
        RECT 2530.100 15.310 2530.360 15.630 ;
        RECT 2530.160 2.400 2530.300 15.310 ;
        RECT 2529.950 -4.800 2530.510 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2462.910 20.300 2463.230 20.360 ;
        RECT 2548.010 20.300 2548.330 20.360 ;
        RECT 2462.910 20.160 2548.330 20.300 ;
        RECT 2462.910 20.100 2463.230 20.160 ;
        RECT 2548.010 20.100 2548.330 20.160 ;
      LAYER via ;
        RECT 2462.940 20.100 2463.200 20.360 ;
        RECT 2548.040 20.100 2548.300 20.360 ;
      LAYER met2 ;
        RECT 2460.100 1700.410 2460.380 1704.000 ;
        RECT 2460.100 1700.270 2463.140 1700.410 ;
        RECT 2460.100 1700.000 2460.380 1700.270 ;
        RECT 2463.000 20.390 2463.140 1700.270 ;
        RECT 2462.940 20.070 2463.200 20.390 ;
        RECT 2548.040 20.070 2548.300 20.390 ;
        RECT 2548.100 2.400 2548.240 20.070 ;
        RECT 2547.890 -4.800 2548.450 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2469.810 20.640 2470.130 20.700 ;
        RECT 2565.950 20.640 2566.270 20.700 ;
        RECT 2469.810 20.500 2566.270 20.640 ;
        RECT 2469.810 20.440 2470.130 20.500 ;
        RECT 2565.950 20.440 2566.270 20.500 ;
      LAYER via ;
        RECT 2469.840 20.440 2470.100 20.700 ;
        RECT 2565.980 20.440 2566.240 20.700 ;
      LAYER met2 ;
        RECT 2469.300 1700.410 2469.580 1704.000 ;
        RECT 2469.300 1700.270 2470.040 1700.410 ;
        RECT 2469.300 1700.000 2469.580 1700.270 ;
        RECT 2469.900 20.730 2470.040 1700.270 ;
        RECT 2469.840 20.410 2470.100 20.730 ;
        RECT 2565.980 20.410 2566.240 20.730 ;
        RECT 2566.040 2.400 2566.180 20.410 ;
        RECT 2565.830 -4.800 2566.390 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2549.005 16.405 2549.175 19.295 ;
      LAYER mcon ;
        RECT 2549.005 19.125 2549.175 19.295 ;
      LAYER met1 ;
        RECT 2478.550 1686.300 2478.870 1686.360 ;
        RECT 2483.610 1686.300 2483.930 1686.360 ;
        RECT 2478.550 1686.160 2483.930 1686.300 ;
        RECT 2478.550 1686.100 2478.870 1686.160 ;
        RECT 2483.610 1686.100 2483.930 1686.160 ;
        RECT 2483.610 19.280 2483.930 19.340 ;
        RECT 2548.945 19.280 2549.235 19.325 ;
        RECT 2483.610 19.140 2549.235 19.280 ;
        RECT 2483.610 19.080 2483.930 19.140 ;
        RECT 2548.945 19.095 2549.235 19.140 ;
        RECT 2548.945 16.560 2549.235 16.605 ;
        RECT 2583.890 16.560 2584.210 16.620 ;
        RECT 2548.945 16.420 2584.210 16.560 ;
        RECT 2548.945 16.375 2549.235 16.420 ;
        RECT 2583.890 16.360 2584.210 16.420 ;
      LAYER via ;
        RECT 2478.580 1686.100 2478.840 1686.360 ;
        RECT 2483.640 1686.100 2483.900 1686.360 ;
        RECT 2483.640 19.080 2483.900 19.340 ;
        RECT 2583.920 16.360 2584.180 16.620 ;
      LAYER met2 ;
        RECT 2478.500 1700.000 2478.780 1704.000 ;
        RECT 2478.640 1686.390 2478.780 1700.000 ;
        RECT 2478.580 1686.070 2478.840 1686.390 ;
        RECT 2483.640 1686.070 2483.900 1686.390 ;
        RECT 2483.700 19.370 2483.840 1686.070 ;
        RECT 2483.640 19.050 2483.900 19.370 ;
        RECT 2583.920 16.330 2584.180 16.650 ;
        RECT 2583.980 2.400 2584.120 16.330 ;
        RECT 2583.770 -4.800 2584.330 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 817.490 34.240 817.810 34.300 ;
        RECT 1567.750 34.240 1568.070 34.300 ;
        RECT 817.490 34.100 1568.070 34.240 ;
        RECT 817.490 34.040 817.810 34.100 ;
        RECT 1567.750 34.040 1568.070 34.100 ;
      LAYER via ;
        RECT 817.520 34.040 817.780 34.300 ;
        RECT 1567.780 34.040 1568.040 34.300 ;
      LAYER met2 ;
        RECT 1569.080 1700.410 1569.360 1704.000 ;
        RECT 1567.840 1700.270 1569.360 1700.410 ;
        RECT 1567.840 34.330 1567.980 1700.270 ;
        RECT 1569.080 1700.000 1569.360 1700.270 ;
        RECT 817.520 34.010 817.780 34.330 ;
        RECT 1567.780 34.010 1568.040 34.330 ;
        RECT 817.580 2.400 817.720 34.010 ;
        RECT 817.370 -4.800 817.930 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2487.750 1689.360 2488.070 1689.420 ;
        RECT 2549.390 1689.360 2549.710 1689.420 ;
        RECT 2487.750 1689.220 2549.710 1689.360 ;
        RECT 2487.750 1689.160 2488.070 1689.220 ;
        RECT 2549.390 1689.160 2549.710 1689.220 ;
        RECT 2549.390 19.280 2549.710 19.340 ;
        RECT 2601.370 19.280 2601.690 19.340 ;
        RECT 2549.390 19.140 2601.690 19.280 ;
        RECT 2549.390 19.080 2549.710 19.140 ;
        RECT 2601.370 19.080 2601.690 19.140 ;
      LAYER via ;
        RECT 2487.780 1689.160 2488.040 1689.420 ;
        RECT 2549.420 1689.160 2549.680 1689.420 ;
        RECT 2549.420 19.080 2549.680 19.340 ;
        RECT 2601.400 19.080 2601.660 19.340 ;
      LAYER met2 ;
        RECT 2487.700 1700.000 2487.980 1704.000 ;
        RECT 2487.840 1689.450 2487.980 1700.000 ;
        RECT 2487.780 1689.130 2488.040 1689.450 ;
        RECT 2549.420 1689.130 2549.680 1689.450 ;
        RECT 2549.480 19.370 2549.620 1689.130 ;
        RECT 2549.420 19.050 2549.680 19.370 ;
        RECT 2601.400 19.050 2601.660 19.370 ;
        RECT 2601.460 2.400 2601.600 19.050 ;
        RECT 2601.250 -4.800 2601.810 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2496.950 17.920 2497.270 17.980 ;
        RECT 2619.310 17.920 2619.630 17.980 ;
        RECT 2496.950 17.780 2619.630 17.920 ;
        RECT 2496.950 17.720 2497.270 17.780 ;
        RECT 2619.310 17.720 2619.630 17.780 ;
      LAYER via ;
        RECT 2496.980 17.720 2497.240 17.980 ;
        RECT 2619.340 17.720 2619.600 17.980 ;
      LAYER met2 ;
        RECT 2496.900 1700.000 2497.180 1704.000 ;
        RECT 2497.040 18.010 2497.180 1700.000 ;
        RECT 2496.980 17.690 2497.240 18.010 ;
        RECT 2619.340 17.690 2619.600 18.010 ;
        RECT 2619.400 2.400 2619.540 17.690 ;
        RECT 2619.190 -4.800 2619.750 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2526.940 1688.880 2532.600 1689.020 ;
        RECT 2506.150 1688.680 2506.470 1688.740 ;
        RECT 2526.940 1688.680 2527.080 1688.880 ;
        RECT 2506.150 1688.540 2527.080 1688.680 ;
        RECT 2532.460 1688.680 2532.600 1688.880 ;
        RECT 2532.460 1688.540 2565.260 1688.680 ;
        RECT 2506.150 1688.480 2506.470 1688.540 ;
        RECT 2565.120 1688.340 2565.260 1688.540 ;
        RECT 2583.890 1688.340 2584.210 1688.400 ;
        RECT 2565.120 1688.200 2584.210 1688.340 ;
        RECT 2583.890 1688.140 2584.210 1688.200 ;
        RECT 2583.430 14.180 2583.750 14.240 ;
        RECT 2637.250 14.180 2637.570 14.240 ;
        RECT 2583.430 14.040 2637.570 14.180 ;
        RECT 2583.430 13.980 2583.750 14.040 ;
        RECT 2637.250 13.980 2637.570 14.040 ;
      LAYER via ;
        RECT 2506.180 1688.480 2506.440 1688.740 ;
        RECT 2583.920 1688.140 2584.180 1688.400 ;
        RECT 2583.460 13.980 2583.720 14.240 ;
        RECT 2637.280 13.980 2637.540 14.240 ;
      LAYER met2 ;
        RECT 2506.100 1700.000 2506.380 1704.000 ;
        RECT 2506.240 1688.770 2506.380 1700.000 ;
        RECT 2506.180 1688.450 2506.440 1688.770 ;
        RECT 2583.920 1688.110 2584.180 1688.430 ;
        RECT 2583.980 24.380 2584.120 1688.110 ;
        RECT 2583.520 24.240 2584.120 24.380 ;
        RECT 2583.520 14.270 2583.660 24.240 ;
        RECT 2583.460 13.950 2583.720 14.270 ;
        RECT 2637.280 13.950 2637.540 14.270 ;
        RECT 2637.340 2.400 2637.480 13.950 ;
        RECT 2637.130 -4.800 2637.690 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2518.570 14.520 2518.890 14.580 ;
        RECT 2655.190 14.520 2655.510 14.580 ;
        RECT 2518.570 14.380 2655.510 14.520 ;
        RECT 2518.570 14.320 2518.890 14.380 ;
        RECT 2655.190 14.320 2655.510 14.380 ;
      LAYER via ;
        RECT 2518.600 14.320 2518.860 14.580 ;
        RECT 2655.220 14.320 2655.480 14.580 ;
      LAYER met2 ;
        RECT 2515.300 1700.410 2515.580 1704.000 ;
        RECT 2515.300 1700.270 2517.880 1700.410 ;
        RECT 2515.300 1700.000 2515.580 1700.270 ;
        RECT 2517.740 1688.850 2517.880 1700.270 ;
        RECT 2517.740 1688.710 2518.340 1688.850 ;
        RECT 2518.200 17.920 2518.340 1688.710 ;
        RECT 2518.200 17.780 2518.800 17.920 ;
        RECT 2518.660 14.610 2518.800 17.780 ;
        RECT 2518.600 14.290 2518.860 14.610 ;
        RECT 2655.220 14.290 2655.480 14.610 ;
        RECT 2655.280 2.400 2655.420 14.290 ;
        RECT 2655.070 -4.800 2655.630 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2524.550 1684.600 2524.870 1684.660 ;
        RECT 2670.370 1684.600 2670.690 1684.660 ;
        RECT 2524.550 1684.460 2670.690 1684.600 ;
        RECT 2524.550 1684.400 2524.870 1684.460 ;
        RECT 2670.370 1684.400 2670.690 1684.460 ;
      LAYER via ;
        RECT 2524.580 1684.400 2524.840 1684.660 ;
        RECT 2670.400 1684.400 2670.660 1684.660 ;
      LAYER met2 ;
        RECT 2524.500 1700.000 2524.780 1704.000 ;
        RECT 2524.640 1684.690 2524.780 1700.000 ;
        RECT 2524.580 1684.370 2524.840 1684.690 ;
        RECT 2670.400 1684.370 2670.660 1684.690 ;
        RECT 2670.460 16.730 2670.600 1684.370 ;
        RECT 2670.460 16.590 2672.900 16.730 ;
        RECT 2672.760 2.400 2672.900 16.590 ;
        RECT 2672.550 -4.800 2673.110 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2533.750 1686.300 2534.070 1686.360 ;
        RECT 2538.810 1686.300 2539.130 1686.360 ;
        RECT 2533.750 1686.160 2539.130 1686.300 ;
        RECT 2533.750 1686.100 2534.070 1686.160 ;
        RECT 2538.810 1686.100 2539.130 1686.160 ;
        RECT 2538.810 15.540 2539.130 15.600 ;
        RECT 2690.610 15.540 2690.930 15.600 ;
        RECT 2538.810 15.400 2690.930 15.540 ;
        RECT 2538.810 15.340 2539.130 15.400 ;
        RECT 2690.610 15.340 2690.930 15.400 ;
      LAYER via ;
        RECT 2533.780 1686.100 2534.040 1686.360 ;
        RECT 2538.840 1686.100 2539.100 1686.360 ;
        RECT 2538.840 15.340 2539.100 15.600 ;
        RECT 2690.640 15.340 2690.900 15.600 ;
      LAYER met2 ;
        RECT 2533.700 1700.000 2533.980 1704.000 ;
        RECT 2533.840 1686.390 2533.980 1700.000 ;
        RECT 2533.780 1686.070 2534.040 1686.390 ;
        RECT 2538.840 1686.070 2539.100 1686.390 ;
        RECT 2538.900 15.630 2539.040 1686.070 ;
        RECT 2538.840 15.310 2539.100 15.630 ;
        RECT 2690.640 15.310 2690.900 15.630 ;
        RECT 2690.700 2.400 2690.840 15.310 ;
        RECT 2690.490 -4.800 2691.050 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2634.105 1687.505 2634.275 1688.355 ;
      LAYER mcon ;
        RECT 2634.105 1688.185 2634.275 1688.355 ;
      LAYER met1 ;
        RECT 2634.045 1688.340 2634.335 1688.385 ;
        RECT 2597.780 1688.200 2634.335 1688.340 ;
        RECT 2542.950 1688.000 2543.270 1688.060 ;
        RECT 2597.780 1688.000 2597.920 1688.200 ;
        RECT 2634.045 1688.155 2634.335 1688.200 ;
        RECT 2542.950 1687.860 2597.920 1688.000 ;
        RECT 2542.950 1687.800 2543.270 1687.860 ;
        RECT 2634.045 1687.660 2634.335 1687.705 ;
        RECT 2644.610 1687.660 2644.930 1687.720 ;
        RECT 2634.045 1687.520 2644.930 1687.660 ;
        RECT 2634.045 1687.475 2634.335 1687.520 ;
        RECT 2644.610 1687.460 2644.930 1687.520 ;
        RECT 2645.990 14.180 2646.310 14.240 ;
        RECT 2708.550 14.180 2708.870 14.240 ;
        RECT 2645.990 14.040 2708.870 14.180 ;
        RECT 2645.990 13.980 2646.310 14.040 ;
        RECT 2708.550 13.980 2708.870 14.040 ;
      LAYER via ;
        RECT 2542.980 1687.800 2543.240 1688.060 ;
        RECT 2644.640 1687.460 2644.900 1687.720 ;
        RECT 2646.020 13.980 2646.280 14.240 ;
        RECT 2708.580 13.980 2708.840 14.240 ;
      LAYER met2 ;
        RECT 2542.900 1700.000 2543.180 1704.000 ;
        RECT 2543.040 1688.090 2543.180 1700.000 ;
        RECT 2542.980 1687.770 2543.240 1688.090 ;
        RECT 2644.700 1688.030 2646.220 1688.170 ;
        RECT 2644.700 1687.750 2644.840 1688.030 ;
        RECT 2644.640 1687.430 2644.900 1687.750 ;
        RECT 2646.080 14.270 2646.220 1688.030 ;
        RECT 2646.020 13.950 2646.280 14.270 ;
        RECT 2708.580 13.950 2708.840 14.270 ;
        RECT 2708.640 2.400 2708.780 13.950 ;
        RECT 2708.430 -4.800 2708.990 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2584.885 16.065 2585.055 20.315 ;
      LAYER mcon ;
        RECT 2584.885 20.145 2585.055 20.315 ;
      LAYER met1 ;
        RECT 2552.610 20.300 2552.930 20.360 ;
        RECT 2584.825 20.300 2585.115 20.345 ;
        RECT 2552.610 20.160 2585.115 20.300 ;
        RECT 2552.610 20.100 2552.930 20.160 ;
        RECT 2584.825 20.115 2585.115 20.160 ;
        RECT 2584.825 16.220 2585.115 16.265 ;
        RECT 2584.825 16.080 2694.980 16.220 ;
        RECT 2584.825 16.035 2585.115 16.080 ;
        RECT 2694.840 15.880 2694.980 16.080 ;
        RECT 2726.490 15.880 2726.810 15.940 ;
        RECT 2694.840 15.740 2726.810 15.880 ;
        RECT 2726.490 15.680 2726.810 15.740 ;
      LAYER via ;
        RECT 2552.640 20.100 2552.900 20.360 ;
        RECT 2726.520 15.680 2726.780 15.940 ;
      LAYER met2 ;
        RECT 2552.100 1700.410 2552.380 1704.000 ;
        RECT 2552.100 1700.270 2552.840 1700.410 ;
        RECT 2552.100 1700.000 2552.380 1700.270 ;
        RECT 2552.700 20.390 2552.840 1700.270 ;
        RECT 2552.640 20.070 2552.900 20.390 ;
        RECT 2726.520 15.650 2726.780 15.970 ;
        RECT 2726.580 2.400 2726.720 15.650 ;
        RECT 2726.370 -4.800 2726.930 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2561.350 1690.380 2561.670 1690.440 ;
        RECT 2735.690 1690.380 2736.010 1690.440 ;
        RECT 2561.350 1690.240 2736.010 1690.380 ;
        RECT 2561.350 1690.180 2561.670 1690.240 ;
        RECT 2735.690 1690.180 2736.010 1690.240 ;
        RECT 2735.690 15.880 2736.010 15.940 ;
        RECT 2744.430 15.880 2744.750 15.940 ;
        RECT 2735.690 15.740 2744.750 15.880 ;
        RECT 2735.690 15.680 2736.010 15.740 ;
        RECT 2744.430 15.680 2744.750 15.740 ;
      LAYER via ;
        RECT 2561.380 1690.180 2561.640 1690.440 ;
        RECT 2735.720 1690.180 2735.980 1690.440 ;
        RECT 2735.720 15.680 2735.980 15.940 ;
        RECT 2744.460 15.680 2744.720 15.940 ;
      LAYER met2 ;
        RECT 2561.300 1700.000 2561.580 1704.000 ;
        RECT 2561.440 1690.470 2561.580 1700.000 ;
        RECT 2561.380 1690.150 2561.640 1690.470 ;
        RECT 2735.720 1690.150 2735.980 1690.470 ;
        RECT 2735.780 15.970 2735.920 1690.150 ;
        RECT 2735.720 15.650 2735.980 15.970 ;
        RECT 2744.460 15.650 2744.720 15.970 ;
        RECT 2744.520 2.400 2744.660 15.650 ;
        RECT 2744.310 -4.800 2744.870 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2573.310 16.900 2573.630 16.960 ;
        RECT 2761.910 16.900 2762.230 16.960 ;
        RECT 2573.310 16.760 2762.230 16.900 ;
        RECT 2573.310 16.700 2573.630 16.760 ;
        RECT 2761.910 16.700 2762.230 16.760 ;
      LAYER via ;
        RECT 2573.340 16.700 2573.600 16.960 ;
        RECT 2761.940 16.700 2762.200 16.960 ;
      LAYER met2 ;
        RECT 2570.040 1701.090 2570.320 1704.000 ;
        RECT 2570.040 1700.950 2573.080 1701.090 ;
        RECT 2570.040 1700.000 2570.320 1700.950 ;
        RECT 2572.940 1688.340 2573.080 1700.950 ;
        RECT 2572.940 1688.200 2573.540 1688.340 ;
        RECT 2573.400 16.990 2573.540 1688.200 ;
        RECT 2573.340 16.670 2573.600 16.990 ;
        RECT 2761.940 16.670 2762.200 16.990 ;
        RECT 2762.000 2.400 2762.140 16.670 ;
        RECT 2761.790 -4.800 2762.350 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1573.270 1689.360 1573.590 1689.420 ;
        RECT 1576.950 1689.360 1577.270 1689.420 ;
        RECT 1573.270 1689.220 1577.270 1689.360 ;
        RECT 1573.270 1689.160 1573.590 1689.220 ;
        RECT 1576.950 1689.160 1577.270 1689.220 ;
        RECT 835.430 30.500 835.750 30.560 ;
        RECT 1572.810 30.500 1573.130 30.560 ;
        RECT 835.430 30.360 1573.130 30.500 ;
        RECT 835.430 30.300 835.750 30.360 ;
        RECT 1572.810 30.300 1573.130 30.360 ;
      LAYER via ;
        RECT 1573.300 1689.160 1573.560 1689.420 ;
        RECT 1576.980 1689.160 1577.240 1689.420 ;
        RECT 835.460 30.300 835.720 30.560 ;
        RECT 1572.840 30.300 1573.100 30.560 ;
      LAYER met2 ;
        RECT 1578.280 1700.410 1578.560 1704.000 ;
        RECT 1577.040 1700.270 1578.560 1700.410 ;
        RECT 1577.040 1689.450 1577.180 1700.270 ;
        RECT 1578.280 1700.000 1578.560 1700.270 ;
        RECT 1573.300 1689.130 1573.560 1689.450 ;
        RECT 1576.980 1689.130 1577.240 1689.450 ;
        RECT 1573.360 31.010 1573.500 1689.130 ;
        RECT 1572.900 30.870 1573.500 31.010 ;
        RECT 1572.900 30.590 1573.040 30.870 ;
        RECT 835.460 30.270 835.720 30.590 ;
        RECT 1572.840 30.270 1573.100 30.590 ;
        RECT 835.520 2.400 835.660 30.270 ;
        RECT 835.310 -4.800 835.870 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2579.290 1689.020 2579.610 1689.080 ;
        RECT 2774.330 1689.020 2774.650 1689.080 ;
        RECT 2579.290 1688.880 2774.650 1689.020 ;
        RECT 2579.290 1688.820 2579.610 1688.880 ;
        RECT 2774.330 1688.820 2774.650 1688.880 ;
      LAYER via ;
        RECT 2579.320 1688.820 2579.580 1689.080 ;
        RECT 2774.360 1688.820 2774.620 1689.080 ;
      LAYER met2 ;
        RECT 2579.240 1700.000 2579.520 1704.000 ;
        RECT 2579.380 1689.110 2579.520 1700.000 ;
        RECT 2579.320 1688.790 2579.580 1689.110 ;
        RECT 2774.360 1688.790 2774.620 1689.110 ;
        RECT 2774.420 16.730 2774.560 1688.790 ;
        RECT 2774.420 16.590 2780.080 16.730 ;
        RECT 2779.940 2.400 2780.080 16.590 ;
        RECT 2779.730 -4.800 2780.290 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2588.490 1684.940 2588.810 1685.000 ;
        RECT 2594.010 1684.940 2594.330 1685.000 ;
        RECT 2588.490 1684.800 2594.330 1684.940 ;
        RECT 2588.490 1684.740 2588.810 1684.800 ;
        RECT 2594.010 1684.740 2594.330 1684.800 ;
        RECT 2594.010 20.300 2594.330 20.360 ;
        RECT 2797.790 20.300 2798.110 20.360 ;
        RECT 2594.010 20.160 2798.110 20.300 ;
        RECT 2594.010 20.100 2594.330 20.160 ;
        RECT 2797.790 20.100 2798.110 20.160 ;
      LAYER via ;
        RECT 2588.520 1684.740 2588.780 1685.000 ;
        RECT 2594.040 1684.740 2594.300 1685.000 ;
        RECT 2594.040 20.100 2594.300 20.360 ;
        RECT 2797.820 20.100 2798.080 20.360 ;
      LAYER met2 ;
        RECT 2588.440 1700.000 2588.720 1704.000 ;
        RECT 2588.580 1685.030 2588.720 1700.000 ;
        RECT 2588.520 1684.710 2588.780 1685.030 ;
        RECT 2594.040 1684.710 2594.300 1685.030 ;
        RECT 2594.100 20.390 2594.240 1684.710 ;
        RECT 2594.040 20.070 2594.300 20.390 ;
        RECT 2797.820 20.070 2798.080 20.390 ;
        RECT 2797.880 2.400 2798.020 20.070 ;
        RECT 2797.670 -4.800 2798.230 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2815.730 1688.340 2816.050 1688.400 ;
        RECT 2646.080 1688.200 2816.050 1688.340 ;
        RECT 2646.080 1687.660 2646.220 1688.200 ;
        RECT 2815.730 1688.140 2816.050 1688.200 ;
        RECT 2645.160 1687.520 2646.220 1687.660 ;
        RECT 2597.690 1687.320 2598.010 1687.380 ;
        RECT 2645.160 1687.320 2645.300 1687.520 ;
        RECT 2597.690 1687.180 2645.300 1687.320 ;
        RECT 2597.690 1687.120 2598.010 1687.180 ;
      LAYER via ;
        RECT 2815.760 1688.140 2816.020 1688.400 ;
        RECT 2597.720 1687.120 2597.980 1687.380 ;
      LAYER met2 ;
        RECT 2597.640 1700.000 2597.920 1704.000 ;
        RECT 2597.780 1687.410 2597.920 1700.000 ;
        RECT 2815.760 1688.110 2816.020 1688.430 ;
        RECT 2597.720 1687.090 2597.980 1687.410 ;
        RECT 2815.820 2.400 2815.960 1688.110 ;
        RECT 2815.610 -4.800 2816.170 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2607.810 19.280 2608.130 19.340 ;
        RECT 2833.670 19.280 2833.990 19.340 ;
        RECT 2607.810 19.140 2833.990 19.280 ;
        RECT 2607.810 19.080 2608.130 19.140 ;
        RECT 2833.670 19.080 2833.990 19.140 ;
      LAYER via ;
        RECT 2607.840 19.080 2608.100 19.340 ;
        RECT 2833.700 19.080 2833.960 19.340 ;
      LAYER met2 ;
        RECT 2606.840 1700.410 2607.120 1704.000 ;
        RECT 2606.840 1700.270 2608.040 1700.410 ;
        RECT 2606.840 1700.000 2607.120 1700.270 ;
        RECT 2607.900 19.370 2608.040 1700.270 ;
        RECT 2607.840 19.050 2608.100 19.370 ;
        RECT 2833.700 19.050 2833.960 19.370 ;
        RECT 2833.760 2.400 2833.900 19.050 ;
        RECT 2833.550 -4.800 2834.110 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2647.370 1687.320 2647.690 1687.380 ;
        RECT 2846.090 1687.320 2846.410 1687.380 ;
        RECT 2647.370 1687.180 2846.410 1687.320 ;
        RECT 2647.370 1687.120 2647.690 1687.180 ;
        RECT 2846.090 1687.120 2846.410 1687.180 ;
        RECT 2846.090 17.580 2846.410 17.640 ;
        RECT 2851.150 17.580 2851.470 17.640 ;
        RECT 2846.090 17.440 2851.470 17.580 ;
        RECT 2846.090 17.380 2846.410 17.440 ;
        RECT 2851.150 17.380 2851.470 17.440 ;
      LAYER via ;
        RECT 2647.400 1687.120 2647.660 1687.380 ;
        RECT 2846.120 1687.120 2846.380 1687.380 ;
        RECT 2846.120 17.380 2846.380 17.640 ;
        RECT 2851.180 17.380 2851.440 17.640 ;
      LAYER met2 ;
        RECT 2616.040 1700.000 2616.320 1704.000 ;
        RECT 2616.180 1688.965 2616.320 1700.000 ;
        RECT 2616.110 1688.595 2616.390 1688.965 ;
        RECT 2647.390 1688.595 2647.670 1688.965 ;
        RECT 2647.460 1687.410 2647.600 1688.595 ;
        RECT 2647.400 1687.090 2647.660 1687.410 ;
        RECT 2846.120 1687.090 2846.380 1687.410 ;
        RECT 2846.180 17.670 2846.320 1687.090 ;
        RECT 2846.120 17.350 2846.380 17.670 ;
        RECT 2851.180 17.350 2851.440 17.670 ;
        RECT 2851.240 2.400 2851.380 17.350 ;
        RECT 2851.030 -4.800 2851.590 2.400 ;
      LAYER via2 ;
        RECT 2616.110 1688.640 2616.390 1688.920 ;
        RECT 2647.390 1688.640 2647.670 1688.920 ;
      LAYER met3 ;
        RECT 2616.085 1688.930 2616.415 1688.945 ;
        RECT 2647.365 1688.930 2647.695 1688.945 ;
        RECT 2616.085 1688.630 2647.695 1688.930 ;
        RECT 2616.085 1688.615 2616.415 1688.630 ;
        RECT 2647.365 1688.615 2647.695 1688.630 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2627.590 17.920 2627.910 17.980 ;
        RECT 2627.590 17.780 2852.760 17.920 ;
        RECT 2627.590 17.720 2627.910 17.780 ;
        RECT 2852.620 17.580 2852.760 17.780 ;
        RECT 2869.090 17.580 2869.410 17.640 ;
        RECT 2852.620 17.440 2869.410 17.580 ;
        RECT 2869.090 17.380 2869.410 17.440 ;
      LAYER via ;
        RECT 2627.620 17.720 2627.880 17.980 ;
        RECT 2869.120 17.380 2869.380 17.640 ;
      LAYER met2 ;
        RECT 2625.240 1700.410 2625.520 1704.000 ;
        RECT 2625.240 1700.270 2627.820 1700.410 ;
        RECT 2625.240 1700.000 2625.520 1700.270 ;
        RECT 2627.680 18.010 2627.820 1700.270 ;
        RECT 2627.620 17.690 2627.880 18.010 ;
        RECT 2869.120 17.350 2869.380 17.670 ;
        RECT 2869.180 2.400 2869.320 17.350 ;
        RECT 2868.970 -4.800 2869.530 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2645.145 1688.185 2647.155 1688.355 ;
        RECT 2646.985 1686.145 2647.155 1688.185 ;
        RECT 2657.105 1686.145 2657.275 1686.995 ;
      LAYER mcon ;
        RECT 2657.105 1686.825 2657.275 1686.995 ;
      LAYER met1 ;
        RECT 2634.490 1688.340 2634.810 1688.400 ;
        RECT 2645.085 1688.340 2645.375 1688.385 ;
        RECT 2634.490 1688.200 2645.375 1688.340 ;
        RECT 2634.490 1688.140 2634.810 1688.200 ;
        RECT 2645.085 1688.155 2645.375 1688.200 ;
        RECT 2657.045 1686.980 2657.335 1687.025 ;
        RECT 2859.890 1686.980 2860.210 1687.040 ;
        RECT 2657.045 1686.840 2860.210 1686.980 ;
        RECT 2657.045 1686.795 2657.335 1686.840 ;
        RECT 2859.890 1686.780 2860.210 1686.840 ;
        RECT 2646.925 1686.300 2647.215 1686.345 ;
        RECT 2657.045 1686.300 2657.335 1686.345 ;
        RECT 2646.925 1686.160 2657.335 1686.300 ;
        RECT 2646.925 1686.115 2647.215 1686.160 ;
        RECT 2657.045 1686.115 2657.335 1686.160 ;
        RECT 2859.890 15.200 2860.210 15.260 ;
        RECT 2887.030 15.200 2887.350 15.260 ;
        RECT 2859.890 15.060 2887.350 15.200 ;
        RECT 2859.890 15.000 2860.210 15.060 ;
        RECT 2887.030 15.000 2887.350 15.060 ;
      LAYER via ;
        RECT 2634.520 1688.140 2634.780 1688.400 ;
        RECT 2859.920 1686.780 2860.180 1687.040 ;
        RECT 2859.920 15.000 2860.180 15.260 ;
        RECT 2887.060 15.000 2887.320 15.260 ;
      LAYER met2 ;
        RECT 2634.440 1700.000 2634.720 1704.000 ;
        RECT 2634.580 1688.430 2634.720 1700.000 ;
        RECT 2634.520 1688.110 2634.780 1688.430 ;
        RECT 2859.920 1686.750 2860.180 1687.070 ;
        RECT 2859.980 15.290 2860.120 1686.750 ;
        RECT 2859.920 14.970 2860.180 15.290 ;
        RECT 2887.060 14.970 2887.320 15.290 ;
        RECT 2887.120 2.400 2887.260 14.970 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2643.690 1683.920 2644.010 1683.980 ;
        RECT 2649.210 1683.920 2649.530 1683.980 ;
        RECT 2643.690 1683.780 2649.530 1683.920 ;
        RECT 2643.690 1683.720 2644.010 1683.780 ;
        RECT 2649.210 1683.720 2649.530 1683.780 ;
        RECT 2649.210 17.240 2649.530 17.300 ;
        RECT 2904.970 17.240 2905.290 17.300 ;
        RECT 2649.210 17.100 2905.290 17.240 ;
        RECT 2649.210 17.040 2649.530 17.100 ;
        RECT 2904.970 17.040 2905.290 17.100 ;
      LAYER via ;
        RECT 2643.720 1683.720 2643.980 1683.980 ;
        RECT 2649.240 1683.720 2649.500 1683.980 ;
        RECT 2649.240 17.040 2649.500 17.300 ;
        RECT 2905.000 17.040 2905.260 17.300 ;
      LAYER met2 ;
        RECT 2643.640 1700.000 2643.920 1704.000 ;
        RECT 2643.780 1684.010 2643.920 1700.000 ;
        RECT 2643.720 1683.690 2643.980 1684.010 ;
        RECT 2649.240 1683.690 2649.500 1684.010 ;
        RECT 2649.300 17.330 2649.440 1683.690 ;
        RECT 2649.240 17.010 2649.500 17.330 ;
        RECT 2905.000 17.010 2905.260 17.330 ;
        RECT 2905.060 2.400 2905.200 17.010 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 852.910 30.160 853.230 30.220 ;
        RECT 1587.070 30.160 1587.390 30.220 ;
        RECT 852.910 30.020 1587.390 30.160 ;
        RECT 852.910 29.960 853.230 30.020 ;
        RECT 1587.070 29.960 1587.390 30.020 ;
      LAYER via ;
        RECT 852.940 29.960 853.200 30.220 ;
        RECT 1587.100 29.960 1587.360 30.220 ;
      LAYER met2 ;
        RECT 1587.480 1700.410 1587.760 1704.000 ;
        RECT 1587.160 1700.270 1587.760 1700.410 ;
        RECT 1587.160 30.250 1587.300 1700.270 ;
        RECT 1587.480 1700.000 1587.760 1700.270 ;
        RECT 852.940 29.930 853.200 30.250 ;
        RECT 1587.100 29.930 1587.360 30.250 ;
        RECT 853.000 2.400 853.140 29.930 ;
        RECT 852.790 -4.800 853.350 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 870.850 29.820 871.170 29.880 ;
        RECT 870.850 29.680 1576.720 29.820 ;
        RECT 870.850 29.620 871.170 29.680 ;
        RECT 1576.580 29.480 1576.720 29.680 ;
        RECT 1594.430 29.480 1594.750 29.540 ;
        RECT 1576.580 29.340 1594.750 29.480 ;
        RECT 1594.430 29.280 1594.750 29.340 ;
      LAYER via ;
        RECT 870.880 29.620 871.140 29.880 ;
        RECT 1594.460 29.280 1594.720 29.540 ;
      LAYER met2 ;
        RECT 1596.680 1700.410 1596.960 1704.000 ;
        RECT 1594.060 1700.270 1596.960 1700.410 ;
        RECT 1594.060 34.410 1594.200 1700.270 ;
        RECT 1596.680 1700.000 1596.960 1700.270 ;
        RECT 1594.060 34.270 1594.660 34.410 ;
        RECT 870.880 29.590 871.140 29.910 ;
        RECT 870.940 2.400 871.080 29.590 ;
        RECT 1594.520 29.570 1594.660 34.270 ;
        RECT 1594.460 29.250 1594.720 29.570 ;
        RECT 870.730 -4.800 871.290 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1576.105 29.325 1576.275 33.915 ;
      LAYER mcon ;
        RECT 1576.105 33.745 1576.275 33.915 ;
      LAYER met1 ;
        RECT 1600.870 1689.700 1601.190 1689.760 ;
        RECT 1604.550 1689.700 1604.870 1689.760 ;
        RECT 1600.870 1689.560 1604.870 1689.700 ;
        RECT 1600.870 1689.500 1601.190 1689.560 ;
        RECT 1604.550 1689.500 1604.870 1689.560 ;
        RECT 1576.045 33.900 1576.335 33.945 ;
        RECT 1600.870 33.900 1601.190 33.960 ;
        RECT 1576.045 33.760 1601.190 33.900 ;
        RECT 1576.045 33.715 1576.335 33.760 ;
        RECT 1600.870 33.700 1601.190 33.760 ;
        RECT 888.790 29.480 889.110 29.540 ;
        RECT 1576.045 29.480 1576.335 29.525 ;
        RECT 888.790 29.340 1576.335 29.480 ;
        RECT 888.790 29.280 889.110 29.340 ;
        RECT 1576.045 29.295 1576.335 29.340 ;
      LAYER via ;
        RECT 1600.900 1689.500 1601.160 1689.760 ;
        RECT 1604.580 1689.500 1604.840 1689.760 ;
        RECT 1600.900 33.700 1601.160 33.960 ;
        RECT 888.820 29.280 889.080 29.540 ;
      LAYER met2 ;
        RECT 1605.880 1700.410 1606.160 1704.000 ;
        RECT 1604.640 1700.270 1606.160 1700.410 ;
        RECT 1604.640 1689.790 1604.780 1700.270 ;
        RECT 1605.880 1700.000 1606.160 1700.270 ;
        RECT 1600.900 1689.470 1601.160 1689.790 ;
        RECT 1604.580 1689.470 1604.840 1689.790 ;
        RECT 1600.960 33.990 1601.100 1689.470 ;
        RECT 1600.900 33.670 1601.160 33.990 ;
        RECT 888.820 29.250 889.080 29.570 ;
        RECT 888.880 2.400 889.020 29.250 ;
        RECT 888.670 -4.800 889.230 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1611.065 28.985 1611.235 30.175 ;
      LAYER mcon ;
        RECT 1611.065 30.005 1611.235 30.175 ;
      LAYER met1 ;
        RECT 1611.005 30.160 1611.295 30.205 ;
        RECT 1614.670 30.160 1614.990 30.220 ;
        RECT 1611.005 30.020 1614.990 30.160 ;
        RECT 1611.005 29.975 1611.295 30.020 ;
        RECT 1614.670 29.960 1614.990 30.020 ;
        RECT 906.730 29.140 907.050 29.200 ;
        RECT 1611.005 29.140 1611.295 29.185 ;
        RECT 906.730 29.000 1611.295 29.140 ;
        RECT 906.730 28.940 907.050 29.000 ;
        RECT 1611.005 28.955 1611.295 29.000 ;
      LAYER via ;
        RECT 1614.700 29.960 1614.960 30.220 ;
        RECT 906.760 28.940 907.020 29.200 ;
      LAYER met2 ;
        RECT 1615.080 1700.410 1615.360 1704.000 ;
        RECT 1614.760 1700.270 1615.360 1700.410 ;
        RECT 1614.760 30.250 1614.900 1700.270 ;
        RECT 1615.080 1700.000 1615.360 1700.270 ;
        RECT 1614.700 29.930 1614.960 30.250 ;
        RECT 906.760 28.910 907.020 29.230 ;
        RECT 906.820 2.400 906.960 28.910 ;
        RECT 906.610 -4.800 907.170 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 924.210 28.800 924.530 28.860 ;
        RECT 1621.570 28.800 1621.890 28.860 ;
        RECT 924.210 28.660 1621.890 28.800 ;
        RECT 924.210 28.600 924.530 28.660 ;
        RECT 1621.570 28.600 1621.890 28.660 ;
      LAYER via ;
        RECT 924.240 28.600 924.500 28.860 ;
        RECT 1621.600 28.600 1621.860 28.860 ;
      LAYER met2 ;
        RECT 1624.280 1700.410 1624.560 1704.000 ;
        RECT 1621.660 1700.270 1624.560 1700.410 ;
        RECT 1621.660 28.890 1621.800 1700.270 ;
        RECT 1624.280 1700.000 1624.560 1700.270 ;
        RECT 924.240 28.570 924.500 28.890 ;
        RECT 1621.600 28.570 1621.860 28.890 ;
        RECT 924.300 2.400 924.440 28.570 ;
        RECT 924.090 -4.800 924.650 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1628.470 1678.140 1628.790 1678.200 ;
        RECT 1632.150 1678.140 1632.470 1678.200 ;
        RECT 1628.470 1678.000 1632.470 1678.140 ;
        RECT 1628.470 1677.940 1628.790 1678.000 ;
        RECT 1632.150 1677.940 1632.470 1678.000 ;
        RECT 942.150 28.460 942.470 28.520 ;
        RECT 1628.470 28.460 1628.790 28.520 ;
        RECT 942.150 28.320 1628.790 28.460 ;
        RECT 942.150 28.260 942.470 28.320 ;
        RECT 1628.470 28.260 1628.790 28.320 ;
      LAYER via ;
        RECT 1628.500 1677.940 1628.760 1678.200 ;
        RECT 1632.180 1677.940 1632.440 1678.200 ;
        RECT 942.180 28.260 942.440 28.520 ;
        RECT 1628.500 28.260 1628.760 28.520 ;
      LAYER met2 ;
        RECT 1633.480 1700.410 1633.760 1704.000 ;
        RECT 1632.240 1700.270 1633.760 1700.410 ;
        RECT 1632.240 1678.230 1632.380 1700.270 ;
        RECT 1633.480 1700.000 1633.760 1700.270 ;
        RECT 1628.500 1677.910 1628.760 1678.230 ;
        RECT 1632.180 1677.910 1632.440 1678.230 ;
        RECT 1628.560 28.550 1628.700 1677.910 ;
        RECT 942.180 28.230 942.440 28.550 ;
        RECT 1628.500 28.230 1628.760 28.550 ;
        RECT 942.240 2.400 942.380 28.230 ;
        RECT 942.030 -4.800 942.590 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 960.090 28.120 960.410 28.180 ;
        RECT 1642.270 28.120 1642.590 28.180 ;
        RECT 960.090 27.980 1642.590 28.120 ;
        RECT 960.090 27.920 960.410 27.980 ;
        RECT 1642.270 27.920 1642.590 27.980 ;
      LAYER via ;
        RECT 960.120 27.920 960.380 28.180 ;
        RECT 1642.300 27.920 1642.560 28.180 ;
      LAYER met2 ;
        RECT 1642.680 1700.410 1642.960 1704.000 ;
        RECT 1642.360 1700.270 1642.960 1700.410 ;
        RECT 1642.360 28.210 1642.500 1700.270 ;
        RECT 1642.680 1700.000 1642.960 1700.270 ;
        RECT 960.120 27.890 960.380 28.210 ;
        RECT 1642.300 27.890 1642.560 28.210 ;
        RECT 960.180 2.400 960.320 27.890 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 978.030 27.780 978.350 27.840 ;
        RECT 1649.170 27.780 1649.490 27.840 ;
        RECT 978.030 27.640 1649.490 27.780 ;
        RECT 978.030 27.580 978.350 27.640 ;
        RECT 1649.170 27.580 1649.490 27.640 ;
      LAYER via ;
        RECT 978.060 27.580 978.320 27.840 ;
        RECT 1649.200 27.580 1649.460 27.840 ;
      LAYER met2 ;
        RECT 1651.880 1700.410 1652.160 1704.000 ;
        RECT 1649.260 1700.270 1652.160 1700.410 ;
        RECT 1649.260 27.870 1649.400 1700.270 ;
        RECT 1651.880 1700.000 1652.160 1700.270 ;
        RECT 978.060 27.550 978.320 27.870 ;
        RECT 1649.200 27.550 1649.460 27.870 ;
        RECT 978.120 2.400 978.260 27.550 ;
        RECT 977.910 -4.800 978.470 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 662.010 65.860 662.330 65.920 ;
        RECT 1484.490 65.860 1484.810 65.920 ;
        RECT 662.010 65.720 1484.810 65.860 ;
        RECT 662.010 65.660 662.330 65.720 ;
        RECT 1484.490 65.660 1484.810 65.720 ;
      LAYER via ;
        RECT 662.040 65.660 662.300 65.920 ;
        RECT 1484.520 65.660 1484.780 65.920 ;
      LAYER met2 ;
        RECT 1486.740 1700.410 1487.020 1704.000 ;
        RECT 1484.580 1700.270 1487.020 1700.410 ;
        RECT 1484.580 65.950 1484.720 1700.270 ;
        RECT 1486.740 1700.000 1487.020 1700.270 ;
        RECT 662.040 65.630 662.300 65.950 ;
        RECT 1484.520 65.630 1484.780 65.950 ;
        RECT 662.100 17.410 662.240 65.630 ;
        RECT 657.040 17.270 662.240 17.410 ;
        RECT 657.040 2.400 657.180 17.270 ;
        RECT 656.830 -4.800 657.390 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1656.605 1138.745 1656.775 1159.315 ;
        RECT 1657.065 737.205 1657.235 772.735 ;
        RECT 1657.065 241.485 1657.235 324.275 ;
      LAYER mcon ;
        RECT 1656.605 1159.145 1656.775 1159.315 ;
        RECT 1657.065 772.565 1657.235 772.735 ;
        RECT 1657.065 324.105 1657.235 324.275 ;
      LAYER met1 ;
        RECT 1657.450 1642.440 1657.770 1642.500 ;
        RECT 1658.370 1642.440 1658.690 1642.500 ;
        RECT 1657.450 1642.300 1658.690 1642.440 ;
        RECT 1657.450 1642.240 1657.770 1642.300 ;
        RECT 1658.370 1642.240 1658.690 1642.300 ;
        RECT 1656.990 1497.260 1657.310 1497.320 ;
        RECT 1657.450 1497.260 1657.770 1497.320 ;
        RECT 1656.990 1497.120 1657.770 1497.260 ;
        RECT 1656.990 1497.060 1657.310 1497.120 ;
        RECT 1657.450 1497.060 1657.770 1497.120 ;
        RECT 1656.990 1400.700 1657.310 1400.760 ;
        RECT 1657.450 1400.700 1657.770 1400.760 ;
        RECT 1656.990 1400.560 1657.770 1400.700 ;
        RECT 1656.990 1400.500 1657.310 1400.560 ;
        RECT 1657.450 1400.500 1657.770 1400.560 ;
        RECT 1656.530 1317.740 1656.850 1317.800 ;
        RECT 1656.530 1317.600 1657.680 1317.740 ;
        RECT 1656.530 1317.540 1656.850 1317.600 ;
        RECT 1657.540 1317.460 1657.680 1317.600 ;
        RECT 1657.450 1317.200 1657.770 1317.460 ;
        RECT 1655.610 1304.140 1655.930 1304.200 ;
        RECT 1657.450 1304.140 1657.770 1304.200 ;
        RECT 1655.610 1304.000 1657.770 1304.140 ;
        RECT 1655.610 1303.940 1655.930 1304.000 ;
        RECT 1657.450 1303.940 1657.770 1304.000 ;
        RECT 1655.610 1207.580 1655.930 1207.640 ;
        RECT 1657.450 1207.580 1657.770 1207.640 ;
        RECT 1655.610 1207.440 1657.770 1207.580 ;
        RECT 1655.610 1207.380 1655.930 1207.440 ;
        RECT 1657.450 1207.380 1657.770 1207.440 ;
        RECT 1656.545 1159.300 1656.835 1159.345 ;
        RECT 1657.450 1159.300 1657.770 1159.360 ;
        RECT 1656.545 1159.160 1657.770 1159.300 ;
        RECT 1656.545 1159.115 1656.835 1159.160 ;
        RECT 1657.450 1159.100 1657.770 1159.160 ;
        RECT 1656.530 1138.900 1656.850 1138.960 ;
        RECT 1656.335 1138.760 1656.850 1138.900 ;
        RECT 1656.530 1138.700 1656.850 1138.760 ;
        RECT 1655.610 1048.800 1655.930 1048.860 ;
        RECT 1656.530 1048.800 1656.850 1048.860 ;
        RECT 1655.610 1048.660 1656.850 1048.800 ;
        RECT 1655.610 1048.600 1655.930 1048.660 ;
        RECT 1656.530 1048.600 1656.850 1048.660 ;
        RECT 1656.990 917.900 1657.310 917.960 ;
        RECT 1657.450 917.900 1657.770 917.960 ;
        RECT 1656.990 917.760 1657.770 917.900 ;
        RECT 1656.990 917.700 1657.310 917.760 ;
        RECT 1657.450 917.700 1657.770 917.760 ;
        RECT 1657.450 910.760 1657.770 910.820 ;
        RECT 1657.910 910.760 1658.230 910.820 ;
        RECT 1657.450 910.620 1658.230 910.760 ;
        RECT 1657.450 910.560 1657.770 910.620 ;
        RECT 1657.910 910.560 1658.230 910.620 ;
        RECT 1656.990 772.720 1657.310 772.780 ;
        RECT 1656.795 772.580 1657.310 772.720 ;
        RECT 1656.990 772.520 1657.310 772.580 ;
        RECT 1657.005 737.360 1657.295 737.405 ;
        RECT 1657.450 737.360 1657.770 737.420 ;
        RECT 1657.005 737.220 1657.770 737.360 ;
        RECT 1657.005 737.175 1657.295 737.220 ;
        RECT 1657.450 737.160 1657.770 737.220 ;
        RECT 1656.530 435.100 1656.850 435.160 ;
        RECT 1656.990 435.100 1657.310 435.160 ;
        RECT 1656.530 434.960 1657.310 435.100 ;
        RECT 1656.530 434.900 1656.850 434.960 ;
        RECT 1656.990 434.900 1657.310 434.960 ;
        RECT 1656.990 338.680 1657.310 338.940 ;
        RECT 1657.080 338.260 1657.220 338.680 ;
        RECT 1656.990 338.000 1657.310 338.260 ;
        RECT 1656.990 324.260 1657.310 324.320 ;
        RECT 1656.795 324.120 1657.310 324.260 ;
        RECT 1656.990 324.060 1657.310 324.120 ;
        RECT 1657.005 241.640 1657.295 241.685 ;
        RECT 1657.450 241.640 1657.770 241.700 ;
        RECT 1657.005 241.500 1657.770 241.640 ;
        RECT 1657.005 241.455 1657.295 241.500 ;
        RECT 1657.450 241.440 1657.770 241.500 ;
        RECT 1656.990 186.560 1657.310 186.620 ;
        RECT 1657.450 186.560 1657.770 186.620 ;
        RECT 1656.990 186.420 1657.770 186.560 ;
        RECT 1656.990 186.360 1657.310 186.420 ;
        RECT 1657.450 186.360 1657.770 186.420 ;
        RECT 1656.530 137.940 1656.850 138.000 ;
        RECT 1656.990 137.940 1657.310 138.000 ;
        RECT 1656.530 137.800 1657.310 137.940 ;
        RECT 1656.530 137.740 1656.850 137.800 ;
        RECT 1656.990 137.740 1657.310 137.800 ;
        RECT 1000.110 65.180 1000.430 65.240 ;
        RECT 1656.530 65.180 1656.850 65.240 ;
        RECT 1000.110 65.040 1656.850 65.180 ;
        RECT 1000.110 64.980 1000.430 65.040 ;
        RECT 1656.530 64.980 1656.850 65.040 ;
      LAYER via ;
        RECT 1657.480 1642.240 1657.740 1642.500 ;
        RECT 1658.400 1642.240 1658.660 1642.500 ;
        RECT 1657.020 1497.060 1657.280 1497.320 ;
        RECT 1657.480 1497.060 1657.740 1497.320 ;
        RECT 1657.020 1400.500 1657.280 1400.760 ;
        RECT 1657.480 1400.500 1657.740 1400.760 ;
        RECT 1656.560 1317.540 1656.820 1317.800 ;
        RECT 1657.480 1317.200 1657.740 1317.460 ;
        RECT 1655.640 1303.940 1655.900 1304.200 ;
        RECT 1657.480 1303.940 1657.740 1304.200 ;
        RECT 1655.640 1207.380 1655.900 1207.640 ;
        RECT 1657.480 1207.380 1657.740 1207.640 ;
        RECT 1657.480 1159.100 1657.740 1159.360 ;
        RECT 1656.560 1138.700 1656.820 1138.960 ;
        RECT 1655.640 1048.600 1655.900 1048.860 ;
        RECT 1656.560 1048.600 1656.820 1048.860 ;
        RECT 1657.020 917.700 1657.280 917.960 ;
        RECT 1657.480 917.700 1657.740 917.960 ;
        RECT 1657.480 910.560 1657.740 910.820 ;
        RECT 1657.940 910.560 1658.200 910.820 ;
        RECT 1657.020 772.520 1657.280 772.780 ;
        RECT 1657.480 737.160 1657.740 737.420 ;
        RECT 1656.560 434.900 1656.820 435.160 ;
        RECT 1657.020 434.900 1657.280 435.160 ;
        RECT 1657.020 338.680 1657.280 338.940 ;
        RECT 1657.020 338.000 1657.280 338.260 ;
        RECT 1657.020 324.060 1657.280 324.320 ;
        RECT 1657.480 241.440 1657.740 241.700 ;
        RECT 1657.020 186.360 1657.280 186.620 ;
        RECT 1657.480 186.360 1657.740 186.620 ;
        RECT 1656.560 137.740 1656.820 138.000 ;
        RECT 1657.020 137.740 1657.280 138.000 ;
        RECT 1000.140 64.980 1000.400 65.240 ;
        RECT 1656.560 64.980 1656.820 65.240 ;
      LAYER met2 ;
        RECT 1661.080 1701.090 1661.360 1704.000 ;
        RECT 1658.460 1700.950 1661.360 1701.090 ;
        RECT 1658.460 1642.530 1658.600 1700.950 ;
        RECT 1661.080 1700.000 1661.360 1700.950 ;
        RECT 1657.480 1642.210 1657.740 1642.530 ;
        RECT 1658.400 1642.210 1658.660 1642.530 ;
        RECT 1657.540 1546.050 1657.680 1642.210 ;
        RECT 1657.080 1545.910 1657.680 1546.050 ;
        RECT 1657.080 1521.570 1657.220 1545.910 ;
        RECT 1656.620 1521.430 1657.220 1521.570 ;
        RECT 1656.620 1510.010 1656.760 1521.430 ;
        RECT 1656.620 1509.870 1657.680 1510.010 ;
        RECT 1657.540 1497.350 1657.680 1509.870 ;
        RECT 1657.020 1497.030 1657.280 1497.350 ;
        RECT 1657.480 1497.030 1657.740 1497.350 ;
        RECT 1657.080 1450.285 1657.220 1497.030 ;
        RECT 1657.010 1449.915 1657.290 1450.285 ;
        RECT 1656.550 1448.555 1656.830 1448.925 ;
        RECT 1656.620 1414.130 1656.760 1448.555 ;
        RECT 1656.620 1413.990 1657.680 1414.130 ;
        RECT 1657.540 1400.790 1657.680 1413.990 ;
        RECT 1657.020 1400.470 1657.280 1400.790 ;
        RECT 1657.480 1400.470 1657.740 1400.790 ;
        RECT 1657.080 1353.725 1657.220 1400.470 ;
        RECT 1657.010 1353.355 1657.290 1353.725 ;
        RECT 1656.550 1351.995 1656.830 1352.365 ;
        RECT 1656.620 1317.830 1656.760 1351.995 ;
        RECT 1656.560 1317.510 1656.820 1317.830 ;
        RECT 1657.480 1317.170 1657.740 1317.490 ;
        RECT 1657.540 1304.230 1657.680 1317.170 ;
        RECT 1655.640 1303.910 1655.900 1304.230 ;
        RECT 1657.480 1303.910 1657.740 1304.230 ;
        RECT 1655.700 1256.485 1655.840 1303.910 ;
        RECT 1655.630 1256.115 1655.910 1256.485 ;
        RECT 1655.630 1255.435 1655.910 1255.805 ;
        RECT 1655.700 1207.670 1655.840 1255.435 ;
        RECT 1655.640 1207.350 1655.900 1207.670 ;
        RECT 1657.480 1207.350 1657.740 1207.670 ;
        RECT 1657.540 1159.390 1657.680 1207.350 ;
        RECT 1657.480 1159.070 1657.740 1159.390 ;
        RECT 1656.560 1138.670 1656.820 1138.990 ;
        RECT 1656.620 1048.890 1656.760 1138.670 ;
        RECT 1655.640 1048.570 1655.900 1048.890 ;
        RECT 1656.560 1048.570 1656.820 1048.890 ;
        RECT 1655.700 1000.805 1655.840 1048.570 ;
        RECT 1655.630 1000.435 1655.910 1000.805 ;
        RECT 1657.010 1000.435 1657.290 1000.805 ;
        RECT 1657.080 917.990 1657.220 1000.435 ;
        RECT 1657.020 917.670 1657.280 917.990 ;
        RECT 1657.480 917.670 1657.740 917.990 ;
        RECT 1657.540 910.850 1657.680 917.670 ;
        RECT 1657.480 910.530 1657.740 910.850 ;
        RECT 1657.940 910.530 1658.200 910.850 ;
        RECT 1658.000 773.005 1658.140 910.530 ;
        RECT 1657.010 772.635 1657.290 773.005 ;
        RECT 1657.930 772.635 1658.210 773.005 ;
        RECT 1657.020 772.490 1657.280 772.635 ;
        RECT 1657.480 737.130 1657.740 737.450 ;
        RECT 1657.540 669.530 1657.680 737.130 ;
        RECT 1657.080 669.390 1657.680 669.530 ;
        RECT 1657.080 640.970 1657.220 669.390 ;
        RECT 1657.080 640.830 1657.680 640.970 ;
        RECT 1657.540 596.770 1657.680 640.830 ;
        RECT 1657.540 596.630 1658.140 596.770 ;
        RECT 1658.000 554.610 1658.140 596.630 ;
        RECT 1657.540 554.470 1658.140 554.610 ;
        RECT 1657.540 498.170 1657.680 554.470 ;
        RECT 1657.080 498.030 1657.680 498.170 ;
        RECT 1657.080 483.210 1657.220 498.030 ;
        RECT 1657.080 483.070 1657.680 483.210 ;
        RECT 1657.540 482.530 1657.680 483.070 ;
        RECT 1656.620 482.390 1657.680 482.530 ;
        RECT 1656.620 435.190 1656.760 482.390 ;
        RECT 1656.560 434.870 1656.820 435.190 ;
        RECT 1657.020 434.870 1657.280 435.190 ;
        RECT 1657.080 338.970 1657.220 434.870 ;
        RECT 1657.020 338.650 1657.280 338.970 ;
        RECT 1657.020 337.970 1657.280 338.290 ;
        RECT 1657.080 324.350 1657.220 337.970 ;
        RECT 1657.020 324.030 1657.280 324.350 ;
        RECT 1657.480 241.410 1657.740 241.730 ;
        RECT 1657.540 186.650 1657.680 241.410 ;
        RECT 1657.020 186.330 1657.280 186.650 ;
        RECT 1657.480 186.330 1657.740 186.650 ;
        RECT 1657.080 138.030 1657.220 186.330 ;
        RECT 1656.560 137.710 1656.820 138.030 ;
        RECT 1657.020 137.710 1657.280 138.030 ;
        RECT 1656.620 65.270 1656.760 137.710 ;
        RECT 1000.140 64.950 1000.400 65.270 ;
        RECT 1656.560 64.950 1656.820 65.270 ;
        RECT 1000.200 17.410 1000.340 64.950 ;
        RECT 996.060 17.270 1000.340 17.410 ;
        RECT 996.060 2.400 996.200 17.270 ;
        RECT 995.850 -4.800 996.410 2.400 ;
      LAYER via2 ;
        RECT 1657.010 1449.960 1657.290 1450.240 ;
        RECT 1656.550 1448.600 1656.830 1448.880 ;
        RECT 1657.010 1353.400 1657.290 1353.680 ;
        RECT 1656.550 1352.040 1656.830 1352.320 ;
        RECT 1655.630 1256.160 1655.910 1256.440 ;
        RECT 1655.630 1255.480 1655.910 1255.760 ;
        RECT 1655.630 1000.480 1655.910 1000.760 ;
        RECT 1657.010 1000.480 1657.290 1000.760 ;
        RECT 1657.010 772.680 1657.290 772.960 ;
        RECT 1657.930 772.680 1658.210 772.960 ;
      LAYER met3 ;
        RECT 1656.985 1450.250 1657.315 1450.265 ;
        RECT 1656.310 1449.950 1657.315 1450.250 ;
        RECT 1656.310 1448.905 1656.610 1449.950 ;
        RECT 1656.985 1449.935 1657.315 1449.950 ;
        RECT 1656.310 1448.590 1656.855 1448.905 ;
        RECT 1656.525 1448.575 1656.855 1448.590 ;
        RECT 1656.985 1353.690 1657.315 1353.705 ;
        RECT 1656.310 1353.390 1657.315 1353.690 ;
        RECT 1656.310 1352.345 1656.610 1353.390 ;
        RECT 1656.985 1353.375 1657.315 1353.390 ;
        RECT 1656.310 1352.030 1656.855 1352.345 ;
        RECT 1656.525 1352.015 1656.855 1352.030 ;
        RECT 1655.605 1256.450 1655.935 1256.465 ;
        RECT 1655.605 1256.150 1656.610 1256.450 ;
        RECT 1655.605 1256.135 1655.935 1256.150 ;
        RECT 1655.605 1255.770 1655.935 1255.785 ;
        RECT 1656.310 1255.770 1656.610 1256.150 ;
        RECT 1655.605 1255.470 1656.610 1255.770 ;
        RECT 1655.605 1255.455 1655.935 1255.470 ;
        RECT 1655.605 1000.770 1655.935 1000.785 ;
        RECT 1656.985 1000.770 1657.315 1000.785 ;
        RECT 1655.605 1000.470 1657.315 1000.770 ;
        RECT 1655.605 1000.455 1655.935 1000.470 ;
        RECT 1656.985 1000.455 1657.315 1000.470 ;
        RECT 1656.985 772.970 1657.315 772.985 ;
        RECT 1657.905 772.970 1658.235 772.985 ;
        RECT 1656.985 772.670 1658.235 772.970 ;
        RECT 1656.985 772.655 1657.315 772.670 ;
        RECT 1657.905 772.655 1658.235 772.670 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1670.330 1677.120 1670.650 1677.180 ;
        RECT 1670.330 1676.980 1671.020 1677.120 ;
        RECT 1670.330 1676.920 1670.650 1676.980 ;
        RECT 1670.880 1676.160 1671.020 1676.980 ;
        RECT 1670.790 1675.900 1671.110 1676.160 ;
        RECT 1013.910 68.920 1014.230 68.980 ;
        RECT 1670.790 68.920 1671.110 68.980 ;
        RECT 1013.910 68.780 1671.110 68.920 ;
        RECT 1013.910 68.720 1014.230 68.780 ;
        RECT 1670.790 68.720 1671.110 68.780 ;
      LAYER via ;
        RECT 1670.360 1676.920 1670.620 1677.180 ;
        RECT 1670.820 1675.900 1671.080 1676.160 ;
        RECT 1013.940 68.720 1014.200 68.980 ;
        RECT 1670.820 68.720 1671.080 68.980 ;
      LAYER met2 ;
        RECT 1670.280 1700.000 1670.560 1704.000 ;
        RECT 1670.420 1677.210 1670.560 1700.000 ;
        RECT 1670.360 1676.890 1670.620 1677.210 ;
        RECT 1670.820 1675.870 1671.080 1676.190 ;
        RECT 1670.880 69.010 1671.020 1675.870 ;
        RECT 1013.940 68.690 1014.200 69.010 ;
        RECT 1670.820 68.690 1671.080 69.010 ;
        RECT 1014.000 17.410 1014.140 68.690 ;
        RECT 1013.540 17.270 1014.140 17.410 ;
        RECT 1013.540 2.400 1013.680 17.270 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1034.610 64.840 1034.930 64.900 ;
        RECT 1677.230 64.840 1677.550 64.900 ;
        RECT 1034.610 64.700 1677.550 64.840 ;
        RECT 1034.610 64.640 1034.930 64.700 ;
        RECT 1677.230 64.640 1677.550 64.700 ;
        RECT 1031.390 2.960 1031.710 3.020 ;
        RECT 1034.610 2.960 1034.930 3.020 ;
        RECT 1031.390 2.820 1034.930 2.960 ;
        RECT 1031.390 2.760 1031.710 2.820 ;
        RECT 1034.610 2.760 1034.930 2.820 ;
      LAYER via ;
        RECT 1034.640 64.640 1034.900 64.900 ;
        RECT 1677.260 64.640 1677.520 64.900 ;
        RECT 1031.420 2.760 1031.680 3.020 ;
        RECT 1034.640 2.760 1034.900 3.020 ;
      LAYER met2 ;
        RECT 1679.480 1700.410 1679.760 1704.000 ;
        RECT 1677.320 1700.270 1679.760 1700.410 ;
        RECT 1677.320 64.930 1677.460 1700.270 ;
        RECT 1679.480 1700.000 1679.760 1700.270 ;
        RECT 1034.640 64.610 1034.900 64.930 ;
        RECT 1677.260 64.610 1677.520 64.930 ;
        RECT 1034.700 3.050 1034.840 64.610 ;
        RECT 1031.420 2.730 1031.680 3.050 ;
        RECT 1034.640 2.730 1034.900 3.050 ;
        RECT 1031.480 2.400 1031.620 2.730 ;
        RECT 1031.270 -4.800 1031.830 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1684.205 1014.305 1684.375 1028.415 ;
        RECT 1684.205 882.725 1684.375 910.775 ;
      LAYER mcon ;
        RECT 1684.205 1028.245 1684.375 1028.415 ;
        RECT 1684.205 910.605 1684.375 910.775 ;
      LAYER met1 ;
        RECT 1684.590 1642.440 1684.910 1642.500 ;
        RECT 1685.970 1642.440 1686.290 1642.500 ;
        RECT 1684.590 1642.300 1686.290 1642.440 ;
        RECT 1684.590 1642.240 1684.910 1642.300 ;
        RECT 1685.970 1642.240 1686.290 1642.300 ;
        RECT 1684.130 1545.880 1684.450 1545.940 ;
        RECT 1684.590 1545.880 1684.910 1545.940 ;
        RECT 1684.130 1545.740 1684.910 1545.880 ;
        RECT 1684.130 1545.680 1684.450 1545.740 ;
        RECT 1684.590 1545.680 1684.910 1545.740 ;
        RECT 1684.130 1028.400 1684.450 1028.460 ;
        RECT 1683.935 1028.260 1684.450 1028.400 ;
        RECT 1684.130 1028.200 1684.450 1028.260 ;
        RECT 1684.130 1014.460 1684.450 1014.520 ;
        RECT 1683.935 1014.320 1684.450 1014.460 ;
        RECT 1684.130 1014.260 1684.450 1014.320 ;
        RECT 1683.670 966.180 1683.990 966.240 ;
        RECT 1684.130 966.180 1684.450 966.240 ;
        RECT 1683.670 966.040 1684.450 966.180 ;
        RECT 1683.670 965.980 1683.990 966.040 ;
        RECT 1684.130 965.980 1684.450 966.040 ;
        RECT 1683.670 917.900 1683.990 917.960 ;
        RECT 1684.130 917.900 1684.450 917.960 ;
        RECT 1683.670 917.760 1684.450 917.900 ;
        RECT 1683.670 917.700 1683.990 917.760 ;
        RECT 1684.130 917.700 1684.450 917.760 ;
        RECT 1684.130 910.760 1684.450 910.820 ;
        RECT 1683.935 910.620 1684.450 910.760 ;
        RECT 1684.130 910.560 1684.450 910.620 ;
        RECT 1684.130 882.880 1684.450 882.940 ;
        RECT 1683.935 882.740 1684.450 882.880 ;
        RECT 1684.130 882.680 1684.450 882.740 ;
        RECT 1684.130 593.340 1684.450 593.600 ;
        RECT 1684.220 592.920 1684.360 593.340 ;
        RECT 1684.130 592.660 1684.450 592.920 ;
        RECT 1684.130 400.220 1684.450 400.480 ;
        RECT 1684.220 399.800 1684.360 400.220 ;
        RECT 1684.130 399.540 1684.450 399.800 ;
        RECT 1682.750 76.060 1683.070 76.120 ;
        RECT 1684.130 76.060 1684.450 76.120 ;
        RECT 1682.750 75.920 1684.450 76.060 ;
        RECT 1682.750 75.860 1683.070 75.920 ;
        RECT 1684.130 75.860 1684.450 75.920 ;
        RECT 1055.310 64.160 1055.630 64.220 ;
        RECT 1684.130 64.160 1684.450 64.220 ;
        RECT 1055.310 64.020 1684.450 64.160 ;
        RECT 1055.310 63.960 1055.630 64.020 ;
        RECT 1684.130 63.960 1684.450 64.020 ;
        RECT 1049.330 20.980 1049.650 21.040 ;
        RECT 1055.310 20.980 1055.630 21.040 ;
        RECT 1049.330 20.840 1055.630 20.980 ;
        RECT 1049.330 20.780 1049.650 20.840 ;
        RECT 1055.310 20.780 1055.630 20.840 ;
      LAYER via ;
        RECT 1684.620 1642.240 1684.880 1642.500 ;
        RECT 1686.000 1642.240 1686.260 1642.500 ;
        RECT 1684.160 1545.680 1684.420 1545.940 ;
        RECT 1684.620 1545.680 1684.880 1545.940 ;
        RECT 1684.160 1028.200 1684.420 1028.460 ;
        RECT 1684.160 1014.260 1684.420 1014.520 ;
        RECT 1683.700 965.980 1683.960 966.240 ;
        RECT 1684.160 965.980 1684.420 966.240 ;
        RECT 1683.700 917.700 1683.960 917.960 ;
        RECT 1684.160 917.700 1684.420 917.960 ;
        RECT 1684.160 910.560 1684.420 910.820 ;
        RECT 1684.160 882.680 1684.420 882.940 ;
        RECT 1684.160 593.340 1684.420 593.600 ;
        RECT 1684.160 592.660 1684.420 592.920 ;
        RECT 1684.160 400.220 1684.420 400.480 ;
        RECT 1684.160 399.540 1684.420 399.800 ;
        RECT 1682.780 75.860 1683.040 76.120 ;
        RECT 1684.160 75.860 1684.420 76.120 ;
        RECT 1055.340 63.960 1055.600 64.220 ;
        RECT 1684.160 63.960 1684.420 64.220 ;
        RECT 1049.360 20.780 1049.620 21.040 ;
        RECT 1055.340 20.780 1055.600 21.040 ;
      LAYER met2 ;
        RECT 1688.680 1701.090 1688.960 1704.000 ;
        RECT 1686.060 1700.950 1688.960 1701.090 ;
        RECT 1686.060 1642.530 1686.200 1700.950 ;
        RECT 1688.680 1700.000 1688.960 1700.950 ;
        RECT 1684.620 1642.210 1684.880 1642.530 ;
        RECT 1686.000 1642.210 1686.260 1642.530 ;
        RECT 1684.680 1545.970 1684.820 1642.210 ;
        RECT 1684.160 1545.650 1684.420 1545.970 ;
        RECT 1684.620 1545.650 1684.880 1545.970 ;
        RECT 1684.220 1511.370 1684.360 1545.650 ;
        RECT 1683.760 1511.230 1684.360 1511.370 ;
        RECT 1683.760 1510.690 1683.900 1511.230 ;
        RECT 1683.760 1510.550 1684.360 1510.690 ;
        RECT 1684.220 1414.810 1684.360 1510.550 ;
        RECT 1683.760 1414.670 1684.360 1414.810 ;
        RECT 1683.760 1414.130 1683.900 1414.670 ;
        RECT 1683.760 1413.990 1684.360 1414.130 ;
        RECT 1684.220 1318.250 1684.360 1413.990 ;
        RECT 1683.760 1318.110 1684.360 1318.250 ;
        RECT 1683.760 1317.570 1683.900 1318.110 ;
        RECT 1683.760 1317.430 1684.360 1317.570 ;
        RECT 1684.220 1221.690 1684.360 1317.430 ;
        RECT 1683.760 1221.550 1684.360 1221.690 ;
        RECT 1683.760 1221.010 1683.900 1221.550 ;
        RECT 1683.760 1220.870 1684.360 1221.010 ;
        RECT 1684.220 1125.130 1684.360 1220.870 ;
        RECT 1683.760 1124.990 1684.360 1125.130 ;
        RECT 1683.760 1124.450 1683.900 1124.990 ;
        RECT 1683.760 1124.310 1684.360 1124.450 ;
        RECT 1684.220 1028.490 1684.360 1124.310 ;
        RECT 1684.160 1028.170 1684.420 1028.490 ;
        RECT 1684.160 1014.230 1684.420 1014.550 ;
        RECT 1684.220 966.270 1684.360 1014.230 ;
        RECT 1683.700 965.950 1683.960 966.270 ;
        RECT 1684.160 965.950 1684.420 966.270 ;
        RECT 1683.760 917.990 1683.900 965.950 ;
        RECT 1683.700 917.670 1683.960 917.990 ;
        RECT 1684.160 917.670 1684.420 917.990 ;
        RECT 1684.220 910.850 1684.360 917.670 ;
        RECT 1684.160 910.530 1684.420 910.850 ;
        RECT 1684.160 882.650 1684.420 882.970 ;
        RECT 1684.220 690.610 1684.360 882.650 ;
        RECT 1683.760 690.470 1684.360 690.610 ;
        RECT 1683.760 689.930 1683.900 690.470 ;
        RECT 1683.760 689.790 1684.360 689.930 ;
        RECT 1684.220 593.630 1684.360 689.790 ;
        RECT 1684.160 593.310 1684.420 593.630 ;
        RECT 1684.160 592.630 1684.420 592.950 ;
        RECT 1684.220 400.510 1684.360 592.630 ;
        RECT 1684.160 400.190 1684.420 400.510 ;
        RECT 1684.160 399.510 1684.420 399.830 ;
        RECT 1684.220 303.690 1684.360 399.510 ;
        RECT 1683.760 303.550 1684.360 303.690 ;
        RECT 1683.760 303.010 1683.900 303.550 ;
        RECT 1683.760 302.870 1684.360 303.010 ;
        RECT 1684.220 138.450 1684.360 302.870 ;
        RECT 1683.760 138.310 1684.360 138.450 ;
        RECT 1683.760 124.285 1683.900 138.310 ;
        RECT 1682.770 123.915 1683.050 124.285 ;
        RECT 1683.690 123.915 1683.970 124.285 ;
        RECT 1682.840 76.150 1682.980 123.915 ;
        RECT 1682.780 75.830 1683.040 76.150 ;
        RECT 1684.160 75.830 1684.420 76.150 ;
        RECT 1684.220 64.250 1684.360 75.830 ;
        RECT 1055.340 63.930 1055.600 64.250 ;
        RECT 1684.160 63.930 1684.420 64.250 ;
        RECT 1055.400 21.070 1055.540 63.930 ;
        RECT 1049.360 20.750 1049.620 21.070 ;
        RECT 1055.340 20.750 1055.600 21.070 ;
        RECT 1049.420 2.400 1049.560 20.750 ;
        RECT 1049.210 -4.800 1049.770 2.400 ;
      LAYER via2 ;
        RECT 1682.770 123.960 1683.050 124.240 ;
        RECT 1683.690 123.960 1683.970 124.240 ;
      LAYER met3 ;
        RECT 1682.745 124.250 1683.075 124.265 ;
        RECT 1683.665 124.250 1683.995 124.265 ;
        RECT 1682.745 123.950 1683.995 124.250 ;
        RECT 1682.745 123.935 1683.075 123.950 ;
        RECT 1683.665 123.935 1683.995 123.950 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1069.110 64.500 1069.430 64.560 ;
        RECT 1698.390 64.500 1698.710 64.560 ;
        RECT 1069.110 64.360 1698.710 64.500 ;
        RECT 1069.110 64.300 1069.430 64.360 ;
        RECT 1698.390 64.300 1698.710 64.360 ;
      LAYER via ;
        RECT 1069.140 64.300 1069.400 64.560 ;
        RECT 1698.420 64.300 1698.680 64.560 ;
      LAYER met2 ;
        RECT 1697.880 1700.410 1698.160 1704.000 ;
        RECT 1697.880 1700.270 1698.620 1700.410 ;
        RECT 1697.880 1700.000 1698.160 1700.270 ;
        RECT 1698.480 64.590 1698.620 1700.270 ;
        RECT 1069.140 64.270 1069.400 64.590 ;
        RECT 1698.420 64.270 1698.680 64.590 ;
        RECT 1069.200 17.410 1069.340 64.270 ;
        RECT 1067.360 17.270 1069.340 17.410 ;
        RECT 1067.360 2.400 1067.500 17.270 ;
        RECT 1067.150 -4.800 1067.710 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1089.810 63.820 1090.130 63.880 ;
        RECT 1704.830 63.820 1705.150 63.880 ;
        RECT 1089.810 63.680 1705.150 63.820 ;
        RECT 1089.810 63.620 1090.130 63.680 ;
        RECT 1704.830 63.620 1705.150 63.680 ;
      LAYER via ;
        RECT 1089.840 63.620 1090.100 63.880 ;
        RECT 1704.860 63.620 1705.120 63.880 ;
      LAYER met2 ;
        RECT 1707.080 1700.410 1707.360 1704.000 ;
        RECT 1704.920 1700.270 1707.360 1700.410 ;
        RECT 1704.920 63.910 1705.060 1700.270 ;
        RECT 1707.080 1700.000 1707.360 1700.270 ;
        RECT 1089.840 63.590 1090.100 63.910 ;
        RECT 1704.860 63.590 1705.120 63.910 ;
        RECT 1089.900 17.410 1090.040 63.590 ;
        RECT 1085.300 17.270 1090.040 17.410 ;
        RECT 1085.300 2.400 1085.440 17.270 ;
        RECT 1085.090 -4.800 1085.650 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1712.265 1497.785 1712.435 1545.215 ;
        RECT 1712.725 1401.225 1712.895 1414.655 ;
        RECT 1712.725 1304.325 1712.895 1318.095 ;
        RECT 1712.265 1256.045 1712.435 1303.815 ;
        RECT 1711.805 814.385 1711.975 862.495 ;
        RECT 1713.185 572.645 1713.355 620.755 ;
        RECT 1712.725 399.925 1712.895 434.775 ;
        RECT 1712.265 227.885 1712.435 275.995 ;
        RECT 1711.805 96.645 1711.975 162.095 ;
      LAYER mcon ;
        RECT 1712.265 1545.045 1712.435 1545.215 ;
        RECT 1712.725 1414.485 1712.895 1414.655 ;
        RECT 1712.725 1317.925 1712.895 1318.095 ;
        RECT 1712.265 1303.645 1712.435 1303.815 ;
        RECT 1711.805 862.325 1711.975 862.495 ;
        RECT 1713.185 620.585 1713.355 620.755 ;
        RECT 1712.725 434.605 1712.895 434.775 ;
        RECT 1712.265 275.825 1712.435 275.995 ;
        RECT 1711.805 161.925 1711.975 162.095 ;
      LAYER met1 ;
        RECT 1713.110 1642.440 1713.430 1642.500 ;
        RECT 1714.950 1642.440 1715.270 1642.500 ;
        RECT 1713.110 1642.300 1715.270 1642.440 ;
        RECT 1713.110 1642.240 1713.430 1642.300 ;
        RECT 1714.950 1642.240 1715.270 1642.300 ;
        RECT 1713.110 1546.220 1713.430 1546.280 ;
        RECT 1712.280 1546.080 1713.430 1546.220 ;
        RECT 1712.280 1545.940 1712.420 1546.080 ;
        RECT 1713.110 1546.020 1713.430 1546.080 ;
        RECT 1712.190 1545.680 1712.510 1545.940 ;
        RECT 1712.190 1545.200 1712.510 1545.260 ;
        RECT 1711.995 1545.060 1712.510 1545.200 ;
        RECT 1712.190 1545.000 1712.510 1545.060 ;
        RECT 1712.205 1497.940 1712.495 1497.985 ;
        RECT 1712.650 1497.940 1712.970 1498.000 ;
        RECT 1712.205 1497.800 1712.970 1497.940 ;
        RECT 1712.205 1497.755 1712.495 1497.800 ;
        RECT 1712.650 1497.740 1712.970 1497.800 ;
        RECT 1712.650 1414.640 1712.970 1414.700 ;
        RECT 1712.455 1414.500 1712.970 1414.640 ;
        RECT 1712.650 1414.440 1712.970 1414.500 ;
        RECT 1712.650 1401.380 1712.970 1401.440 ;
        RECT 1712.455 1401.240 1712.970 1401.380 ;
        RECT 1712.650 1401.180 1712.970 1401.240 ;
        RECT 1712.650 1318.080 1712.970 1318.140 ;
        RECT 1712.455 1317.940 1712.970 1318.080 ;
        RECT 1712.650 1317.880 1712.970 1317.940 ;
        RECT 1712.650 1304.480 1712.970 1304.540 ;
        RECT 1712.455 1304.340 1712.970 1304.480 ;
        RECT 1712.650 1304.280 1712.970 1304.340 ;
        RECT 1712.205 1303.800 1712.495 1303.845 ;
        RECT 1712.650 1303.800 1712.970 1303.860 ;
        RECT 1712.205 1303.660 1712.970 1303.800 ;
        RECT 1712.205 1303.615 1712.495 1303.660 ;
        RECT 1712.650 1303.600 1712.970 1303.660 ;
        RECT 1712.190 1256.200 1712.510 1256.260 ;
        RECT 1711.995 1256.060 1712.510 1256.200 ;
        RECT 1712.190 1256.000 1712.510 1256.060 ;
        RECT 1713.570 983.180 1713.890 983.240 ;
        RECT 1714.490 983.180 1714.810 983.240 ;
        RECT 1713.570 983.040 1714.810 983.180 ;
        RECT 1713.570 982.980 1713.890 983.040 ;
        RECT 1714.490 982.980 1714.810 983.040 ;
        RECT 1711.745 862.480 1712.035 862.525 ;
        RECT 1712.650 862.480 1712.970 862.540 ;
        RECT 1711.745 862.340 1712.970 862.480 ;
        RECT 1711.745 862.295 1712.035 862.340 ;
        RECT 1712.650 862.280 1712.970 862.340 ;
        RECT 1711.730 814.540 1712.050 814.600 ;
        RECT 1711.535 814.400 1712.050 814.540 ;
        RECT 1711.730 814.340 1712.050 814.400 ;
        RECT 1712.190 627.880 1712.510 627.940 ;
        RECT 1713.110 627.880 1713.430 627.940 ;
        RECT 1712.190 627.740 1713.430 627.880 ;
        RECT 1712.190 627.680 1712.510 627.740 ;
        RECT 1713.110 627.680 1713.430 627.740 ;
        RECT 1713.110 620.740 1713.430 620.800 ;
        RECT 1712.915 620.600 1713.430 620.740 ;
        RECT 1713.110 620.540 1713.430 620.600 ;
        RECT 1713.110 572.800 1713.430 572.860 ;
        RECT 1712.915 572.660 1713.430 572.800 ;
        RECT 1713.110 572.600 1713.430 572.660 ;
        RECT 1712.650 531.660 1712.970 531.720 ;
        RECT 1713.110 531.660 1713.430 531.720 ;
        RECT 1712.650 531.520 1713.430 531.660 ;
        RECT 1712.650 531.460 1712.970 531.520 ;
        RECT 1713.110 531.460 1713.430 531.520 ;
        RECT 1712.190 448.840 1712.510 449.100 ;
        RECT 1712.280 448.420 1712.420 448.840 ;
        RECT 1712.190 448.160 1712.510 448.420 ;
        RECT 1712.650 434.760 1712.970 434.820 ;
        RECT 1712.455 434.620 1712.970 434.760 ;
        RECT 1712.650 434.560 1712.970 434.620 ;
        RECT 1712.650 400.080 1712.970 400.140 ;
        RECT 1712.455 399.940 1712.970 400.080 ;
        RECT 1712.650 399.880 1712.970 399.940 ;
        RECT 1712.205 275.980 1712.495 276.025 ;
        RECT 1712.650 275.980 1712.970 276.040 ;
        RECT 1712.205 275.840 1712.970 275.980 ;
        RECT 1712.205 275.795 1712.495 275.840 ;
        RECT 1712.650 275.780 1712.970 275.840 ;
        RECT 1712.190 228.040 1712.510 228.100 ;
        RECT 1711.995 227.900 1712.510 228.040 ;
        RECT 1712.190 227.840 1712.510 227.900 ;
        RECT 1711.745 162.080 1712.035 162.125 ;
        RECT 1712.190 162.080 1712.510 162.140 ;
        RECT 1711.745 161.940 1712.510 162.080 ;
        RECT 1711.745 161.895 1712.035 161.940 ;
        RECT 1712.190 161.880 1712.510 161.940 ;
        RECT 1711.730 96.800 1712.050 96.860 ;
        RECT 1711.535 96.660 1712.050 96.800 ;
        RECT 1711.730 96.600 1712.050 96.660 ;
        RECT 1103.610 63.480 1103.930 63.540 ;
        RECT 1711.730 63.480 1712.050 63.540 ;
        RECT 1103.610 63.340 1712.050 63.480 ;
        RECT 1103.610 63.280 1103.930 63.340 ;
        RECT 1711.730 63.280 1712.050 63.340 ;
        RECT 1102.690 2.960 1103.010 3.020 ;
        RECT 1103.610 2.960 1103.930 3.020 ;
        RECT 1102.690 2.820 1103.930 2.960 ;
        RECT 1102.690 2.760 1103.010 2.820 ;
        RECT 1103.610 2.760 1103.930 2.820 ;
      LAYER via ;
        RECT 1713.140 1642.240 1713.400 1642.500 ;
        RECT 1714.980 1642.240 1715.240 1642.500 ;
        RECT 1713.140 1546.020 1713.400 1546.280 ;
        RECT 1712.220 1545.680 1712.480 1545.940 ;
        RECT 1712.220 1545.000 1712.480 1545.260 ;
        RECT 1712.680 1497.740 1712.940 1498.000 ;
        RECT 1712.680 1414.440 1712.940 1414.700 ;
        RECT 1712.680 1401.180 1712.940 1401.440 ;
        RECT 1712.680 1317.880 1712.940 1318.140 ;
        RECT 1712.680 1304.280 1712.940 1304.540 ;
        RECT 1712.680 1303.600 1712.940 1303.860 ;
        RECT 1712.220 1256.000 1712.480 1256.260 ;
        RECT 1713.600 982.980 1713.860 983.240 ;
        RECT 1714.520 982.980 1714.780 983.240 ;
        RECT 1712.680 862.280 1712.940 862.540 ;
        RECT 1711.760 814.340 1712.020 814.600 ;
        RECT 1712.220 627.680 1712.480 627.940 ;
        RECT 1713.140 627.680 1713.400 627.940 ;
        RECT 1713.140 620.540 1713.400 620.800 ;
        RECT 1713.140 572.600 1713.400 572.860 ;
        RECT 1712.680 531.460 1712.940 531.720 ;
        RECT 1713.140 531.460 1713.400 531.720 ;
        RECT 1712.220 448.840 1712.480 449.100 ;
        RECT 1712.220 448.160 1712.480 448.420 ;
        RECT 1712.680 434.560 1712.940 434.820 ;
        RECT 1712.680 399.880 1712.940 400.140 ;
        RECT 1712.680 275.780 1712.940 276.040 ;
        RECT 1712.220 227.840 1712.480 228.100 ;
        RECT 1712.220 161.880 1712.480 162.140 ;
        RECT 1711.760 96.600 1712.020 96.860 ;
        RECT 1103.640 63.280 1103.900 63.540 ;
        RECT 1711.760 63.280 1712.020 63.540 ;
        RECT 1102.720 2.760 1102.980 3.020 ;
        RECT 1103.640 2.760 1103.900 3.020 ;
      LAYER met2 ;
        RECT 1716.280 1700.410 1716.560 1704.000 ;
        RECT 1715.040 1700.270 1716.560 1700.410 ;
        RECT 1715.040 1642.530 1715.180 1700.270 ;
        RECT 1716.280 1700.000 1716.560 1700.270 ;
        RECT 1713.140 1642.210 1713.400 1642.530 ;
        RECT 1714.980 1642.210 1715.240 1642.530 ;
        RECT 1713.200 1546.310 1713.340 1642.210 ;
        RECT 1713.140 1545.990 1713.400 1546.310 ;
        RECT 1712.220 1545.650 1712.480 1545.970 ;
        RECT 1712.280 1545.290 1712.420 1545.650 ;
        RECT 1712.220 1544.970 1712.480 1545.290 ;
        RECT 1712.680 1497.710 1712.940 1498.030 ;
        RECT 1712.740 1497.260 1712.880 1497.710 ;
        RECT 1712.740 1497.120 1713.800 1497.260 ;
        RECT 1713.660 1449.490 1713.800 1497.120 ;
        RECT 1712.740 1449.350 1713.800 1449.490 ;
        RECT 1712.740 1414.730 1712.880 1449.350 ;
        RECT 1712.680 1414.410 1712.940 1414.730 ;
        RECT 1712.680 1401.150 1712.940 1401.470 ;
        RECT 1712.740 1400.700 1712.880 1401.150 ;
        RECT 1712.740 1400.560 1713.800 1400.700 ;
        RECT 1713.660 1352.930 1713.800 1400.560 ;
        RECT 1712.740 1352.790 1713.800 1352.930 ;
        RECT 1712.740 1318.170 1712.880 1352.790 ;
        RECT 1712.680 1317.850 1712.940 1318.170 ;
        RECT 1712.680 1304.250 1712.940 1304.570 ;
        RECT 1712.740 1303.890 1712.880 1304.250 ;
        RECT 1712.680 1303.570 1712.940 1303.890 ;
        RECT 1712.220 1255.970 1712.480 1256.290 ;
        RECT 1712.280 1255.805 1712.420 1255.970 ;
        RECT 1712.210 1255.435 1712.490 1255.805 ;
        RECT 1713.130 1255.435 1713.410 1255.805 ;
        RECT 1713.200 1207.580 1713.340 1255.435 ;
        RECT 1713.200 1207.440 1713.800 1207.580 ;
        RECT 1713.660 1172.730 1713.800 1207.440 ;
        RECT 1712.280 1172.590 1713.800 1172.730 ;
        RECT 1712.280 1159.245 1712.420 1172.590 ;
        RECT 1712.210 1158.875 1712.490 1159.245 ;
        RECT 1713.590 1158.875 1713.870 1159.245 ;
        RECT 1713.660 1064.045 1713.800 1158.875 ;
        RECT 1713.590 1063.675 1713.870 1064.045 ;
        RECT 1712.210 1062.485 1712.490 1062.855 ;
        RECT 1712.280 1039.450 1712.420 1062.485 ;
        RECT 1712.280 1039.310 1713.800 1039.450 ;
        RECT 1713.660 983.270 1713.800 1039.310 ;
        RECT 1713.600 982.950 1713.860 983.270 ;
        RECT 1714.520 982.950 1714.780 983.270 ;
        RECT 1714.580 959.325 1714.720 982.950 ;
        RECT 1713.590 958.955 1713.870 959.325 ;
        RECT 1714.510 958.955 1714.790 959.325 ;
        RECT 1713.660 934.730 1713.800 958.955 ;
        RECT 1713.660 934.590 1714.720 934.730 ;
        RECT 1714.580 862.765 1714.720 934.590 ;
        RECT 1712.670 862.395 1712.950 862.765 ;
        RECT 1714.510 862.395 1714.790 862.765 ;
        RECT 1712.680 862.250 1712.940 862.395 ;
        RECT 1711.760 814.310 1712.020 814.630 ;
        RECT 1711.820 773.005 1711.960 814.310 ;
        RECT 1711.750 772.635 1712.030 773.005 ;
        RECT 1712.670 772.635 1712.950 773.005 ;
        RECT 1712.740 690.610 1712.880 772.635 ;
        RECT 1712.280 690.470 1712.880 690.610 ;
        RECT 1712.280 689.930 1712.420 690.470 ;
        RECT 1712.280 689.790 1712.880 689.930 ;
        RECT 1712.740 651.850 1712.880 689.790 ;
        RECT 1712.280 651.710 1712.880 651.850 ;
        RECT 1712.280 627.970 1712.420 651.710 ;
        RECT 1712.220 627.650 1712.480 627.970 ;
        RECT 1713.140 627.650 1713.400 627.970 ;
        RECT 1713.200 620.830 1713.340 627.650 ;
        RECT 1713.140 620.510 1713.400 620.830 ;
        RECT 1713.140 572.570 1713.400 572.890 ;
        RECT 1713.200 531.750 1713.340 572.570 ;
        RECT 1712.680 531.430 1712.940 531.750 ;
        RECT 1713.140 531.430 1713.400 531.750 ;
        RECT 1712.740 497.490 1712.880 531.430 ;
        RECT 1712.280 497.350 1712.880 497.490 ;
        RECT 1712.280 449.130 1712.420 497.350 ;
        RECT 1712.220 448.810 1712.480 449.130 ;
        RECT 1712.220 448.130 1712.480 448.450 ;
        RECT 1712.280 434.930 1712.420 448.130 ;
        RECT 1712.280 434.850 1712.880 434.930 ;
        RECT 1712.280 434.790 1712.940 434.850 ;
        RECT 1712.680 434.530 1712.940 434.790 ;
        RECT 1712.680 399.850 1712.940 400.170 ;
        RECT 1712.740 303.690 1712.880 399.850 ;
        RECT 1712.280 303.550 1712.880 303.690 ;
        RECT 1712.280 303.010 1712.420 303.550 ;
        RECT 1712.280 302.870 1712.880 303.010 ;
        RECT 1712.740 276.070 1712.880 302.870 ;
        RECT 1712.680 275.750 1712.940 276.070 ;
        RECT 1712.220 227.810 1712.480 228.130 ;
        RECT 1712.280 227.530 1712.420 227.810 ;
        RECT 1711.820 227.390 1712.420 227.530 ;
        RECT 1711.820 186.050 1711.960 227.390 ;
        RECT 1711.820 185.910 1712.420 186.050 ;
        RECT 1712.280 162.170 1712.420 185.910 ;
        RECT 1712.220 161.850 1712.480 162.170 ;
        RECT 1711.760 96.570 1712.020 96.890 ;
        RECT 1711.820 63.570 1711.960 96.570 ;
        RECT 1103.640 63.250 1103.900 63.570 ;
        RECT 1711.760 63.250 1712.020 63.570 ;
        RECT 1103.700 3.050 1103.840 63.250 ;
        RECT 1102.720 2.730 1102.980 3.050 ;
        RECT 1103.640 2.730 1103.900 3.050 ;
        RECT 1102.780 2.400 1102.920 2.730 ;
        RECT 1102.570 -4.800 1103.130 2.400 ;
      LAYER via2 ;
        RECT 1712.210 1255.480 1712.490 1255.760 ;
        RECT 1713.130 1255.480 1713.410 1255.760 ;
        RECT 1712.210 1158.920 1712.490 1159.200 ;
        RECT 1713.590 1158.920 1713.870 1159.200 ;
        RECT 1713.590 1063.720 1713.870 1064.000 ;
        RECT 1712.210 1062.530 1712.490 1062.810 ;
        RECT 1713.590 959.000 1713.870 959.280 ;
        RECT 1714.510 959.000 1714.790 959.280 ;
        RECT 1712.670 862.440 1712.950 862.720 ;
        RECT 1714.510 862.440 1714.790 862.720 ;
        RECT 1711.750 772.680 1712.030 772.960 ;
        RECT 1712.670 772.680 1712.950 772.960 ;
      LAYER met3 ;
        RECT 1712.185 1255.770 1712.515 1255.785 ;
        RECT 1713.105 1255.770 1713.435 1255.785 ;
        RECT 1712.185 1255.470 1713.435 1255.770 ;
        RECT 1712.185 1255.455 1712.515 1255.470 ;
        RECT 1713.105 1255.455 1713.435 1255.470 ;
        RECT 1712.185 1159.210 1712.515 1159.225 ;
        RECT 1713.565 1159.210 1713.895 1159.225 ;
        RECT 1712.185 1158.910 1713.895 1159.210 ;
        RECT 1712.185 1158.895 1712.515 1158.910 ;
        RECT 1713.565 1158.895 1713.895 1158.910 ;
        RECT 1713.565 1064.010 1713.895 1064.025 ;
        RECT 1711.510 1063.710 1713.895 1064.010 ;
        RECT 1711.510 1062.820 1711.810 1063.710 ;
        RECT 1713.565 1063.695 1713.895 1063.710 ;
        RECT 1712.185 1062.820 1712.515 1062.835 ;
        RECT 1711.510 1062.520 1712.515 1062.820 ;
        RECT 1712.185 1062.505 1712.515 1062.520 ;
        RECT 1713.565 959.290 1713.895 959.305 ;
        RECT 1714.485 959.290 1714.815 959.305 ;
        RECT 1713.565 958.990 1714.815 959.290 ;
        RECT 1713.565 958.975 1713.895 958.990 ;
        RECT 1714.485 958.975 1714.815 958.990 ;
        RECT 1712.645 862.730 1712.975 862.745 ;
        RECT 1714.485 862.730 1714.815 862.745 ;
        RECT 1712.645 862.430 1714.815 862.730 ;
        RECT 1712.645 862.415 1712.975 862.430 ;
        RECT 1714.485 862.415 1714.815 862.430 ;
        RECT 1711.725 772.970 1712.055 772.985 ;
        RECT 1712.645 772.970 1712.975 772.985 ;
        RECT 1711.725 772.670 1712.975 772.970 ;
        RECT 1711.725 772.655 1712.055 772.670 ;
        RECT 1712.645 772.655 1712.975 772.670 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1120.630 35.940 1120.950 36.000 ;
        RECT 1725.530 35.940 1725.850 36.000 ;
        RECT 1120.630 35.800 1725.850 35.940 ;
        RECT 1120.630 35.740 1120.950 35.800 ;
        RECT 1725.530 35.740 1725.850 35.800 ;
      LAYER via ;
        RECT 1120.660 35.740 1120.920 36.000 ;
        RECT 1725.560 35.740 1725.820 36.000 ;
      LAYER met2 ;
        RECT 1725.480 1700.000 1725.760 1704.000 ;
        RECT 1725.620 36.030 1725.760 1700.000 ;
        RECT 1120.660 35.710 1120.920 36.030 ;
        RECT 1725.560 35.710 1725.820 36.030 ;
        RECT 1120.720 2.400 1120.860 35.710 ;
        RECT 1120.510 -4.800 1121.070 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1138.570 35.600 1138.890 35.660 ;
        RECT 1731.970 35.600 1732.290 35.660 ;
        RECT 1138.570 35.460 1732.290 35.600 ;
        RECT 1138.570 35.400 1138.890 35.460 ;
        RECT 1731.970 35.400 1732.290 35.460 ;
      LAYER via ;
        RECT 1138.600 35.400 1138.860 35.660 ;
        RECT 1732.000 35.400 1732.260 35.660 ;
      LAYER met2 ;
        RECT 1734.680 1700.410 1734.960 1704.000 ;
        RECT 1732.060 1700.270 1734.960 1700.410 ;
        RECT 1732.060 35.690 1732.200 1700.270 ;
        RECT 1734.680 1700.000 1734.960 1700.270 ;
        RECT 1138.600 35.370 1138.860 35.690 ;
        RECT 1732.000 35.370 1732.260 35.690 ;
        RECT 1138.660 2.400 1138.800 35.370 ;
        RECT 1138.450 -4.800 1139.010 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1739.865 1442.025 1740.035 1490.475 ;
        RECT 1740.325 1207.425 1740.495 1250.435 ;
        RECT 1739.865 814.385 1740.035 903.975 ;
        RECT 1740.325 565.845 1740.495 572.815 ;
        RECT 1739.405 96.985 1739.575 131.155 ;
      LAYER mcon ;
        RECT 1739.865 1490.305 1740.035 1490.475 ;
        RECT 1740.325 1250.265 1740.495 1250.435 ;
        RECT 1739.865 903.805 1740.035 903.975 ;
        RECT 1740.325 572.645 1740.495 572.815 ;
        RECT 1739.405 130.985 1739.575 131.155 ;
      LAYER met1 ;
        RECT 1739.790 1683.920 1740.110 1683.980 ;
        RECT 1743.930 1683.920 1744.250 1683.980 ;
        RECT 1739.790 1683.780 1744.250 1683.920 ;
        RECT 1739.790 1683.720 1740.110 1683.780 ;
        RECT 1743.930 1683.720 1744.250 1683.780 ;
        RECT 1740.250 1621.700 1740.570 1621.760 ;
        RECT 1741.170 1621.700 1741.490 1621.760 ;
        RECT 1740.250 1621.560 1741.490 1621.700 ;
        RECT 1740.250 1621.500 1740.570 1621.560 ;
        RECT 1741.170 1621.500 1741.490 1621.560 ;
        RECT 1740.250 1608.100 1740.570 1608.160 ;
        RECT 1739.880 1607.960 1740.570 1608.100 ;
        RECT 1739.880 1607.820 1740.020 1607.960 ;
        RECT 1740.250 1607.900 1740.570 1607.960 ;
        RECT 1739.790 1607.560 1740.110 1607.820 ;
        RECT 1739.790 1497.740 1740.110 1498.000 ;
        RECT 1739.880 1496.980 1740.020 1497.740 ;
        RECT 1739.790 1496.720 1740.110 1496.980 ;
        RECT 1739.790 1490.460 1740.110 1490.520 ;
        RECT 1739.595 1490.320 1740.110 1490.460 ;
        RECT 1739.790 1490.260 1740.110 1490.320 ;
        RECT 1739.805 1442.180 1740.095 1442.225 ;
        RECT 1740.250 1442.180 1740.570 1442.240 ;
        RECT 1739.805 1442.040 1740.570 1442.180 ;
        RECT 1739.805 1441.995 1740.095 1442.040 ;
        RECT 1740.250 1441.980 1740.570 1442.040 ;
        RECT 1740.250 1400.700 1740.570 1400.760 ;
        RECT 1740.710 1400.700 1741.030 1400.760 ;
        RECT 1740.250 1400.560 1741.030 1400.700 ;
        RECT 1740.250 1400.500 1740.570 1400.560 ;
        RECT 1740.710 1400.500 1741.030 1400.560 ;
        RECT 1739.330 1338.820 1739.650 1338.880 ;
        RECT 1741.170 1338.820 1741.490 1338.880 ;
        RECT 1739.330 1338.680 1741.490 1338.820 ;
        RECT 1739.330 1338.620 1739.650 1338.680 ;
        RECT 1741.170 1338.620 1741.490 1338.680 ;
        RECT 1740.250 1250.420 1740.570 1250.480 ;
        RECT 1740.055 1250.280 1740.570 1250.420 ;
        RECT 1740.250 1250.220 1740.570 1250.280 ;
        RECT 1740.250 1207.580 1740.570 1207.640 ;
        RECT 1740.055 1207.440 1740.570 1207.580 ;
        RECT 1740.250 1207.380 1740.570 1207.440 ;
        RECT 1739.790 1152.840 1740.110 1152.900 ;
        RECT 1740.250 1152.840 1740.570 1152.900 ;
        RECT 1739.790 1152.700 1740.570 1152.840 ;
        RECT 1739.790 1152.640 1740.110 1152.700 ;
        RECT 1740.250 1152.640 1740.570 1152.700 ;
        RECT 1739.790 1124.760 1740.110 1125.020 ;
        RECT 1739.880 1124.280 1740.020 1124.760 ;
        RECT 1740.250 1124.280 1740.570 1124.340 ;
        RECT 1739.880 1124.140 1740.570 1124.280 ;
        RECT 1740.250 1124.080 1740.570 1124.140 ;
        RECT 1739.790 1062.740 1740.110 1062.800 ;
        RECT 1740.710 1062.740 1741.030 1062.800 ;
        RECT 1739.790 1062.600 1741.030 1062.740 ;
        RECT 1739.790 1062.540 1740.110 1062.600 ;
        RECT 1740.710 1062.540 1741.030 1062.600 ;
        RECT 1739.790 1028.200 1740.110 1028.460 ;
        RECT 1739.880 1028.060 1740.020 1028.200 ;
        RECT 1740.250 1028.060 1740.570 1028.120 ;
        RECT 1739.880 1027.920 1740.570 1028.060 ;
        RECT 1740.250 1027.860 1740.570 1027.920 ;
        RECT 1739.790 966.180 1740.110 966.240 ;
        RECT 1740.710 966.180 1741.030 966.240 ;
        RECT 1739.790 966.040 1741.030 966.180 ;
        RECT 1739.790 965.980 1740.110 966.040 ;
        RECT 1740.710 965.980 1741.030 966.040 ;
        RECT 1739.790 917.900 1740.110 917.960 ;
        RECT 1740.250 917.900 1740.570 917.960 ;
        RECT 1739.790 917.760 1740.570 917.900 ;
        RECT 1739.790 917.700 1740.110 917.760 ;
        RECT 1740.250 917.700 1740.570 917.760 ;
        RECT 1739.805 903.960 1740.095 904.005 ;
        RECT 1740.250 903.960 1740.570 904.020 ;
        RECT 1739.805 903.820 1740.570 903.960 ;
        RECT 1739.805 903.775 1740.095 903.820 ;
        RECT 1740.250 903.760 1740.570 903.820 ;
        RECT 1739.790 814.540 1740.110 814.600 ;
        RECT 1739.595 814.400 1740.110 814.540 ;
        RECT 1739.790 814.340 1740.110 814.400 ;
        RECT 1739.790 724.440 1740.110 724.500 ;
        RECT 1740.250 724.440 1740.570 724.500 ;
        RECT 1739.790 724.300 1740.570 724.440 ;
        RECT 1739.790 724.240 1740.110 724.300 ;
        RECT 1740.250 724.240 1740.570 724.300 ;
        RECT 1739.790 628.020 1740.110 628.280 ;
        RECT 1739.880 627.540 1740.020 628.020 ;
        RECT 1740.250 627.540 1740.570 627.600 ;
        RECT 1739.880 627.400 1740.570 627.540 ;
        RECT 1740.250 627.340 1740.570 627.400 ;
        RECT 1740.250 572.800 1740.570 572.860 ;
        RECT 1740.055 572.660 1740.570 572.800 ;
        RECT 1740.250 572.600 1740.570 572.660 ;
        RECT 1740.250 566.000 1740.570 566.060 ;
        RECT 1740.055 565.860 1740.570 566.000 ;
        RECT 1740.250 565.800 1740.570 565.860 ;
        RECT 1739.330 524.520 1739.650 524.580 ;
        RECT 1740.250 524.520 1740.570 524.580 ;
        RECT 1739.330 524.380 1740.570 524.520 ;
        RECT 1739.330 524.320 1739.650 524.380 ;
        RECT 1740.250 524.320 1740.570 524.380 ;
        RECT 1739.330 427.960 1739.650 428.020 ;
        RECT 1740.250 427.960 1740.570 428.020 ;
        RECT 1739.330 427.820 1740.570 427.960 ;
        RECT 1739.330 427.760 1739.650 427.820 ;
        RECT 1740.250 427.760 1740.570 427.820 ;
        RECT 1740.250 386.820 1740.570 386.880 ;
        RECT 1739.880 386.680 1740.570 386.820 ;
        RECT 1739.880 386.540 1740.020 386.680 ;
        RECT 1740.250 386.620 1740.570 386.680 ;
        RECT 1739.790 386.280 1740.110 386.540 ;
        RECT 1739.790 304.000 1740.110 304.260 ;
        RECT 1739.880 303.580 1740.020 304.000 ;
        RECT 1739.790 303.320 1740.110 303.580 ;
        RECT 1739.790 234.840 1740.110 234.900 ;
        RECT 1740.710 234.840 1741.030 234.900 ;
        RECT 1739.790 234.700 1741.030 234.840 ;
        RECT 1739.790 234.640 1740.110 234.700 ;
        RECT 1740.710 234.640 1741.030 234.700 ;
        RECT 1739.330 179.760 1739.650 179.820 ;
        RECT 1740.710 179.760 1741.030 179.820 ;
        RECT 1739.330 179.620 1741.030 179.760 ;
        RECT 1739.330 179.560 1739.650 179.620 ;
        RECT 1740.710 179.560 1741.030 179.620 ;
        RECT 1739.330 131.140 1739.650 131.200 ;
        RECT 1739.135 131.000 1739.650 131.140 ;
        RECT 1739.330 130.940 1739.650 131.000 ;
        RECT 1739.345 97.140 1739.635 97.185 ;
        RECT 1739.790 97.140 1740.110 97.200 ;
        RECT 1739.345 97.000 1740.110 97.140 ;
        RECT 1739.345 96.955 1739.635 97.000 ;
        RECT 1739.790 96.940 1740.110 97.000 ;
        RECT 1739.790 62.460 1740.110 62.520 ;
        RECT 1739.420 62.320 1740.110 62.460 ;
        RECT 1739.420 62.180 1739.560 62.320 ;
        RECT 1739.790 62.260 1740.110 62.320 ;
        RECT 1739.330 61.920 1739.650 62.180 ;
        RECT 1156.510 37.980 1156.830 38.040 ;
        RECT 1739.330 37.980 1739.650 38.040 ;
        RECT 1156.510 37.840 1739.650 37.980 ;
        RECT 1156.510 37.780 1156.830 37.840 ;
        RECT 1739.330 37.780 1739.650 37.840 ;
      LAYER via ;
        RECT 1739.820 1683.720 1740.080 1683.980 ;
        RECT 1743.960 1683.720 1744.220 1683.980 ;
        RECT 1740.280 1621.500 1740.540 1621.760 ;
        RECT 1741.200 1621.500 1741.460 1621.760 ;
        RECT 1740.280 1607.900 1740.540 1608.160 ;
        RECT 1739.820 1607.560 1740.080 1607.820 ;
        RECT 1739.820 1497.740 1740.080 1498.000 ;
        RECT 1739.820 1496.720 1740.080 1496.980 ;
        RECT 1739.820 1490.260 1740.080 1490.520 ;
        RECT 1740.280 1441.980 1740.540 1442.240 ;
        RECT 1740.280 1400.500 1740.540 1400.760 ;
        RECT 1740.740 1400.500 1741.000 1400.760 ;
        RECT 1739.360 1338.620 1739.620 1338.880 ;
        RECT 1741.200 1338.620 1741.460 1338.880 ;
        RECT 1740.280 1250.220 1740.540 1250.480 ;
        RECT 1740.280 1207.380 1740.540 1207.640 ;
        RECT 1739.820 1152.640 1740.080 1152.900 ;
        RECT 1740.280 1152.640 1740.540 1152.900 ;
        RECT 1739.820 1124.760 1740.080 1125.020 ;
        RECT 1740.280 1124.080 1740.540 1124.340 ;
        RECT 1739.820 1062.540 1740.080 1062.800 ;
        RECT 1740.740 1062.540 1741.000 1062.800 ;
        RECT 1739.820 1028.200 1740.080 1028.460 ;
        RECT 1740.280 1027.860 1740.540 1028.120 ;
        RECT 1739.820 965.980 1740.080 966.240 ;
        RECT 1740.740 965.980 1741.000 966.240 ;
        RECT 1739.820 917.700 1740.080 917.960 ;
        RECT 1740.280 917.700 1740.540 917.960 ;
        RECT 1740.280 903.760 1740.540 904.020 ;
        RECT 1739.820 814.340 1740.080 814.600 ;
        RECT 1739.820 724.240 1740.080 724.500 ;
        RECT 1740.280 724.240 1740.540 724.500 ;
        RECT 1739.820 628.020 1740.080 628.280 ;
        RECT 1740.280 627.340 1740.540 627.600 ;
        RECT 1740.280 572.600 1740.540 572.860 ;
        RECT 1740.280 565.800 1740.540 566.060 ;
        RECT 1739.360 524.320 1739.620 524.580 ;
        RECT 1740.280 524.320 1740.540 524.580 ;
        RECT 1739.360 427.760 1739.620 428.020 ;
        RECT 1740.280 427.760 1740.540 428.020 ;
        RECT 1740.280 386.620 1740.540 386.880 ;
        RECT 1739.820 386.280 1740.080 386.540 ;
        RECT 1739.820 304.000 1740.080 304.260 ;
        RECT 1739.820 303.320 1740.080 303.580 ;
        RECT 1739.820 234.640 1740.080 234.900 ;
        RECT 1740.740 234.640 1741.000 234.900 ;
        RECT 1739.360 179.560 1739.620 179.820 ;
        RECT 1740.740 179.560 1741.000 179.820 ;
        RECT 1739.360 130.940 1739.620 131.200 ;
        RECT 1739.820 96.940 1740.080 97.200 ;
        RECT 1739.820 62.260 1740.080 62.520 ;
        RECT 1739.360 61.920 1739.620 62.180 ;
        RECT 1156.540 37.780 1156.800 38.040 ;
        RECT 1739.360 37.780 1739.620 38.040 ;
      LAYER met2 ;
        RECT 1743.880 1700.000 1744.160 1704.000 ;
        RECT 1744.020 1684.010 1744.160 1700.000 ;
        RECT 1739.820 1683.690 1740.080 1684.010 ;
        RECT 1743.960 1683.690 1744.220 1684.010 ;
        RECT 1739.880 1669.925 1740.020 1683.690 ;
        RECT 1739.810 1669.555 1740.090 1669.925 ;
        RECT 1741.190 1669.555 1741.470 1669.925 ;
        RECT 1741.260 1621.790 1741.400 1669.555 ;
        RECT 1740.280 1621.470 1740.540 1621.790 ;
        RECT 1741.200 1621.470 1741.460 1621.790 ;
        RECT 1740.340 1608.190 1740.480 1621.470 ;
        RECT 1740.280 1607.870 1740.540 1608.190 ;
        RECT 1739.820 1607.530 1740.080 1607.850 ;
        RECT 1739.880 1498.030 1740.020 1607.530 ;
        RECT 1739.820 1497.710 1740.080 1498.030 ;
        RECT 1739.820 1496.690 1740.080 1497.010 ;
        RECT 1739.880 1490.550 1740.020 1496.690 ;
        RECT 1739.820 1490.230 1740.080 1490.550 ;
        RECT 1740.280 1441.950 1740.540 1442.270 ;
        RECT 1740.340 1400.790 1740.480 1441.950 ;
        RECT 1740.280 1400.470 1740.540 1400.790 ;
        RECT 1740.740 1400.470 1741.000 1400.790 ;
        RECT 1740.800 1352.930 1740.940 1400.470 ;
        RECT 1740.800 1352.790 1741.400 1352.930 ;
        RECT 1741.260 1338.910 1741.400 1352.790 ;
        RECT 1739.360 1338.765 1739.620 1338.910 ;
        RECT 1738.430 1338.395 1738.710 1338.765 ;
        RECT 1739.350 1338.395 1739.630 1338.765 ;
        RECT 1741.200 1338.590 1741.460 1338.910 ;
        RECT 1738.500 1290.485 1738.640 1338.395 ;
        RECT 1738.430 1290.115 1738.710 1290.485 ;
        RECT 1740.270 1290.115 1740.550 1290.485 ;
        RECT 1740.340 1250.510 1740.480 1290.115 ;
        RECT 1740.280 1250.190 1740.540 1250.510 ;
        RECT 1740.280 1207.350 1740.540 1207.670 ;
        RECT 1740.340 1152.930 1740.480 1207.350 ;
        RECT 1739.820 1152.610 1740.080 1152.930 ;
        RECT 1740.280 1152.610 1740.540 1152.930 ;
        RECT 1739.880 1125.050 1740.020 1152.610 ;
        RECT 1739.820 1124.730 1740.080 1125.050 ;
        RECT 1740.280 1124.050 1740.540 1124.370 ;
        RECT 1740.340 1087.050 1740.480 1124.050 ;
        RECT 1740.340 1086.910 1740.940 1087.050 ;
        RECT 1740.800 1062.830 1740.940 1086.910 ;
        RECT 1739.820 1062.510 1740.080 1062.830 ;
        RECT 1740.740 1062.510 1741.000 1062.830 ;
        RECT 1739.880 1028.490 1740.020 1062.510 ;
        RECT 1739.820 1028.170 1740.080 1028.490 ;
        RECT 1740.280 1027.830 1740.540 1028.150 ;
        RECT 1740.340 990.490 1740.480 1027.830 ;
        RECT 1740.340 990.350 1740.940 990.490 ;
        RECT 1740.800 966.270 1740.940 990.350 ;
        RECT 1739.820 965.950 1740.080 966.270 ;
        RECT 1740.740 965.950 1741.000 966.270 ;
        RECT 1739.880 917.990 1740.020 965.950 ;
        RECT 1739.820 917.670 1740.080 917.990 ;
        RECT 1740.280 917.670 1740.540 917.990 ;
        RECT 1740.340 904.050 1740.480 917.670 ;
        RECT 1740.280 903.730 1740.540 904.050 ;
        RECT 1739.820 814.310 1740.080 814.630 ;
        RECT 1739.880 766.090 1740.020 814.310 ;
        RECT 1739.880 765.950 1740.480 766.090 ;
        RECT 1740.340 724.530 1740.480 765.950 ;
        RECT 1739.820 724.210 1740.080 724.530 ;
        RECT 1740.280 724.210 1740.540 724.530 ;
        RECT 1739.880 670.325 1740.020 724.210 ;
        RECT 1739.810 669.955 1740.090 670.325 ;
        RECT 1739.810 669.275 1740.090 669.645 ;
        RECT 1739.880 628.310 1740.020 669.275 ;
        RECT 1739.820 627.990 1740.080 628.310 ;
        RECT 1740.280 627.310 1740.540 627.630 ;
        RECT 1740.340 572.890 1740.480 627.310 ;
        RECT 1740.280 572.570 1740.540 572.890 ;
        RECT 1740.280 565.770 1740.540 566.090 ;
        RECT 1740.340 524.610 1740.480 565.770 ;
        RECT 1739.360 524.290 1739.620 524.610 ;
        RECT 1740.280 524.290 1740.540 524.610 ;
        RECT 1739.420 428.050 1739.560 524.290 ;
        RECT 1739.360 427.730 1739.620 428.050 ;
        RECT 1740.280 427.730 1740.540 428.050 ;
        RECT 1740.340 386.910 1740.480 427.730 ;
        RECT 1740.280 386.590 1740.540 386.910 ;
        RECT 1739.820 386.250 1740.080 386.570 ;
        RECT 1739.880 304.290 1740.020 386.250 ;
        RECT 1739.820 303.970 1740.080 304.290 ;
        RECT 1739.820 303.290 1740.080 303.610 ;
        RECT 1739.880 234.930 1740.020 303.290 ;
        RECT 1739.820 234.610 1740.080 234.930 ;
        RECT 1740.740 234.610 1741.000 234.930 ;
        RECT 1740.800 179.850 1740.940 234.610 ;
        RECT 1739.360 179.530 1739.620 179.850 ;
        RECT 1740.740 179.530 1741.000 179.850 ;
        RECT 1739.420 131.230 1739.560 179.530 ;
        RECT 1739.360 130.910 1739.620 131.230 ;
        RECT 1739.820 96.910 1740.080 97.230 ;
        RECT 1739.880 62.550 1740.020 96.910 ;
        RECT 1739.820 62.230 1740.080 62.550 ;
        RECT 1739.360 61.890 1739.620 62.210 ;
        RECT 1739.420 38.070 1739.560 61.890 ;
        RECT 1156.540 37.750 1156.800 38.070 ;
        RECT 1739.360 37.750 1739.620 38.070 ;
        RECT 1156.600 2.400 1156.740 37.750 ;
        RECT 1156.390 -4.800 1156.950 2.400 ;
      LAYER via2 ;
        RECT 1739.810 1669.600 1740.090 1669.880 ;
        RECT 1741.190 1669.600 1741.470 1669.880 ;
        RECT 1738.430 1338.440 1738.710 1338.720 ;
        RECT 1739.350 1338.440 1739.630 1338.720 ;
        RECT 1738.430 1290.160 1738.710 1290.440 ;
        RECT 1740.270 1290.160 1740.550 1290.440 ;
        RECT 1739.810 670.000 1740.090 670.280 ;
        RECT 1739.810 669.320 1740.090 669.600 ;
      LAYER met3 ;
        RECT 1739.785 1669.890 1740.115 1669.905 ;
        RECT 1741.165 1669.890 1741.495 1669.905 ;
        RECT 1739.785 1669.590 1741.495 1669.890 ;
        RECT 1739.785 1669.575 1740.115 1669.590 ;
        RECT 1741.165 1669.575 1741.495 1669.590 ;
        RECT 1738.405 1338.730 1738.735 1338.745 ;
        RECT 1739.325 1338.730 1739.655 1338.745 ;
        RECT 1738.405 1338.430 1739.655 1338.730 ;
        RECT 1738.405 1338.415 1738.735 1338.430 ;
        RECT 1739.325 1338.415 1739.655 1338.430 ;
        RECT 1738.405 1290.450 1738.735 1290.465 ;
        RECT 1740.245 1290.450 1740.575 1290.465 ;
        RECT 1738.405 1290.150 1740.575 1290.450 ;
        RECT 1738.405 1290.135 1738.735 1290.150 ;
        RECT 1740.245 1290.135 1740.575 1290.150 ;
        RECT 1739.785 670.290 1740.115 670.305 ;
        RECT 1739.785 669.975 1740.330 670.290 ;
        RECT 1740.030 669.625 1740.330 669.975 ;
        RECT 1739.785 669.310 1740.330 669.625 ;
        RECT 1739.785 669.295 1740.115 669.310 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1491.925 1435.225 1492.095 1483.335 ;
        RECT 1491.465 917.745 1491.635 932.195 ;
        RECT 1491.465 786.505 1491.635 814.215 ;
        RECT 1491.005 559.045 1491.175 593.895 ;
        RECT 1491.925 510.765 1492.095 558.535 ;
        RECT 1491.925 468.945 1492.095 497.335 ;
        RECT 1492.845 421.005 1493.015 444.975 ;
      LAYER mcon ;
        RECT 1491.925 1483.165 1492.095 1483.335 ;
        RECT 1491.465 932.025 1491.635 932.195 ;
        RECT 1491.465 814.045 1491.635 814.215 ;
        RECT 1491.005 593.725 1491.175 593.895 ;
        RECT 1491.925 558.365 1492.095 558.535 ;
        RECT 1491.925 497.165 1492.095 497.335 ;
        RECT 1492.845 444.805 1493.015 444.975 ;
      LAYER met1 ;
        RECT 1491.390 1511.340 1491.710 1511.600 ;
        RECT 1491.480 1510.520 1491.620 1511.340 ;
        RECT 1491.850 1510.520 1492.170 1510.580 ;
        RECT 1491.480 1510.380 1492.170 1510.520 ;
        RECT 1491.850 1510.320 1492.170 1510.380 ;
        RECT 1491.850 1483.320 1492.170 1483.380 ;
        RECT 1491.655 1483.180 1492.170 1483.320 ;
        RECT 1491.850 1483.120 1492.170 1483.180 ;
        RECT 1491.865 1435.380 1492.155 1435.425 ;
        RECT 1492.310 1435.380 1492.630 1435.440 ;
        RECT 1491.865 1435.240 1492.630 1435.380 ;
        RECT 1491.865 1435.195 1492.155 1435.240 ;
        RECT 1492.310 1435.180 1492.630 1435.240 ;
        RECT 1492.310 1400.700 1492.630 1400.760 ;
        RECT 1491.480 1400.560 1492.630 1400.700 ;
        RECT 1491.480 1400.420 1491.620 1400.560 ;
        RECT 1492.310 1400.500 1492.630 1400.560 ;
        RECT 1491.390 1400.160 1491.710 1400.420 ;
        RECT 1491.390 1255.860 1491.710 1255.920 ;
        RECT 1492.770 1255.860 1493.090 1255.920 ;
        RECT 1491.390 1255.720 1493.090 1255.860 ;
        RECT 1491.390 1255.660 1491.710 1255.720 ;
        RECT 1492.770 1255.660 1493.090 1255.720 ;
        RECT 1491.390 1159.300 1491.710 1159.360 ;
        RECT 1492.770 1159.300 1493.090 1159.360 ;
        RECT 1491.390 1159.160 1493.090 1159.300 ;
        RECT 1491.390 1159.100 1491.710 1159.160 ;
        RECT 1492.770 1159.100 1493.090 1159.160 ;
        RECT 1491.390 1111.020 1491.710 1111.080 ;
        RECT 1492.770 1111.020 1493.090 1111.080 ;
        RECT 1491.390 1110.880 1493.090 1111.020 ;
        RECT 1491.390 1110.820 1491.710 1110.880 ;
        RECT 1492.770 1110.820 1493.090 1110.880 ;
        RECT 1491.390 1062.740 1491.710 1062.800 ;
        RECT 1492.770 1062.740 1493.090 1062.800 ;
        RECT 1491.390 1062.600 1493.090 1062.740 ;
        RECT 1491.390 1062.540 1491.710 1062.600 ;
        RECT 1492.770 1062.540 1493.090 1062.600 ;
        RECT 1491.390 1028.200 1491.710 1028.460 ;
        RECT 1491.480 1028.060 1491.620 1028.200 ;
        RECT 1491.850 1028.060 1492.170 1028.120 ;
        RECT 1491.480 1027.920 1492.170 1028.060 ;
        RECT 1491.850 1027.860 1492.170 1027.920 ;
        RECT 1491.390 966.180 1491.710 966.240 ;
        RECT 1492.310 966.180 1492.630 966.240 ;
        RECT 1491.390 966.040 1492.630 966.180 ;
        RECT 1491.390 965.980 1491.710 966.040 ;
        RECT 1492.310 965.980 1492.630 966.040 ;
        RECT 1491.390 932.180 1491.710 932.240 ;
        RECT 1491.195 932.040 1491.710 932.180 ;
        RECT 1491.390 931.980 1491.710 932.040 ;
        RECT 1491.390 917.900 1491.710 917.960 ;
        RECT 1491.195 917.760 1491.710 917.900 ;
        RECT 1491.390 917.700 1491.710 917.760 ;
        RECT 1491.390 910.760 1491.710 910.820 ;
        RECT 1492.310 910.760 1492.630 910.820 ;
        RECT 1491.390 910.620 1492.630 910.760 ;
        RECT 1491.390 910.560 1491.710 910.620 ;
        RECT 1492.310 910.560 1492.630 910.620 ;
        RECT 1490.930 821.340 1491.250 821.400 ;
        RECT 1491.390 821.340 1491.710 821.400 ;
        RECT 1490.930 821.200 1491.710 821.340 ;
        RECT 1490.930 821.140 1491.250 821.200 ;
        RECT 1491.390 821.140 1491.710 821.200 ;
        RECT 1491.390 814.200 1491.710 814.260 ;
        RECT 1491.195 814.060 1491.710 814.200 ;
        RECT 1491.390 814.000 1491.710 814.060 ;
        RECT 1491.390 786.660 1491.710 786.720 ;
        RECT 1491.195 786.520 1491.710 786.660 ;
        RECT 1491.390 786.460 1491.710 786.520 ;
        RECT 1491.390 724.440 1491.710 724.500 ;
        RECT 1492.310 724.440 1492.630 724.500 ;
        RECT 1491.390 724.300 1492.630 724.440 ;
        RECT 1491.390 724.240 1491.710 724.300 ;
        RECT 1492.310 724.240 1492.630 724.300 ;
        RECT 1490.945 593.880 1491.235 593.925 ;
        RECT 1491.390 593.880 1491.710 593.940 ;
        RECT 1490.945 593.740 1491.710 593.880 ;
        RECT 1490.945 593.695 1491.235 593.740 ;
        RECT 1491.390 593.680 1491.710 593.740 ;
        RECT 1490.945 559.015 1491.235 559.245 ;
        RECT 1491.020 558.520 1491.160 559.015 ;
        RECT 1491.865 558.520 1492.155 558.565 ;
        RECT 1491.020 558.380 1492.155 558.520 ;
        RECT 1491.865 558.335 1492.155 558.380 ;
        RECT 1491.850 510.920 1492.170 510.980 ;
        RECT 1491.655 510.780 1492.170 510.920 ;
        RECT 1491.850 510.720 1492.170 510.780 ;
        RECT 1491.850 497.320 1492.170 497.380 ;
        RECT 1491.655 497.180 1492.170 497.320 ;
        RECT 1491.850 497.120 1492.170 497.180 ;
        RECT 1491.850 469.100 1492.170 469.160 ;
        RECT 1491.655 468.960 1492.170 469.100 ;
        RECT 1491.850 468.900 1492.170 468.960 ;
        RECT 1491.850 444.960 1492.170 445.020 ;
        RECT 1492.785 444.960 1493.075 445.005 ;
        RECT 1491.850 444.820 1493.075 444.960 ;
        RECT 1491.850 444.760 1492.170 444.820 ;
        RECT 1492.785 444.775 1493.075 444.820 ;
        RECT 1492.770 421.160 1493.090 421.220 ;
        RECT 1492.770 421.020 1493.285 421.160 ;
        RECT 1492.770 420.960 1493.090 421.020 ;
        RECT 1491.390 289.720 1491.710 289.980 ;
        RECT 1491.480 289.240 1491.620 289.720 ;
        RECT 1491.850 289.240 1492.170 289.300 ;
        RECT 1491.480 289.100 1492.170 289.240 ;
        RECT 1491.850 289.040 1492.170 289.100 ;
        RECT 1491.850 275.980 1492.170 276.040 ;
        RECT 1492.310 275.980 1492.630 276.040 ;
        RECT 1491.850 275.840 1492.630 275.980 ;
        RECT 1491.850 275.780 1492.170 275.840 ;
        RECT 1492.310 275.780 1492.630 275.840 ;
      LAYER via ;
        RECT 1491.420 1511.340 1491.680 1511.600 ;
        RECT 1491.880 1510.320 1492.140 1510.580 ;
        RECT 1491.880 1483.120 1492.140 1483.380 ;
        RECT 1492.340 1435.180 1492.600 1435.440 ;
        RECT 1492.340 1400.500 1492.600 1400.760 ;
        RECT 1491.420 1400.160 1491.680 1400.420 ;
        RECT 1491.420 1255.660 1491.680 1255.920 ;
        RECT 1492.800 1255.660 1493.060 1255.920 ;
        RECT 1491.420 1159.100 1491.680 1159.360 ;
        RECT 1492.800 1159.100 1493.060 1159.360 ;
        RECT 1491.420 1110.820 1491.680 1111.080 ;
        RECT 1492.800 1110.820 1493.060 1111.080 ;
        RECT 1491.420 1062.540 1491.680 1062.800 ;
        RECT 1492.800 1062.540 1493.060 1062.800 ;
        RECT 1491.420 1028.200 1491.680 1028.460 ;
        RECT 1491.880 1027.860 1492.140 1028.120 ;
        RECT 1491.420 965.980 1491.680 966.240 ;
        RECT 1492.340 965.980 1492.600 966.240 ;
        RECT 1491.420 931.980 1491.680 932.240 ;
        RECT 1491.420 917.700 1491.680 917.960 ;
        RECT 1491.420 910.560 1491.680 910.820 ;
        RECT 1492.340 910.560 1492.600 910.820 ;
        RECT 1490.960 821.140 1491.220 821.400 ;
        RECT 1491.420 821.140 1491.680 821.400 ;
        RECT 1491.420 814.000 1491.680 814.260 ;
        RECT 1491.420 786.460 1491.680 786.720 ;
        RECT 1491.420 724.240 1491.680 724.500 ;
        RECT 1492.340 724.240 1492.600 724.500 ;
        RECT 1491.420 593.680 1491.680 593.940 ;
        RECT 1491.880 510.720 1492.140 510.980 ;
        RECT 1491.880 497.120 1492.140 497.380 ;
        RECT 1491.880 468.900 1492.140 469.160 ;
        RECT 1491.880 444.760 1492.140 445.020 ;
        RECT 1492.800 420.960 1493.060 421.220 ;
        RECT 1491.420 289.720 1491.680 289.980 ;
        RECT 1491.880 289.040 1492.140 289.300 ;
        RECT 1491.880 275.780 1492.140 276.040 ;
        RECT 1492.340 275.780 1492.600 276.040 ;
      LAYER met2 ;
        RECT 1495.940 1700.410 1496.220 1704.000 ;
        RECT 1493.780 1700.270 1496.220 1700.410 ;
        RECT 1493.780 1656.210 1493.920 1700.270 ;
        RECT 1495.940 1700.000 1496.220 1700.270 ;
        RECT 1491.940 1656.070 1493.920 1656.210 ;
        RECT 1491.940 1559.650 1492.080 1656.070 ;
        RECT 1491.480 1559.510 1492.080 1559.650 ;
        RECT 1491.480 1511.630 1491.620 1559.510 ;
        RECT 1491.420 1511.310 1491.680 1511.630 ;
        RECT 1491.880 1510.290 1492.140 1510.610 ;
        RECT 1491.940 1483.410 1492.080 1510.290 ;
        RECT 1491.880 1483.090 1492.140 1483.410 ;
        RECT 1492.340 1435.150 1492.600 1435.470 ;
        RECT 1492.400 1400.790 1492.540 1435.150 ;
        RECT 1492.340 1400.470 1492.600 1400.790 ;
        RECT 1491.420 1400.130 1491.680 1400.450 ;
        RECT 1491.480 1393.845 1491.620 1400.130 ;
        RECT 1491.410 1393.475 1491.690 1393.845 ;
        RECT 1492.790 1393.475 1493.070 1393.845 ;
        RECT 1492.860 1269.290 1493.000 1393.475 ;
        RECT 1491.480 1269.150 1493.000 1269.290 ;
        RECT 1491.480 1255.950 1491.620 1269.150 ;
        RECT 1491.420 1255.630 1491.680 1255.950 ;
        RECT 1492.800 1255.630 1493.060 1255.950 ;
        RECT 1492.860 1159.390 1493.000 1255.630 ;
        RECT 1491.420 1159.070 1491.680 1159.390 ;
        RECT 1492.800 1159.070 1493.060 1159.390 ;
        RECT 1491.480 1111.110 1491.620 1159.070 ;
        RECT 1491.420 1110.790 1491.680 1111.110 ;
        RECT 1492.800 1110.790 1493.060 1111.110 ;
        RECT 1492.860 1062.830 1493.000 1110.790 ;
        RECT 1491.420 1062.510 1491.680 1062.830 ;
        RECT 1492.800 1062.510 1493.060 1062.830 ;
        RECT 1491.480 1028.490 1491.620 1062.510 ;
        RECT 1491.420 1028.170 1491.680 1028.490 ;
        RECT 1491.880 1027.830 1492.140 1028.150 ;
        RECT 1491.940 990.490 1492.080 1027.830 ;
        RECT 1491.940 990.350 1492.540 990.490 ;
        RECT 1492.400 966.270 1492.540 990.350 ;
        RECT 1491.420 965.950 1491.680 966.270 ;
        RECT 1492.340 965.950 1492.600 966.270 ;
        RECT 1491.480 932.270 1491.620 965.950 ;
        RECT 1491.420 931.950 1491.680 932.270 ;
        RECT 1491.420 917.670 1491.680 917.990 ;
        RECT 1491.480 910.850 1491.620 917.670 ;
        RECT 1491.420 910.530 1491.680 910.850 ;
        RECT 1492.340 910.530 1492.600 910.850 ;
        RECT 1492.400 862.765 1492.540 910.530 ;
        RECT 1490.950 862.395 1491.230 862.765 ;
        RECT 1492.330 862.395 1492.610 862.765 ;
        RECT 1491.020 821.430 1491.160 862.395 ;
        RECT 1490.960 821.110 1491.220 821.430 ;
        RECT 1491.420 821.110 1491.680 821.430 ;
        RECT 1491.480 814.290 1491.620 821.110 ;
        RECT 1491.420 813.970 1491.680 814.290 ;
        RECT 1491.420 786.430 1491.680 786.750 ;
        RECT 1491.480 766.090 1491.620 786.430 ;
        RECT 1491.480 765.950 1492.080 766.090 ;
        RECT 1491.940 749.090 1492.080 765.950 ;
        RECT 1491.940 748.950 1492.540 749.090 ;
        RECT 1492.400 724.725 1492.540 748.950 ;
        RECT 1491.410 724.355 1491.690 724.725 ;
        RECT 1492.330 724.355 1492.610 724.725 ;
        RECT 1491.420 724.210 1491.680 724.355 ;
        RECT 1492.340 724.210 1492.600 724.355 ;
        RECT 1492.400 699.450 1492.540 724.210 ;
        RECT 1491.940 699.310 1492.540 699.450 ;
        RECT 1491.940 621.250 1492.080 699.310 ;
        RECT 1491.480 621.110 1492.080 621.250 ;
        RECT 1491.480 593.970 1491.620 621.110 ;
        RECT 1491.420 593.650 1491.680 593.970 ;
        RECT 1491.880 510.690 1492.140 511.010 ;
        RECT 1491.940 497.410 1492.080 510.690 ;
        RECT 1491.880 497.090 1492.140 497.410 ;
        RECT 1491.880 468.870 1492.140 469.190 ;
        RECT 1491.940 445.050 1492.080 468.870 ;
        RECT 1491.880 444.730 1492.140 445.050 ;
        RECT 1492.800 420.930 1493.060 421.250 ;
        RECT 1492.860 379.965 1493.000 420.930 ;
        RECT 1491.410 379.595 1491.690 379.965 ;
        RECT 1492.790 379.595 1493.070 379.965 ;
        RECT 1491.480 290.010 1491.620 379.595 ;
        RECT 1491.420 289.690 1491.680 290.010 ;
        RECT 1491.880 289.010 1492.140 289.330 ;
        RECT 1491.940 276.070 1492.080 289.010 ;
        RECT 1491.880 275.750 1492.140 276.070 ;
        RECT 1492.340 275.750 1492.600 276.070 ;
        RECT 1492.400 60.930 1492.540 275.750 ;
        RECT 1491.020 60.790 1492.540 60.930 ;
        RECT 1491.020 48.010 1491.160 60.790 ;
        RECT 1491.020 47.870 1491.620 48.010 ;
        RECT 1491.480 37.925 1491.620 47.870 ;
        RECT 674.450 37.555 674.730 37.925 ;
        RECT 1491.410 37.555 1491.690 37.925 ;
        RECT 674.520 2.400 674.660 37.555 ;
        RECT 674.310 -4.800 674.870 2.400 ;
      LAYER via2 ;
        RECT 1491.410 1393.520 1491.690 1393.800 ;
        RECT 1492.790 1393.520 1493.070 1393.800 ;
        RECT 1490.950 862.440 1491.230 862.720 ;
        RECT 1492.330 862.440 1492.610 862.720 ;
        RECT 1491.410 724.400 1491.690 724.680 ;
        RECT 1492.330 724.400 1492.610 724.680 ;
        RECT 1491.410 379.640 1491.690 379.920 ;
        RECT 1492.790 379.640 1493.070 379.920 ;
        RECT 674.450 37.600 674.730 37.880 ;
        RECT 1491.410 37.600 1491.690 37.880 ;
      LAYER met3 ;
        RECT 1491.385 1393.810 1491.715 1393.825 ;
        RECT 1492.765 1393.810 1493.095 1393.825 ;
        RECT 1491.385 1393.510 1493.095 1393.810 ;
        RECT 1491.385 1393.495 1491.715 1393.510 ;
        RECT 1492.765 1393.495 1493.095 1393.510 ;
        RECT 1490.925 862.730 1491.255 862.745 ;
        RECT 1492.305 862.730 1492.635 862.745 ;
        RECT 1490.925 862.430 1492.635 862.730 ;
        RECT 1490.925 862.415 1491.255 862.430 ;
        RECT 1492.305 862.415 1492.635 862.430 ;
        RECT 1491.385 724.690 1491.715 724.705 ;
        RECT 1492.305 724.690 1492.635 724.705 ;
        RECT 1491.385 724.390 1492.635 724.690 ;
        RECT 1491.385 724.375 1491.715 724.390 ;
        RECT 1492.305 724.375 1492.635 724.390 ;
        RECT 1491.385 379.930 1491.715 379.945 ;
        RECT 1492.765 379.930 1493.095 379.945 ;
        RECT 1491.385 379.630 1493.095 379.930 ;
        RECT 1491.385 379.615 1491.715 379.630 ;
        RECT 1492.765 379.615 1493.095 379.630 ;
        RECT 674.425 37.890 674.755 37.905 ;
        RECT 1491.385 37.890 1491.715 37.905 ;
        RECT 674.425 37.590 1491.715 37.890 ;
        RECT 674.425 37.575 674.755 37.590 ;
        RECT 1491.385 37.575 1491.715 37.590 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1173.990 38.320 1174.310 38.380 ;
        RECT 1753.130 38.320 1753.450 38.380 ;
        RECT 1173.990 38.180 1753.450 38.320 ;
        RECT 1173.990 38.120 1174.310 38.180 ;
        RECT 1753.130 38.120 1753.450 38.180 ;
      LAYER via ;
        RECT 1174.020 38.120 1174.280 38.380 ;
        RECT 1753.160 38.120 1753.420 38.380 ;
      LAYER met2 ;
        RECT 1753.080 1700.000 1753.360 1704.000 ;
        RECT 1753.220 38.410 1753.360 1700.000 ;
        RECT 1174.020 38.090 1174.280 38.410 ;
        RECT 1753.160 38.090 1753.420 38.410 ;
        RECT 1174.080 2.400 1174.220 38.090 ;
        RECT 1173.870 -4.800 1174.430 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1191.930 35.260 1192.250 35.320 ;
        RECT 1759.570 35.260 1759.890 35.320 ;
        RECT 1191.930 35.120 1759.890 35.260 ;
        RECT 1191.930 35.060 1192.250 35.120 ;
        RECT 1759.570 35.060 1759.890 35.120 ;
      LAYER via ;
        RECT 1191.960 35.060 1192.220 35.320 ;
        RECT 1759.600 35.060 1759.860 35.320 ;
      LAYER met2 ;
        RECT 1762.280 1700.410 1762.560 1704.000 ;
        RECT 1759.660 1700.270 1762.560 1700.410 ;
        RECT 1759.660 35.350 1759.800 1700.270 ;
        RECT 1762.280 1700.000 1762.560 1700.270 ;
        RECT 1191.960 35.030 1192.220 35.350 ;
        RECT 1759.600 35.030 1759.860 35.350 ;
        RECT 1192.020 2.400 1192.160 35.030 ;
        RECT 1191.810 -4.800 1192.370 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1767.925 1207.425 1768.095 1255.875 ;
        RECT 1767.465 814.385 1767.635 903.975 ;
        RECT 1767.465 620.925 1767.635 669.375 ;
        RECT 1767.465 469.285 1767.635 517.395 ;
        RECT 1767.925 186.065 1768.095 227.715 ;
      LAYER mcon ;
        RECT 1767.925 1255.705 1768.095 1255.875 ;
        RECT 1767.465 903.805 1767.635 903.975 ;
        RECT 1767.465 669.205 1767.635 669.375 ;
        RECT 1767.465 517.225 1767.635 517.395 ;
        RECT 1767.925 227.545 1768.095 227.715 ;
      LAYER met1 ;
        RECT 1767.850 1642.440 1768.170 1642.500 ;
        RECT 1769.690 1642.440 1770.010 1642.500 ;
        RECT 1767.850 1642.300 1770.010 1642.440 ;
        RECT 1767.850 1642.240 1768.170 1642.300 ;
        RECT 1769.690 1642.240 1770.010 1642.300 ;
        RECT 1767.390 1545.880 1767.710 1545.940 ;
        RECT 1767.850 1545.880 1768.170 1545.940 ;
        RECT 1767.390 1545.740 1768.170 1545.880 ;
        RECT 1767.390 1545.680 1767.710 1545.740 ;
        RECT 1767.850 1545.680 1768.170 1545.740 ;
        RECT 1767.390 1497.740 1767.710 1498.000 ;
        RECT 1767.480 1496.980 1767.620 1497.740 ;
        RECT 1767.390 1496.720 1767.710 1496.980 ;
        RECT 1767.390 1490.460 1767.710 1490.520 ;
        RECT 1767.850 1490.460 1768.170 1490.520 ;
        RECT 1767.390 1490.320 1768.170 1490.460 ;
        RECT 1767.390 1490.260 1767.710 1490.320 ;
        RECT 1767.850 1490.260 1768.170 1490.320 ;
        RECT 1767.390 1400.700 1767.710 1400.760 ;
        RECT 1767.850 1400.700 1768.170 1400.760 ;
        RECT 1767.390 1400.560 1768.170 1400.700 ;
        RECT 1767.390 1400.500 1767.710 1400.560 ;
        RECT 1767.850 1400.500 1768.170 1400.560 ;
        RECT 1767.390 1317.880 1767.710 1318.140 ;
        RECT 1767.480 1317.400 1767.620 1317.880 ;
        RECT 1767.850 1317.400 1768.170 1317.460 ;
        RECT 1767.480 1317.260 1768.170 1317.400 ;
        RECT 1767.850 1317.200 1768.170 1317.260 ;
        RECT 1767.850 1255.860 1768.170 1255.920 ;
        RECT 1767.655 1255.720 1768.170 1255.860 ;
        RECT 1767.850 1255.660 1768.170 1255.720 ;
        RECT 1767.850 1207.580 1768.170 1207.640 ;
        RECT 1767.655 1207.440 1768.170 1207.580 ;
        RECT 1767.850 1207.380 1768.170 1207.440 ;
        RECT 1767.390 1152.840 1767.710 1152.900 ;
        RECT 1767.850 1152.840 1768.170 1152.900 ;
        RECT 1767.390 1152.700 1768.170 1152.840 ;
        RECT 1767.390 1152.640 1767.710 1152.700 ;
        RECT 1767.850 1152.640 1768.170 1152.700 ;
        RECT 1767.390 1124.760 1767.710 1125.020 ;
        RECT 1767.480 1124.280 1767.620 1124.760 ;
        RECT 1767.850 1124.280 1768.170 1124.340 ;
        RECT 1767.480 1124.140 1768.170 1124.280 ;
        RECT 1767.850 1124.080 1768.170 1124.140 ;
        RECT 1767.390 1062.740 1767.710 1062.800 ;
        RECT 1768.310 1062.740 1768.630 1062.800 ;
        RECT 1767.390 1062.600 1768.630 1062.740 ;
        RECT 1767.390 1062.540 1767.710 1062.600 ;
        RECT 1768.310 1062.540 1768.630 1062.600 ;
        RECT 1767.390 966.180 1767.710 966.240 ;
        RECT 1768.310 966.180 1768.630 966.240 ;
        RECT 1767.390 966.040 1768.630 966.180 ;
        RECT 1767.390 965.980 1767.710 966.040 ;
        RECT 1768.310 965.980 1768.630 966.040 ;
        RECT 1767.390 917.900 1767.710 917.960 ;
        RECT 1767.850 917.900 1768.170 917.960 ;
        RECT 1767.390 917.760 1768.170 917.900 ;
        RECT 1767.390 917.700 1767.710 917.760 ;
        RECT 1767.850 917.700 1768.170 917.760 ;
        RECT 1767.405 903.960 1767.695 904.005 ;
        RECT 1767.850 903.960 1768.170 904.020 ;
        RECT 1767.405 903.820 1768.170 903.960 ;
        RECT 1767.405 903.775 1767.695 903.820 ;
        RECT 1767.850 903.760 1768.170 903.820 ;
        RECT 1767.390 814.540 1767.710 814.600 ;
        RECT 1767.195 814.400 1767.710 814.540 ;
        RECT 1767.390 814.340 1767.710 814.400 ;
        RECT 1767.390 724.440 1767.710 724.500 ;
        RECT 1767.850 724.440 1768.170 724.500 ;
        RECT 1767.390 724.300 1768.170 724.440 ;
        RECT 1767.390 724.240 1767.710 724.300 ;
        RECT 1767.850 724.240 1768.170 724.300 ;
        RECT 1767.390 669.360 1767.710 669.420 ;
        RECT 1767.195 669.220 1767.710 669.360 ;
        RECT 1767.390 669.160 1767.710 669.220 ;
        RECT 1767.405 621.080 1767.695 621.125 ;
        RECT 1767.850 621.080 1768.170 621.140 ;
        RECT 1767.405 620.940 1768.170 621.080 ;
        RECT 1767.405 620.895 1767.695 620.940 ;
        RECT 1767.850 620.880 1768.170 620.940 ;
        RECT 1767.850 573.140 1768.170 573.200 ;
        RECT 1767.480 573.000 1768.170 573.140 ;
        RECT 1767.480 572.860 1767.620 573.000 ;
        RECT 1767.850 572.940 1768.170 573.000 ;
        RECT 1767.390 572.600 1767.710 572.860 ;
        RECT 1767.405 517.380 1767.695 517.425 ;
        RECT 1767.850 517.380 1768.170 517.440 ;
        RECT 1767.405 517.240 1768.170 517.380 ;
        RECT 1767.405 517.195 1767.695 517.240 ;
        RECT 1767.850 517.180 1768.170 517.240 ;
        RECT 1767.390 469.440 1767.710 469.500 ;
        RECT 1767.195 469.300 1767.710 469.440 ;
        RECT 1767.390 469.240 1767.710 469.300 ;
        RECT 1767.390 420.620 1767.710 420.880 ;
        RECT 1766.930 420.480 1767.250 420.540 ;
        RECT 1767.480 420.480 1767.620 420.620 ;
        RECT 1766.930 420.340 1767.620 420.480 ;
        RECT 1766.930 420.280 1767.250 420.340 ;
        RECT 1767.390 282.780 1767.710 282.840 ;
        RECT 1768.310 282.780 1768.630 282.840 ;
        RECT 1767.390 282.640 1768.630 282.780 ;
        RECT 1767.390 282.580 1767.710 282.640 ;
        RECT 1768.310 282.580 1768.630 282.640 ;
        RECT 1767.850 227.700 1768.170 227.760 ;
        RECT 1767.655 227.560 1768.170 227.700 ;
        RECT 1767.850 227.500 1768.170 227.560 ;
        RECT 1767.850 186.220 1768.170 186.280 ;
        RECT 1767.655 186.080 1768.170 186.220 ;
        RECT 1767.850 186.020 1768.170 186.080 ;
        RECT 1209.870 34.920 1210.190 34.980 ;
        RECT 1766.930 34.920 1767.250 34.980 ;
        RECT 1209.870 34.780 1767.250 34.920 ;
        RECT 1209.870 34.720 1210.190 34.780 ;
        RECT 1766.930 34.720 1767.250 34.780 ;
      LAYER via ;
        RECT 1767.880 1642.240 1768.140 1642.500 ;
        RECT 1769.720 1642.240 1769.980 1642.500 ;
        RECT 1767.420 1545.680 1767.680 1545.940 ;
        RECT 1767.880 1545.680 1768.140 1545.940 ;
        RECT 1767.420 1497.740 1767.680 1498.000 ;
        RECT 1767.420 1496.720 1767.680 1496.980 ;
        RECT 1767.420 1490.260 1767.680 1490.520 ;
        RECT 1767.880 1490.260 1768.140 1490.520 ;
        RECT 1767.420 1400.500 1767.680 1400.760 ;
        RECT 1767.880 1400.500 1768.140 1400.760 ;
        RECT 1767.420 1317.880 1767.680 1318.140 ;
        RECT 1767.880 1317.200 1768.140 1317.460 ;
        RECT 1767.880 1255.660 1768.140 1255.920 ;
        RECT 1767.880 1207.380 1768.140 1207.640 ;
        RECT 1767.420 1152.640 1767.680 1152.900 ;
        RECT 1767.880 1152.640 1768.140 1152.900 ;
        RECT 1767.420 1124.760 1767.680 1125.020 ;
        RECT 1767.880 1124.080 1768.140 1124.340 ;
        RECT 1767.420 1062.540 1767.680 1062.800 ;
        RECT 1768.340 1062.540 1768.600 1062.800 ;
        RECT 1767.420 965.980 1767.680 966.240 ;
        RECT 1768.340 965.980 1768.600 966.240 ;
        RECT 1767.420 917.700 1767.680 917.960 ;
        RECT 1767.880 917.700 1768.140 917.960 ;
        RECT 1767.880 903.760 1768.140 904.020 ;
        RECT 1767.420 814.340 1767.680 814.600 ;
        RECT 1767.420 724.240 1767.680 724.500 ;
        RECT 1767.880 724.240 1768.140 724.500 ;
        RECT 1767.420 669.160 1767.680 669.420 ;
        RECT 1767.880 620.880 1768.140 621.140 ;
        RECT 1767.880 572.940 1768.140 573.200 ;
        RECT 1767.420 572.600 1767.680 572.860 ;
        RECT 1767.880 517.180 1768.140 517.440 ;
        RECT 1767.420 469.240 1767.680 469.500 ;
        RECT 1767.420 420.620 1767.680 420.880 ;
        RECT 1766.960 420.280 1767.220 420.540 ;
        RECT 1767.420 282.580 1767.680 282.840 ;
        RECT 1768.340 282.580 1768.600 282.840 ;
        RECT 1767.880 227.500 1768.140 227.760 ;
        RECT 1767.880 186.020 1768.140 186.280 ;
        RECT 1209.900 34.720 1210.160 34.980 ;
        RECT 1766.960 34.720 1767.220 34.980 ;
      LAYER met2 ;
        RECT 1771.020 1700.410 1771.300 1704.000 ;
        RECT 1769.780 1700.270 1771.300 1700.410 ;
        RECT 1769.780 1642.530 1769.920 1700.270 ;
        RECT 1771.020 1700.000 1771.300 1700.270 ;
        RECT 1767.880 1642.210 1768.140 1642.530 ;
        RECT 1769.720 1642.210 1769.980 1642.530 ;
        RECT 1767.940 1545.970 1768.080 1642.210 ;
        RECT 1767.420 1545.650 1767.680 1545.970 ;
        RECT 1767.880 1545.650 1768.140 1545.970 ;
        RECT 1767.480 1498.030 1767.620 1545.650 ;
        RECT 1767.420 1497.710 1767.680 1498.030 ;
        RECT 1767.420 1496.690 1767.680 1497.010 ;
        RECT 1767.480 1490.550 1767.620 1496.690 ;
        RECT 1767.420 1490.230 1767.680 1490.550 ;
        RECT 1767.880 1490.230 1768.140 1490.550 ;
        RECT 1767.940 1400.790 1768.080 1490.230 ;
        RECT 1767.420 1400.470 1767.680 1400.790 ;
        RECT 1767.880 1400.470 1768.140 1400.790 ;
        RECT 1767.480 1318.170 1767.620 1400.470 ;
        RECT 1767.420 1317.850 1767.680 1318.170 ;
        RECT 1767.880 1317.170 1768.140 1317.490 ;
        RECT 1767.940 1255.950 1768.080 1317.170 ;
        RECT 1767.880 1255.630 1768.140 1255.950 ;
        RECT 1767.880 1207.350 1768.140 1207.670 ;
        RECT 1767.940 1152.930 1768.080 1207.350 ;
        RECT 1767.420 1152.610 1767.680 1152.930 ;
        RECT 1767.880 1152.610 1768.140 1152.930 ;
        RECT 1767.480 1125.050 1767.620 1152.610 ;
        RECT 1767.420 1124.730 1767.680 1125.050 ;
        RECT 1767.880 1124.050 1768.140 1124.370 ;
        RECT 1767.940 1087.050 1768.080 1124.050 ;
        RECT 1767.940 1086.910 1768.540 1087.050 ;
        RECT 1768.400 1062.830 1768.540 1086.910 ;
        RECT 1767.420 1062.570 1767.680 1062.830 ;
        RECT 1767.420 1062.510 1768.080 1062.570 ;
        RECT 1768.340 1062.510 1768.600 1062.830 ;
        RECT 1767.480 1062.430 1768.080 1062.510 ;
        RECT 1767.940 990.490 1768.080 1062.430 ;
        RECT 1767.940 990.350 1768.540 990.490 ;
        RECT 1768.400 966.270 1768.540 990.350 ;
        RECT 1767.420 965.950 1767.680 966.270 ;
        RECT 1768.340 965.950 1768.600 966.270 ;
        RECT 1767.480 917.990 1767.620 965.950 ;
        RECT 1767.420 917.670 1767.680 917.990 ;
        RECT 1767.880 917.670 1768.140 917.990 ;
        RECT 1767.940 904.050 1768.080 917.670 ;
        RECT 1767.880 903.730 1768.140 904.050 ;
        RECT 1767.420 814.310 1767.680 814.630 ;
        RECT 1767.480 766.090 1767.620 814.310 ;
        RECT 1767.480 765.950 1768.080 766.090 ;
        RECT 1767.940 724.530 1768.080 765.950 ;
        RECT 1767.420 724.210 1767.680 724.530 ;
        RECT 1767.880 724.210 1768.140 724.530 ;
        RECT 1767.480 670.325 1767.620 724.210 ;
        RECT 1767.410 669.955 1767.690 670.325 ;
        RECT 1767.410 669.275 1767.690 669.645 ;
        RECT 1767.420 669.130 1767.680 669.275 ;
        RECT 1767.880 620.850 1768.140 621.170 ;
        RECT 1767.940 573.230 1768.080 620.850 ;
        RECT 1767.880 572.910 1768.140 573.230 ;
        RECT 1767.420 572.570 1767.680 572.890 ;
        RECT 1767.480 572.405 1767.620 572.570 ;
        RECT 1767.410 572.035 1767.690 572.405 ;
        RECT 1767.870 571.355 1768.150 571.725 ;
        RECT 1767.940 517.470 1768.080 571.355 ;
        RECT 1767.880 517.150 1768.140 517.470 ;
        RECT 1767.420 469.210 1767.680 469.530 ;
        RECT 1767.480 420.910 1767.620 469.210 ;
        RECT 1767.420 420.590 1767.680 420.910 ;
        RECT 1766.960 420.250 1767.220 420.570 ;
        RECT 1767.020 331.685 1767.160 420.250 ;
        RECT 1766.950 331.315 1767.230 331.685 ;
        RECT 1768.330 329.955 1768.610 330.325 ;
        RECT 1768.400 282.870 1768.540 329.955 ;
        RECT 1767.420 282.550 1767.680 282.870 ;
        RECT 1768.340 282.550 1768.600 282.870 ;
        RECT 1767.480 235.010 1767.620 282.550 ;
        RECT 1767.480 234.870 1768.080 235.010 ;
        RECT 1767.940 227.790 1768.080 234.870 ;
        RECT 1767.880 227.470 1768.140 227.790 ;
        RECT 1767.880 185.990 1768.140 186.310 ;
        RECT 1767.940 162.250 1768.080 185.990 ;
        RECT 1767.940 162.110 1768.540 162.250 ;
        RECT 1768.400 60.930 1768.540 162.110 ;
        RECT 1767.020 60.790 1768.540 60.930 ;
        RECT 1767.020 35.010 1767.160 60.790 ;
        RECT 1209.900 34.690 1210.160 35.010 ;
        RECT 1766.960 34.690 1767.220 35.010 ;
        RECT 1209.960 2.400 1210.100 34.690 ;
        RECT 1209.750 -4.800 1210.310 2.400 ;
      LAYER via2 ;
        RECT 1767.410 670.000 1767.690 670.280 ;
        RECT 1767.410 669.320 1767.690 669.600 ;
        RECT 1767.410 572.080 1767.690 572.360 ;
        RECT 1767.870 571.400 1768.150 571.680 ;
        RECT 1766.950 331.360 1767.230 331.640 ;
        RECT 1768.330 330.000 1768.610 330.280 ;
      LAYER met3 ;
        RECT 1767.385 670.290 1767.715 670.305 ;
        RECT 1767.385 669.975 1767.930 670.290 ;
        RECT 1767.630 669.625 1767.930 669.975 ;
        RECT 1767.385 669.310 1767.930 669.625 ;
        RECT 1767.385 669.295 1767.715 669.310 ;
        RECT 1767.385 572.370 1767.715 572.385 ;
        RECT 1766.710 572.070 1767.715 572.370 ;
        RECT 1766.710 571.690 1767.010 572.070 ;
        RECT 1767.385 572.055 1767.715 572.070 ;
        RECT 1767.845 571.690 1768.175 571.705 ;
        RECT 1766.710 571.390 1768.175 571.690 ;
        RECT 1767.845 571.375 1768.175 571.390 ;
        RECT 1766.925 331.650 1767.255 331.665 ;
        RECT 1766.925 331.350 1767.930 331.650 ;
        RECT 1766.925 331.335 1767.255 331.350 ;
        RECT 1767.630 330.290 1767.930 331.350 ;
        RECT 1768.305 330.290 1768.635 330.305 ;
        RECT 1767.630 329.990 1768.635 330.290 ;
        RECT 1768.305 329.975 1768.635 329.990 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1227.810 38.660 1228.130 38.720 ;
        RECT 1780.730 38.660 1781.050 38.720 ;
        RECT 1227.810 38.520 1781.050 38.660 ;
        RECT 1227.810 38.460 1228.130 38.520 ;
        RECT 1780.730 38.460 1781.050 38.520 ;
      LAYER via ;
        RECT 1227.840 38.460 1228.100 38.720 ;
        RECT 1780.760 38.460 1781.020 38.720 ;
      LAYER met2 ;
        RECT 1780.220 1700.410 1780.500 1704.000 ;
        RECT 1780.220 1700.270 1780.960 1700.410 ;
        RECT 1780.220 1700.000 1780.500 1700.270 ;
        RECT 1780.820 38.750 1780.960 1700.270 ;
        RECT 1227.840 38.430 1228.100 38.750 ;
        RECT 1780.760 38.430 1781.020 38.750 ;
        RECT 1227.900 2.400 1228.040 38.430 ;
        RECT 1227.690 -4.800 1228.250 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1245.750 39.000 1246.070 39.060 ;
        RECT 1787.170 39.000 1787.490 39.060 ;
        RECT 1245.750 38.860 1787.490 39.000 ;
        RECT 1245.750 38.800 1246.070 38.860 ;
        RECT 1787.170 38.800 1787.490 38.860 ;
      LAYER via ;
        RECT 1245.780 38.800 1246.040 39.060 ;
        RECT 1787.200 38.800 1787.460 39.060 ;
      LAYER met2 ;
        RECT 1789.420 1700.410 1789.700 1704.000 ;
        RECT 1787.260 1700.270 1789.700 1700.410 ;
        RECT 1787.260 39.090 1787.400 1700.270 ;
        RECT 1789.420 1700.000 1789.700 1700.270 ;
        RECT 1245.780 38.770 1246.040 39.090 ;
        RECT 1787.200 38.770 1787.460 39.090 ;
        RECT 1245.840 2.400 1245.980 38.770 ;
        RECT 1245.630 -4.800 1246.190 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1795.985 938.485 1796.155 986.595 ;
        RECT 1795.065 389.725 1795.235 420.835 ;
        RECT 1795.985 269.025 1796.155 317.475 ;
        RECT 1795.525 227.885 1795.695 241.995 ;
      LAYER mcon ;
        RECT 1795.985 986.425 1796.155 986.595 ;
        RECT 1795.065 420.665 1795.235 420.835 ;
        RECT 1795.985 317.305 1796.155 317.475 ;
        RECT 1795.525 241.825 1795.695 241.995 ;
      LAYER met1 ;
        RECT 1795.450 1642.440 1795.770 1642.500 ;
        RECT 1797.290 1642.440 1797.610 1642.500 ;
        RECT 1795.450 1642.300 1797.610 1642.440 ;
        RECT 1795.450 1642.240 1795.770 1642.300 ;
        RECT 1797.290 1642.240 1797.610 1642.300 ;
        RECT 1795.450 1608.100 1795.770 1608.160 ;
        RECT 1795.080 1607.960 1795.770 1608.100 ;
        RECT 1795.080 1607.820 1795.220 1607.960 ;
        RECT 1795.450 1607.900 1795.770 1607.960 ;
        RECT 1794.990 1607.560 1795.310 1607.820 ;
        RECT 1794.990 1400.700 1795.310 1400.760 ;
        RECT 1795.450 1400.700 1795.770 1400.760 ;
        RECT 1794.990 1400.560 1795.770 1400.700 ;
        RECT 1794.990 1400.500 1795.310 1400.560 ;
        RECT 1795.450 1400.500 1795.770 1400.560 ;
        RECT 1795.450 1304.480 1795.770 1304.540 ;
        RECT 1795.910 1304.480 1796.230 1304.540 ;
        RECT 1795.450 1304.340 1796.230 1304.480 ;
        RECT 1795.450 1304.280 1795.770 1304.340 ;
        RECT 1795.910 1304.280 1796.230 1304.340 ;
        RECT 1795.450 1249.740 1795.770 1249.800 ;
        RECT 1795.080 1249.600 1795.770 1249.740 ;
        RECT 1795.080 1249.460 1795.220 1249.600 ;
        RECT 1795.450 1249.540 1795.770 1249.600 ;
        RECT 1794.990 1249.200 1795.310 1249.460 ;
        RECT 1795.450 1200.780 1795.770 1200.840 ;
        RECT 1796.370 1200.780 1796.690 1200.840 ;
        RECT 1795.450 1200.640 1796.690 1200.780 ;
        RECT 1795.450 1200.580 1795.770 1200.640 ;
        RECT 1796.370 1200.580 1796.690 1200.640 ;
        RECT 1795.450 1169.500 1795.770 1169.560 ;
        RECT 1796.370 1169.500 1796.690 1169.560 ;
        RECT 1795.450 1169.360 1796.690 1169.500 ;
        RECT 1795.450 1169.300 1795.770 1169.360 ;
        RECT 1796.370 1169.300 1796.690 1169.360 ;
        RECT 1794.530 1104.220 1794.850 1104.280 ;
        RECT 1795.450 1104.220 1795.770 1104.280 ;
        RECT 1794.530 1104.080 1795.770 1104.220 ;
        RECT 1794.530 1104.020 1794.850 1104.080 ;
        RECT 1795.450 1104.020 1795.770 1104.080 ;
        RECT 1794.530 1089.940 1794.850 1090.000 ;
        RECT 1794.990 1089.940 1795.310 1090.000 ;
        RECT 1794.530 1089.800 1795.310 1089.940 ;
        RECT 1794.530 1089.740 1794.850 1089.800 ;
        RECT 1794.990 1089.740 1795.310 1089.800 ;
        RECT 1795.450 986.580 1795.770 986.640 ;
        RECT 1795.925 986.580 1796.215 986.625 ;
        RECT 1795.450 986.440 1796.215 986.580 ;
        RECT 1795.450 986.380 1795.770 986.440 ;
        RECT 1795.925 986.395 1796.215 986.440 ;
        RECT 1795.450 938.640 1795.770 938.700 ;
        RECT 1795.925 938.640 1796.215 938.685 ;
        RECT 1795.450 938.500 1796.215 938.640 ;
        RECT 1795.450 938.440 1795.770 938.500 ;
        RECT 1795.925 938.455 1796.215 938.500 ;
        RECT 1795.450 896.480 1795.770 896.540 ;
        RECT 1795.910 896.480 1796.230 896.540 ;
        RECT 1795.450 896.340 1796.230 896.480 ;
        RECT 1795.450 896.280 1795.770 896.340 ;
        RECT 1795.910 896.280 1796.230 896.340 ;
        RECT 1794.990 724.440 1795.310 724.500 ;
        RECT 1795.910 724.440 1796.230 724.500 ;
        RECT 1794.990 724.300 1796.230 724.440 ;
        RECT 1794.990 724.240 1795.310 724.300 ;
        RECT 1795.910 724.240 1796.230 724.300 ;
        RECT 1794.990 448.360 1795.310 448.420 ;
        RECT 1795.910 448.360 1796.230 448.420 ;
        RECT 1794.990 448.220 1796.230 448.360 ;
        RECT 1794.990 448.160 1795.310 448.220 ;
        RECT 1795.910 448.160 1796.230 448.220 ;
        RECT 1794.990 420.820 1795.310 420.880 ;
        RECT 1794.795 420.680 1795.310 420.820 ;
        RECT 1794.990 420.620 1795.310 420.680 ;
        RECT 1795.005 389.880 1795.295 389.925 ;
        RECT 1796.370 389.880 1796.690 389.940 ;
        RECT 1795.005 389.740 1796.690 389.880 ;
        RECT 1795.005 389.695 1795.295 389.740 ;
        RECT 1796.370 389.680 1796.690 389.740 ;
        RECT 1795.910 365.740 1796.230 365.800 ;
        RECT 1796.370 365.740 1796.690 365.800 ;
        RECT 1795.910 365.600 1796.690 365.740 ;
        RECT 1795.910 365.540 1796.230 365.600 ;
        RECT 1796.370 365.540 1796.690 365.600 ;
        RECT 1795.910 317.460 1796.230 317.520 ;
        RECT 1795.715 317.320 1796.230 317.460 ;
        RECT 1795.910 317.260 1796.230 317.320 ;
        RECT 1795.910 269.180 1796.230 269.240 ;
        RECT 1795.715 269.040 1796.230 269.180 ;
        RECT 1795.910 268.980 1796.230 269.040 ;
        RECT 1795.465 241.980 1795.755 242.025 ;
        RECT 1795.910 241.980 1796.230 242.040 ;
        RECT 1795.465 241.840 1796.230 241.980 ;
        RECT 1795.465 241.795 1795.755 241.840 ;
        RECT 1795.910 241.780 1796.230 241.840 ;
        RECT 1795.450 228.040 1795.770 228.100 ;
        RECT 1795.255 227.900 1795.770 228.040 ;
        RECT 1795.450 227.840 1795.770 227.900 ;
        RECT 1794.530 179.420 1794.850 179.480 ;
        RECT 1795.450 179.420 1795.770 179.480 ;
        RECT 1794.530 179.280 1795.770 179.420 ;
        RECT 1794.530 179.220 1794.850 179.280 ;
        RECT 1795.450 179.220 1795.770 179.280 ;
        RECT 1794.530 130.940 1794.850 131.200 ;
        RECT 1794.620 130.800 1794.760 130.940 ;
        RECT 1794.990 130.800 1795.310 130.860 ;
        RECT 1794.620 130.660 1795.310 130.800 ;
        RECT 1794.990 130.600 1795.310 130.660 ;
        RECT 1794.530 41.720 1794.850 41.780 ;
        RECT 1794.990 41.720 1795.310 41.780 ;
        RECT 1794.530 41.580 1795.310 41.720 ;
        RECT 1794.530 41.520 1794.850 41.580 ;
        RECT 1794.990 41.520 1795.310 41.580 ;
        RECT 1263.230 39.340 1263.550 39.400 ;
        RECT 1794.530 39.340 1794.850 39.400 ;
        RECT 1263.230 39.200 1794.850 39.340 ;
        RECT 1263.230 39.140 1263.550 39.200 ;
        RECT 1794.530 39.140 1794.850 39.200 ;
      LAYER via ;
        RECT 1795.480 1642.240 1795.740 1642.500 ;
        RECT 1797.320 1642.240 1797.580 1642.500 ;
        RECT 1795.480 1607.900 1795.740 1608.160 ;
        RECT 1795.020 1607.560 1795.280 1607.820 ;
        RECT 1795.020 1400.500 1795.280 1400.760 ;
        RECT 1795.480 1400.500 1795.740 1400.760 ;
        RECT 1795.480 1304.280 1795.740 1304.540 ;
        RECT 1795.940 1304.280 1796.200 1304.540 ;
        RECT 1795.480 1249.540 1795.740 1249.800 ;
        RECT 1795.020 1249.200 1795.280 1249.460 ;
        RECT 1795.480 1200.580 1795.740 1200.840 ;
        RECT 1796.400 1200.580 1796.660 1200.840 ;
        RECT 1795.480 1169.300 1795.740 1169.560 ;
        RECT 1796.400 1169.300 1796.660 1169.560 ;
        RECT 1794.560 1104.020 1794.820 1104.280 ;
        RECT 1795.480 1104.020 1795.740 1104.280 ;
        RECT 1794.560 1089.740 1794.820 1090.000 ;
        RECT 1795.020 1089.740 1795.280 1090.000 ;
        RECT 1795.480 986.380 1795.740 986.640 ;
        RECT 1795.480 938.440 1795.740 938.700 ;
        RECT 1795.480 896.280 1795.740 896.540 ;
        RECT 1795.940 896.280 1796.200 896.540 ;
        RECT 1795.020 724.240 1795.280 724.500 ;
        RECT 1795.940 724.240 1796.200 724.500 ;
        RECT 1795.020 448.160 1795.280 448.420 ;
        RECT 1795.940 448.160 1796.200 448.420 ;
        RECT 1795.020 420.620 1795.280 420.880 ;
        RECT 1796.400 389.680 1796.660 389.940 ;
        RECT 1795.940 365.540 1796.200 365.800 ;
        RECT 1796.400 365.540 1796.660 365.800 ;
        RECT 1795.940 317.260 1796.200 317.520 ;
        RECT 1795.940 268.980 1796.200 269.240 ;
        RECT 1795.940 241.780 1796.200 242.040 ;
        RECT 1795.480 227.840 1795.740 228.100 ;
        RECT 1794.560 179.220 1794.820 179.480 ;
        RECT 1795.480 179.220 1795.740 179.480 ;
        RECT 1794.560 130.940 1794.820 131.200 ;
        RECT 1795.020 130.600 1795.280 130.860 ;
        RECT 1794.560 41.520 1794.820 41.780 ;
        RECT 1795.020 41.520 1795.280 41.780 ;
        RECT 1263.260 39.140 1263.520 39.400 ;
        RECT 1794.560 39.140 1794.820 39.400 ;
      LAYER met2 ;
        RECT 1798.620 1700.410 1798.900 1704.000 ;
        RECT 1797.380 1700.270 1798.900 1700.410 ;
        RECT 1797.380 1642.530 1797.520 1700.270 ;
        RECT 1798.620 1700.000 1798.900 1700.270 ;
        RECT 1795.480 1642.210 1795.740 1642.530 ;
        RECT 1797.320 1642.210 1797.580 1642.530 ;
        RECT 1795.540 1608.190 1795.680 1642.210 ;
        RECT 1795.480 1607.870 1795.740 1608.190 ;
        RECT 1795.020 1607.530 1795.280 1607.850 ;
        RECT 1795.080 1593.650 1795.220 1607.530 ;
        RECT 1795.080 1593.510 1795.680 1593.650 ;
        RECT 1795.540 1463.090 1795.680 1593.510 ;
        RECT 1795.080 1462.950 1795.680 1463.090 ;
        RECT 1795.080 1414.130 1795.220 1462.950 ;
        RECT 1795.080 1413.990 1795.680 1414.130 ;
        RECT 1795.540 1400.790 1795.680 1413.990 ;
        RECT 1795.020 1400.470 1795.280 1400.790 ;
        RECT 1795.480 1400.470 1795.740 1400.790 ;
        RECT 1795.080 1353.725 1795.220 1400.470 ;
        RECT 1795.010 1353.355 1795.290 1353.725 ;
        RECT 1795.930 1351.995 1796.210 1352.365 ;
        RECT 1796.000 1304.570 1796.140 1351.995 ;
        RECT 1795.480 1304.250 1795.740 1304.570 ;
        RECT 1795.940 1304.250 1796.200 1304.570 ;
        RECT 1795.540 1249.830 1795.680 1304.250 ;
        RECT 1795.480 1249.510 1795.740 1249.830 ;
        RECT 1795.020 1249.170 1795.280 1249.490 ;
        RECT 1795.080 1249.005 1795.220 1249.170 ;
        RECT 1795.010 1248.635 1795.290 1249.005 ;
        RECT 1796.390 1248.635 1796.670 1249.005 ;
        RECT 1796.460 1200.870 1796.600 1248.635 ;
        RECT 1795.480 1200.550 1795.740 1200.870 ;
        RECT 1796.400 1200.550 1796.660 1200.870 ;
        RECT 1795.540 1169.590 1795.680 1200.550 ;
        RECT 1795.480 1169.270 1795.740 1169.590 ;
        RECT 1796.400 1169.270 1796.660 1169.590 ;
        RECT 1796.460 1145.645 1796.600 1169.270 ;
        RECT 1795.470 1145.275 1795.750 1145.645 ;
        RECT 1796.390 1145.275 1796.670 1145.645 ;
        RECT 1795.540 1104.310 1795.680 1145.275 ;
        RECT 1794.560 1103.990 1794.820 1104.310 ;
        RECT 1795.480 1103.990 1795.740 1104.310 ;
        RECT 1794.620 1090.030 1794.760 1103.990 ;
        RECT 1794.560 1089.710 1794.820 1090.030 ;
        RECT 1795.020 1089.710 1795.280 1090.030 ;
        RECT 1795.080 1048.290 1795.220 1089.710 ;
        RECT 1795.080 1048.150 1796.140 1048.290 ;
        RECT 1796.000 1001.485 1796.140 1048.150 ;
        RECT 1795.930 1001.115 1796.210 1001.485 ;
        RECT 1795.470 993.635 1795.750 994.005 ;
        RECT 1795.540 986.670 1795.680 993.635 ;
        RECT 1795.480 986.350 1795.740 986.670 ;
        RECT 1795.480 938.410 1795.740 938.730 ;
        RECT 1795.540 896.570 1795.680 938.410 ;
        RECT 1795.480 896.250 1795.740 896.570 ;
        RECT 1795.940 896.250 1796.200 896.570 ;
        RECT 1796.000 724.725 1796.140 896.250 ;
        RECT 1795.010 724.355 1795.290 724.725 ;
        RECT 1795.930 724.355 1796.210 724.725 ;
        RECT 1795.020 724.210 1795.280 724.355 ;
        RECT 1795.940 724.210 1796.200 724.355 ;
        RECT 1796.000 699.450 1796.140 724.210 ;
        RECT 1795.540 699.310 1796.140 699.450 ;
        RECT 1795.540 621.365 1795.680 699.310 ;
        RECT 1795.470 620.995 1795.750 621.365 ;
        RECT 1795.930 572.035 1796.210 572.405 ;
        RECT 1796.000 448.450 1796.140 572.035 ;
        RECT 1795.020 448.130 1795.280 448.450 ;
        RECT 1795.940 448.130 1796.200 448.450 ;
        RECT 1795.080 420.910 1795.220 448.130 ;
        RECT 1795.020 420.590 1795.280 420.910 ;
        RECT 1796.400 389.650 1796.660 389.970 ;
        RECT 1796.460 365.830 1796.600 389.650 ;
        RECT 1795.940 365.510 1796.200 365.830 ;
        RECT 1796.400 365.510 1796.660 365.830 ;
        RECT 1796.000 317.550 1796.140 365.510 ;
        RECT 1795.940 317.230 1796.200 317.550 ;
        RECT 1795.940 268.950 1796.200 269.270 ;
        RECT 1796.000 242.070 1796.140 268.950 ;
        RECT 1795.940 241.750 1796.200 242.070 ;
        RECT 1795.480 227.810 1795.740 228.130 ;
        RECT 1795.540 179.510 1795.680 227.810 ;
        RECT 1794.560 179.190 1794.820 179.510 ;
        RECT 1795.480 179.190 1795.740 179.510 ;
        RECT 1794.620 131.230 1794.760 179.190 ;
        RECT 1794.560 130.910 1794.820 131.230 ;
        RECT 1795.020 130.570 1795.280 130.890 ;
        RECT 1795.080 41.810 1795.220 130.570 ;
        RECT 1794.560 41.490 1794.820 41.810 ;
        RECT 1795.020 41.490 1795.280 41.810 ;
        RECT 1794.620 39.430 1794.760 41.490 ;
        RECT 1263.260 39.110 1263.520 39.430 ;
        RECT 1794.560 39.110 1794.820 39.430 ;
        RECT 1263.320 2.400 1263.460 39.110 ;
        RECT 1263.110 -4.800 1263.670 2.400 ;
      LAYER via2 ;
        RECT 1795.010 1353.400 1795.290 1353.680 ;
        RECT 1795.930 1352.040 1796.210 1352.320 ;
        RECT 1795.010 1248.680 1795.290 1248.960 ;
        RECT 1796.390 1248.680 1796.670 1248.960 ;
        RECT 1795.470 1145.320 1795.750 1145.600 ;
        RECT 1796.390 1145.320 1796.670 1145.600 ;
        RECT 1795.930 1001.160 1796.210 1001.440 ;
        RECT 1795.470 993.680 1795.750 993.960 ;
        RECT 1795.010 724.400 1795.290 724.680 ;
        RECT 1795.930 724.400 1796.210 724.680 ;
        RECT 1795.470 621.040 1795.750 621.320 ;
        RECT 1795.930 572.080 1796.210 572.360 ;
      LAYER met3 ;
        RECT 1794.985 1353.690 1795.315 1353.705 ;
        RECT 1794.310 1353.390 1795.315 1353.690 ;
        RECT 1794.310 1352.330 1794.610 1353.390 ;
        RECT 1794.985 1353.375 1795.315 1353.390 ;
        RECT 1795.905 1352.330 1796.235 1352.345 ;
        RECT 1794.310 1352.030 1796.235 1352.330 ;
        RECT 1795.905 1352.015 1796.235 1352.030 ;
        RECT 1794.985 1248.970 1795.315 1248.985 ;
        RECT 1796.365 1248.970 1796.695 1248.985 ;
        RECT 1794.985 1248.670 1796.695 1248.970 ;
        RECT 1794.985 1248.655 1795.315 1248.670 ;
        RECT 1796.365 1248.655 1796.695 1248.670 ;
        RECT 1795.445 1145.610 1795.775 1145.625 ;
        RECT 1796.365 1145.610 1796.695 1145.625 ;
        RECT 1795.445 1145.310 1796.695 1145.610 ;
        RECT 1795.445 1145.295 1795.775 1145.310 ;
        RECT 1796.365 1145.295 1796.695 1145.310 ;
        RECT 1795.190 1001.450 1795.570 1001.460 ;
        RECT 1795.905 1001.450 1796.235 1001.465 ;
        RECT 1795.190 1001.150 1796.235 1001.450 ;
        RECT 1795.190 1001.140 1795.570 1001.150 ;
        RECT 1795.905 1001.135 1796.235 1001.150 ;
        RECT 1795.445 993.980 1795.775 993.985 ;
        RECT 1795.190 993.970 1795.775 993.980 ;
        RECT 1795.190 993.670 1796.000 993.970 ;
        RECT 1795.190 993.660 1795.775 993.670 ;
        RECT 1795.445 993.655 1795.775 993.660 ;
        RECT 1794.985 724.690 1795.315 724.705 ;
        RECT 1795.905 724.690 1796.235 724.705 ;
        RECT 1794.985 724.390 1796.235 724.690 ;
        RECT 1794.985 724.375 1795.315 724.390 ;
        RECT 1795.905 724.375 1796.235 724.390 ;
        RECT 1795.445 621.330 1795.775 621.345 ;
        RECT 1795.230 621.015 1795.775 621.330 ;
        RECT 1795.230 620.660 1795.530 621.015 ;
        RECT 1795.190 620.340 1795.570 620.660 ;
        RECT 1795.190 572.740 1795.570 573.060 ;
        RECT 1795.230 572.370 1795.530 572.740 ;
        RECT 1795.905 572.370 1796.235 572.385 ;
        RECT 1795.230 572.070 1796.235 572.370 ;
        RECT 1795.905 572.055 1796.235 572.070 ;
      LAYER via3 ;
        RECT 1795.220 1001.140 1795.540 1001.460 ;
        RECT 1795.220 993.660 1795.540 993.980 ;
        RECT 1795.220 620.340 1795.540 620.660 ;
        RECT 1795.220 572.740 1795.540 573.060 ;
      LAYER met4 ;
        RECT 1795.215 1001.135 1795.545 1001.465 ;
        RECT 1795.230 993.985 1795.530 1001.135 ;
        RECT 1795.215 993.655 1795.545 993.985 ;
        RECT 1795.215 620.335 1795.545 620.665 ;
        RECT 1795.230 573.065 1795.530 620.335 ;
        RECT 1795.215 572.735 1795.545 573.065 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1281.170 39.680 1281.490 39.740 ;
        RECT 1807.870 39.680 1808.190 39.740 ;
        RECT 1281.170 39.540 1808.190 39.680 ;
        RECT 1281.170 39.480 1281.490 39.540 ;
        RECT 1807.870 39.480 1808.190 39.540 ;
      LAYER via ;
        RECT 1281.200 39.480 1281.460 39.740 ;
        RECT 1807.900 39.480 1808.160 39.740 ;
      LAYER met2 ;
        RECT 1807.820 1700.000 1808.100 1704.000 ;
        RECT 1807.960 39.770 1808.100 1700.000 ;
        RECT 1281.200 39.450 1281.460 39.770 ;
        RECT 1807.900 39.450 1808.160 39.770 ;
        RECT 1281.260 2.400 1281.400 39.450 ;
        RECT 1281.050 -4.800 1281.610 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1299.110 40.020 1299.430 40.080 ;
        RECT 1815.230 40.020 1815.550 40.080 ;
        RECT 1299.110 39.880 1815.550 40.020 ;
        RECT 1299.110 39.820 1299.430 39.880 ;
        RECT 1815.230 39.820 1815.550 39.880 ;
      LAYER via ;
        RECT 1299.140 39.820 1299.400 40.080 ;
        RECT 1815.260 39.820 1815.520 40.080 ;
      LAYER met2 ;
        RECT 1817.020 1700.410 1817.300 1704.000 ;
        RECT 1815.320 1700.270 1817.300 1700.410 ;
        RECT 1815.320 40.110 1815.460 1700.270 ;
        RECT 1817.020 1700.000 1817.300 1700.270 ;
        RECT 1299.140 39.790 1299.400 40.110 ;
        RECT 1815.260 39.790 1815.520 40.110 ;
        RECT 1299.200 2.400 1299.340 39.790 ;
        RECT 1298.990 -4.800 1299.550 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1822.665 1490.645 1822.835 1538.755 ;
        RECT 1822.665 1424.685 1822.835 1456.815 ;
        RECT 1820.825 1041.845 1820.995 1062.755 ;
        RECT 1822.665 931.345 1822.835 952.255 ;
        RECT 1822.665 421.005 1822.835 469.115 ;
        RECT 1822.665 324.445 1822.835 372.555 ;
        RECT 1824.045 87.125 1824.215 131.155 ;
      LAYER mcon ;
        RECT 1822.665 1538.585 1822.835 1538.755 ;
        RECT 1822.665 1456.645 1822.835 1456.815 ;
        RECT 1820.825 1062.585 1820.995 1062.755 ;
        RECT 1822.665 952.085 1822.835 952.255 ;
        RECT 1822.665 468.945 1822.835 469.115 ;
        RECT 1822.665 372.385 1822.835 372.555 ;
        RECT 1824.045 130.985 1824.215 131.155 ;
      LAYER met1 ;
        RECT 1823.050 1642.440 1823.370 1642.500 ;
        RECT 1823.970 1642.440 1824.290 1642.500 ;
        RECT 1823.050 1642.300 1824.290 1642.440 ;
        RECT 1823.050 1642.240 1823.370 1642.300 ;
        RECT 1823.970 1642.240 1824.290 1642.300 ;
        RECT 1822.590 1545.880 1822.910 1545.940 ;
        RECT 1823.050 1545.880 1823.370 1545.940 ;
        RECT 1822.590 1545.740 1823.370 1545.880 ;
        RECT 1822.590 1545.680 1822.910 1545.740 ;
        RECT 1823.050 1545.680 1823.370 1545.740 ;
        RECT 1822.590 1538.740 1822.910 1538.800 ;
        RECT 1822.395 1538.600 1822.910 1538.740 ;
        RECT 1822.590 1538.540 1822.910 1538.600 ;
        RECT 1822.605 1490.800 1822.895 1490.845 ;
        RECT 1823.050 1490.800 1823.370 1490.860 ;
        RECT 1822.605 1490.660 1823.370 1490.800 ;
        RECT 1822.605 1490.615 1822.895 1490.660 ;
        RECT 1823.050 1490.600 1823.370 1490.660 ;
        RECT 1822.590 1456.800 1822.910 1456.860 ;
        RECT 1822.395 1456.660 1822.910 1456.800 ;
        RECT 1822.590 1456.600 1822.910 1456.660 ;
        RECT 1822.605 1424.840 1822.895 1424.885 ;
        RECT 1823.050 1424.840 1823.370 1424.900 ;
        RECT 1822.605 1424.700 1823.370 1424.840 ;
        RECT 1822.605 1424.655 1822.895 1424.700 ;
        RECT 1823.050 1424.640 1823.370 1424.700 ;
        RECT 1822.590 1400.700 1822.910 1400.760 ;
        RECT 1823.050 1400.700 1823.370 1400.760 ;
        RECT 1822.590 1400.560 1823.370 1400.700 ;
        RECT 1822.590 1400.500 1822.910 1400.560 ;
        RECT 1823.050 1400.500 1823.370 1400.560 ;
        RECT 1822.590 1249.400 1822.910 1249.460 ;
        RECT 1823.050 1249.400 1823.370 1249.460 ;
        RECT 1822.590 1249.260 1823.370 1249.400 ;
        RECT 1822.590 1249.200 1822.910 1249.260 ;
        RECT 1823.050 1249.200 1823.370 1249.260 ;
        RECT 1822.590 1221.320 1822.910 1221.580 ;
        RECT 1822.680 1220.840 1822.820 1221.320 ;
        RECT 1823.050 1220.840 1823.370 1220.900 ;
        RECT 1822.680 1220.700 1823.370 1220.840 ;
        RECT 1823.050 1220.640 1823.370 1220.700 ;
        RECT 1823.050 1159.100 1823.370 1159.360 ;
        RECT 1822.590 1158.960 1822.910 1159.020 ;
        RECT 1823.140 1158.960 1823.280 1159.100 ;
        RECT 1822.590 1158.820 1823.280 1158.960 ;
        RECT 1822.590 1158.760 1822.910 1158.820 ;
        RECT 1822.130 1104.220 1822.450 1104.280 ;
        RECT 1823.510 1104.220 1823.830 1104.280 ;
        RECT 1822.130 1104.080 1823.830 1104.220 ;
        RECT 1822.130 1104.020 1822.450 1104.080 ;
        RECT 1823.510 1104.020 1823.830 1104.080 ;
        RECT 1820.765 1062.740 1821.055 1062.785 ;
        RECT 1822.130 1062.740 1822.450 1062.800 ;
        RECT 1820.765 1062.600 1822.450 1062.740 ;
        RECT 1820.765 1062.555 1821.055 1062.600 ;
        RECT 1822.130 1062.540 1822.450 1062.600 ;
        RECT 1820.750 1042.000 1821.070 1042.060 ;
        RECT 1820.555 1041.860 1821.070 1042.000 ;
        RECT 1820.750 1041.800 1821.070 1041.860 ;
        RECT 1820.750 1014.460 1821.070 1014.520 ;
        RECT 1823.050 1014.460 1823.370 1014.520 ;
        RECT 1820.750 1014.320 1823.370 1014.460 ;
        RECT 1820.750 1014.260 1821.070 1014.320 ;
        RECT 1823.050 1014.260 1823.370 1014.320 ;
        RECT 1823.050 980.460 1823.370 980.520 ;
        RECT 1823.970 980.460 1824.290 980.520 ;
        RECT 1823.050 980.320 1824.290 980.460 ;
        RECT 1823.050 980.260 1823.370 980.320 ;
        RECT 1823.970 980.260 1824.290 980.320 ;
        RECT 1822.590 952.240 1822.910 952.300 ;
        RECT 1822.395 952.100 1822.910 952.240 ;
        RECT 1822.590 952.040 1822.910 952.100 ;
        RECT 1822.590 931.500 1822.910 931.560 ;
        RECT 1822.395 931.360 1822.910 931.500 ;
        RECT 1822.590 931.300 1822.910 931.360 ;
        RECT 1823.050 883.700 1823.370 883.960 ;
        RECT 1823.140 883.280 1823.280 883.700 ;
        RECT 1823.050 883.020 1823.370 883.280 ;
        RECT 1822.590 738.180 1822.910 738.440 ;
        RECT 1822.680 738.040 1822.820 738.180 ;
        RECT 1823.050 738.040 1823.370 738.100 ;
        RECT 1822.680 737.900 1823.370 738.040 ;
        RECT 1823.050 737.840 1823.370 737.900 ;
        RECT 1822.590 724.440 1822.910 724.500 ;
        RECT 1823.050 724.440 1823.370 724.500 ;
        RECT 1822.590 724.300 1823.370 724.440 ;
        RECT 1822.590 724.240 1822.910 724.300 ;
        RECT 1823.050 724.240 1823.370 724.300 ;
        RECT 1822.590 628.020 1822.910 628.280 ;
        RECT 1822.680 627.540 1822.820 628.020 ;
        RECT 1823.050 627.540 1823.370 627.600 ;
        RECT 1822.680 627.400 1823.370 627.540 ;
        RECT 1823.050 627.340 1823.370 627.400 ;
        RECT 1822.590 545.600 1822.910 545.660 ;
        RECT 1823.510 545.600 1823.830 545.660 ;
        RECT 1822.590 545.460 1823.830 545.600 ;
        RECT 1822.590 545.400 1822.910 545.460 ;
        RECT 1823.510 545.400 1823.830 545.460 ;
        RECT 1822.590 518.740 1822.910 518.800 ;
        RECT 1823.510 518.740 1823.830 518.800 ;
        RECT 1822.590 518.600 1823.830 518.740 ;
        RECT 1822.590 518.540 1822.910 518.600 ;
        RECT 1823.510 518.540 1823.830 518.600 ;
        RECT 1822.605 469.100 1822.895 469.145 ;
        RECT 1823.510 469.100 1823.830 469.160 ;
        RECT 1822.605 468.960 1823.830 469.100 ;
        RECT 1822.605 468.915 1822.895 468.960 ;
        RECT 1823.510 468.900 1823.830 468.960 ;
        RECT 1822.590 421.160 1822.910 421.220 ;
        RECT 1822.395 421.020 1822.910 421.160 ;
        RECT 1822.590 420.960 1822.910 421.020 ;
        RECT 1822.590 372.540 1822.910 372.600 ;
        RECT 1822.395 372.400 1822.910 372.540 ;
        RECT 1822.590 372.340 1822.910 372.400 ;
        RECT 1822.590 324.600 1822.910 324.660 ;
        RECT 1822.395 324.460 1822.910 324.600 ;
        RECT 1822.590 324.400 1822.910 324.460 ;
        RECT 1823.050 180.100 1823.370 180.160 ;
        RECT 1822.680 179.960 1823.370 180.100 ;
        RECT 1822.680 179.820 1822.820 179.960 ;
        RECT 1823.050 179.900 1823.370 179.960 ;
        RECT 1822.590 179.560 1822.910 179.820 ;
        RECT 1823.970 131.140 1824.290 131.200 ;
        RECT 1823.775 131.000 1824.290 131.140 ;
        RECT 1823.970 130.940 1824.290 131.000 ;
        RECT 1823.970 87.280 1824.290 87.340 ;
        RECT 1823.775 87.140 1824.290 87.280 ;
        RECT 1823.970 87.080 1824.290 87.140 ;
        RECT 1822.130 41.720 1822.450 41.780 ;
        RECT 1823.970 41.720 1824.290 41.780 ;
        RECT 1822.130 41.580 1824.290 41.720 ;
        RECT 1822.130 41.520 1822.450 41.580 ;
        RECT 1823.970 41.520 1824.290 41.580 ;
        RECT 1317.050 40.360 1317.370 40.420 ;
        RECT 1822.130 40.360 1822.450 40.420 ;
        RECT 1317.050 40.220 1822.450 40.360 ;
        RECT 1317.050 40.160 1317.370 40.220 ;
        RECT 1822.130 40.160 1822.450 40.220 ;
      LAYER via ;
        RECT 1823.080 1642.240 1823.340 1642.500 ;
        RECT 1824.000 1642.240 1824.260 1642.500 ;
        RECT 1822.620 1545.680 1822.880 1545.940 ;
        RECT 1823.080 1545.680 1823.340 1545.940 ;
        RECT 1822.620 1538.540 1822.880 1538.800 ;
        RECT 1823.080 1490.600 1823.340 1490.860 ;
        RECT 1822.620 1456.600 1822.880 1456.860 ;
        RECT 1823.080 1424.640 1823.340 1424.900 ;
        RECT 1822.620 1400.500 1822.880 1400.760 ;
        RECT 1823.080 1400.500 1823.340 1400.760 ;
        RECT 1822.620 1249.200 1822.880 1249.460 ;
        RECT 1823.080 1249.200 1823.340 1249.460 ;
        RECT 1822.620 1221.320 1822.880 1221.580 ;
        RECT 1823.080 1220.640 1823.340 1220.900 ;
        RECT 1823.080 1159.100 1823.340 1159.360 ;
        RECT 1822.620 1158.760 1822.880 1159.020 ;
        RECT 1822.160 1104.020 1822.420 1104.280 ;
        RECT 1823.540 1104.020 1823.800 1104.280 ;
        RECT 1822.160 1062.540 1822.420 1062.800 ;
        RECT 1820.780 1041.800 1821.040 1042.060 ;
        RECT 1820.780 1014.260 1821.040 1014.520 ;
        RECT 1823.080 1014.260 1823.340 1014.520 ;
        RECT 1823.080 980.260 1823.340 980.520 ;
        RECT 1824.000 980.260 1824.260 980.520 ;
        RECT 1822.620 952.040 1822.880 952.300 ;
        RECT 1822.620 931.300 1822.880 931.560 ;
        RECT 1823.080 883.700 1823.340 883.960 ;
        RECT 1823.080 883.020 1823.340 883.280 ;
        RECT 1822.620 738.180 1822.880 738.440 ;
        RECT 1823.080 737.840 1823.340 738.100 ;
        RECT 1822.620 724.240 1822.880 724.500 ;
        RECT 1823.080 724.240 1823.340 724.500 ;
        RECT 1822.620 628.020 1822.880 628.280 ;
        RECT 1823.080 627.340 1823.340 627.600 ;
        RECT 1822.620 545.400 1822.880 545.660 ;
        RECT 1823.540 545.400 1823.800 545.660 ;
        RECT 1822.620 518.540 1822.880 518.800 ;
        RECT 1823.540 518.540 1823.800 518.800 ;
        RECT 1823.540 468.900 1823.800 469.160 ;
        RECT 1822.620 420.960 1822.880 421.220 ;
        RECT 1822.620 372.340 1822.880 372.600 ;
        RECT 1822.620 324.400 1822.880 324.660 ;
        RECT 1823.080 179.900 1823.340 180.160 ;
        RECT 1822.620 179.560 1822.880 179.820 ;
        RECT 1824.000 130.940 1824.260 131.200 ;
        RECT 1824.000 87.080 1824.260 87.340 ;
        RECT 1822.160 41.520 1822.420 41.780 ;
        RECT 1824.000 41.520 1824.260 41.780 ;
        RECT 1317.080 40.160 1317.340 40.420 ;
        RECT 1822.160 40.160 1822.420 40.420 ;
      LAYER met2 ;
        RECT 1826.220 1701.090 1826.500 1704.000 ;
        RECT 1824.060 1700.950 1826.500 1701.090 ;
        RECT 1824.060 1642.530 1824.200 1700.950 ;
        RECT 1826.220 1700.000 1826.500 1700.950 ;
        RECT 1823.080 1642.210 1823.340 1642.530 ;
        RECT 1824.000 1642.210 1824.260 1642.530 ;
        RECT 1823.140 1545.970 1823.280 1642.210 ;
        RECT 1822.620 1545.650 1822.880 1545.970 ;
        RECT 1823.080 1545.650 1823.340 1545.970 ;
        RECT 1822.680 1538.830 1822.820 1545.650 ;
        RECT 1822.620 1538.510 1822.880 1538.830 ;
        RECT 1823.080 1490.570 1823.340 1490.890 ;
        RECT 1823.140 1490.290 1823.280 1490.570 ;
        RECT 1822.680 1490.150 1823.280 1490.290 ;
        RECT 1822.680 1456.890 1822.820 1490.150 ;
        RECT 1822.620 1456.570 1822.880 1456.890 ;
        RECT 1823.080 1424.610 1823.340 1424.930 ;
        RECT 1823.140 1400.790 1823.280 1424.610 ;
        RECT 1822.620 1400.470 1822.880 1400.790 ;
        RECT 1823.080 1400.470 1823.340 1400.790 ;
        RECT 1822.680 1353.725 1822.820 1400.470 ;
        RECT 1822.610 1353.355 1822.890 1353.725 ;
        RECT 1823.070 1351.995 1823.350 1352.365 ;
        RECT 1823.140 1249.490 1823.280 1351.995 ;
        RECT 1822.620 1249.170 1822.880 1249.490 ;
        RECT 1823.080 1249.170 1823.340 1249.490 ;
        RECT 1822.680 1221.610 1822.820 1249.170 ;
        RECT 1822.620 1221.290 1822.880 1221.610 ;
        RECT 1823.080 1220.610 1823.340 1220.930 ;
        RECT 1823.140 1159.390 1823.280 1220.610 ;
        RECT 1823.080 1159.070 1823.340 1159.390 ;
        RECT 1822.620 1158.730 1822.880 1159.050 ;
        RECT 1822.680 1145.530 1822.820 1158.730 ;
        RECT 1822.680 1145.390 1823.740 1145.530 ;
        RECT 1823.600 1104.310 1823.740 1145.390 ;
        RECT 1822.160 1103.990 1822.420 1104.310 ;
        RECT 1823.540 1103.990 1823.800 1104.310 ;
        RECT 1822.220 1062.830 1822.360 1103.990 ;
        RECT 1822.160 1062.510 1822.420 1062.830 ;
        RECT 1820.780 1041.770 1821.040 1042.090 ;
        RECT 1820.840 1014.550 1820.980 1041.770 ;
        RECT 1820.780 1014.230 1821.040 1014.550 ;
        RECT 1823.080 1014.230 1823.340 1014.550 ;
        RECT 1823.140 980.550 1823.280 1014.230 ;
        RECT 1823.080 980.230 1823.340 980.550 ;
        RECT 1824.000 980.230 1824.260 980.550 ;
        RECT 1824.060 952.525 1824.200 980.230 ;
        RECT 1823.070 952.410 1823.350 952.525 ;
        RECT 1822.680 952.330 1823.350 952.410 ;
        RECT 1822.620 952.270 1823.350 952.330 ;
        RECT 1822.620 952.010 1822.880 952.270 ;
        RECT 1823.070 952.155 1823.350 952.270 ;
        RECT 1823.990 952.155 1824.270 952.525 ;
        RECT 1822.680 951.855 1822.820 952.010 ;
        RECT 1822.620 931.270 1822.880 931.590 ;
        RECT 1822.680 904.130 1822.820 931.270 ;
        RECT 1822.680 903.990 1823.280 904.130 ;
        RECT 1823.140 883.990 1823.280 903.990 ;
        RECT 1823.080 883.670 1823.340 883.990 ;
        RECT 1823.080 882.990 1823.340 883.310 ;
        RECT 1823.140 783.770 1823.280 882.990 ;
        RECT 1822.680 783.630 1823.280 783.770 ;
        RECT 1822.680 738.470 1822.820 783.630 ;
        RECT 1822.620 738.150 1822.880 738.470 ;
        RECT 1823.080 737.810 1823.340 738.130 ;
        RECT 1823.140 724.530 1823.280 737.810 ;
        RECT 1822.620 724.210 1822.880 724.530 ;
        RECT 1823.080 724.210 1823.340 724.530 ;
        RECT 1822.680 628.310 1822.820 724.210 ;
        RECT 1822.620 627.990 1822.880 628.310 ;
        RECT 1823.080 627.310 1823.340 627.630 ;
        RECT 1823.140 572.290 1823.280 627.310 ;
        RECT 1823.140 572.150 1823.740 572.290 ;
        RECT 1823.600 545.690 1823.740 572.150 ;
        RECT 1822.620 545.370 1822.880 545.690 ;
        RECT 1823.540 545.370 1823.800 545.690 ;
        RECT 1822.680 518.830 1822.820 545.370 ;
        RECT 1822.620 518.510 1822.880 518.830 ;
        RECT 1823.540 518.510 1823.800 518.830 ;
        RECT 1823.600 469.190 1823.740 518.510 ;
        RECT 1823.540 468.870 1823.800 469.190 ;
        RECT 1822.620 420.930 1822.880 421.250 ;
        RECT 1822.680 372.630 1822.820 420.930 ;
        RECT 1822.620 372.310 1822.880 372.630 ;
        RECT 1822.620 324.370 1822.880 324.690 ;
        RECT 1822.680 304.370 1822.820 324.370 ;
        RECT 1822.680 304.230 1823.280 304.370 ;
        RECT 1823.140 298.930 1823.280 304.230 ;
        RECT 1822.680 298.790 1823.280 298.930 ;
        RECT 1822.680 265.610 1822.820 298.790 ;
        RECT 1822.680 265.470 1823.280 265.610 ;
        RECT 1823.140 180.190 1823.280 265.470 ;
        RECT 1823.080 179.870 1823.340 180.190 ;
        RECT 1822.620 179.530 1822.880 179.850 ;
        RECT 1822.680 155.450 1822.820 179.530 ;
        RECT 1822.680 155.310 1824.200 155.450 ;
        RECT 1824.060 131.230 1824.200 155.310 ;
        RECT 1824.000 130.910 1824.260 131.230 ;
        RECT 1824.000 87.050 1824.260 87.370 ;
        RECT 1824.060 41.810 1824.200 87.050 ;
        RECT 1822.160 41.490 1822.420 41.810 ;
        RECT 1824.000 41.490 1824.260 41.810 ;
        RECT 1822.220 40.450 1822.360 41.490 ;
        RECT 1317.080 40.130 1317.340 40.450 ;
        RECT 1822.160 40.130 1822.420 40.450 ;
        RECT 1317.140 2.400 1317.280 40.130 ;
        RECT 1316.930 -4.800 1317.490 2.400 ;
      LAYER via2 ;
        RECT 1822.610 1353.400 1822.890 1353.680 ;
        RECT 1823.070 1352.040 1823.350 1352.320 ;
        RECT 1823.070 952.200 1823.350 952.480 ;
        RECT 1823.990 952.200 1824.270 952.480 ;
      LAYER met3 ;
        RECT 1822.585 1353.690 1822.915 1353.705 ;
        RECT 1821.910 1353.390 1822.915 1353.690 ;
        RECT 1821.910 1352.330 1822.210 1353.390 ;
        RECT 1822.585 1353.375 1822.915 1353.390 ;
        RECT 1823.045 1352.330 1823.375 1352.345 ;
        RECT 1821.910 1352.030 1823.375 1352.330 ;
        RECT 1823.045 1352.015 1823.375 1352.030 ;
        RECT 1823.045 952.490 1823.375 952.505 ;
        RECT 1823.965 952.490 1824.295 952.505 ;
        RECT 1823.045 952.190 1824.295 952.490 ;
        RECT 1823.045 952.175 1823.375 952.190 ;
        RECT 1823.965 952.175 1824.295 952.190 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1334.990 40.700 1335.310 40.760 ;
        RECT 1835.470 40.700 1835.790 40.760 ;
        RECT 1334.990 40.560 1835.790 40.700 ;
        RECT 1334.990 40.500 1335.310 40.560 ;
        RECT 1835.470 40.500 1835.790 40.560 ;
      LAYER via ;
        RECT 1335.020 40.500 1335.280 40.760 ;
        RECT 1835.500 40.500 1835.760 40.760 ;
      LAYER met2 ;
        RECT 1835.420 1700.000 1835.700 1704.000 ;
        RECT 1835.560 40.790 1835.700 1700.000 ;
        RECT 1335.020 40.470 1335.280 40.790 ;
        RECT 1835.500 40.470 1835.760 40.790 ;
        RECT 1335.080 2.400 1335.220 40.470 ;
        RECT 1334.870 -4.800 1335.430 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 692.370 36.620 692.690 36.680 ;
        RECT 1504.270 36.620 1504.590 36.680 ;
        RECT 692.370 36.480 1504.590 36.620 ;
        RECT 692.370 36.420 692.690 36.480 ;
        RECT 1504.270 36.420 1504.590 36.480 ;
      LAYER via ;
        RECT 692.400 36.420 692.660 36.680 ;
        RECT 1504.300 36.420 1504.560 36.680 ;
      LAYER met2 ;
        RECT 1504.680 1700.410 1504.960 1704.000 ;
        RECT 1504.360 1700.270 1504.960 1700.410 ;
        RECT 1504.360 36.710 1504.500 1700.270 ;
        RECT 1504.680 1700.000 1504.960 1700.270 ;
        RECT 692.400 36.390 692.660 36.710 ;
        RECT 1504.300 36.390 1504.560 36.710 ;
        RECT 692.460 2.400 692.600 36.390 ;
        RECT 692.250 -4.800 692.810 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1352.470 41.040 1352.790 41.100 ;
        RECT 1842.830 41.040 1843.150 41.100 ;
        RECT 1352.470 40.900 1843.150 41.040 ;
        RECT 1352.470 40.840 1352.790 40.900 ;
        RECT 1842.830 40.840 1843.150 40.900 ;
      LAYER via ;
        RECT 1352.500 40.840 1352.760 41.100 ;
        RECT 1842.860 40.840 1843.120 41.100 ;
      LAYER met2 ;
        RECT 1844.620 1700.410 1844.900 1704.000 ;
        RECT 1842.920 1700.270 1844.900 1700.410 ;
        RECT 1842.920 41.130 1843.060 1700.270 ;
        RECT 1844.620 1700.000 1844.900 1700.270 ;
        RECT 1352.500 40.810 1352.760 41.130 ;
        RECT 1842.860 40.810 1843.120 41.130 ;
        RECT 1352.560 2.400 1352.700 40.810 ;
        RECT 1352.350 -4.800 1352.910 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1850.265 1442.025 1850.435 1490.475 ;
        RECT 1850.265 1242.445 1850.435 1270.155 ;
        RECT 1849.805 1014.305 1849.975 1062.415 ;
        RECT 1849.805 965.685 1849.975 1007.335 ;
        RECT 1850.265 772.905 1850.435 821.015 ;
        RECT 1849.805 41.225 1849.975 48.195 ;
      LAYER mcon ;
        RECT 1850.265 1490.305 1850.435 1490.475 ;
        RECT 1850.265 1269.985 1850.435 1270.155 ;
        RECT 1849.805 1062.245 1849.975 1062.415 ;
        RECT 1849.805 1007.165 1849.975 1007.335 ;
        RECT 1850.265 820.845 1850.435 821.015 ;
        RECT 1849.805 48.025 1849.975 48.195 ;
      LAYER met1 ;
        RECT 1850.650 1642.440 1850.970 1642.500 ;
        RECT 1851.570 1642.440 1851.890 1642.500 ;
        RECT 1850.650 1642.300 1851.890 1642.440 ;
        RECT 1850.650 1642.240 1850.970 1642.300 ;
        RECT 1851.570 1642.240 1851.890 1642.300 ;
        RECT 1850.190 1497.260 1850.510 1497.320 ;
        RECT 1850.650 1497.260 1850.970 1497.320 ;
        RECT 1850.190 1497.120 1850.970 1497.260 ;
        RECT 1850.190 1497.060 1850.510 1497.120 ;
        RECT 1850.650 1497.060 1850.970 1497.120 ;
        RECT 1850.190 1490.460 1850.510 1490.520 ;
        RECT 1849.995 1490.320 1850.510 1490.460 ;
        RECT 1850.190 1490.260 1850.510 1490.320 ;
        RECT 1850.190 1442.180 1850.510 1442.240 ;
        RECT 1849.995 1442.040 1850.510 1442.180 ;
        RECT 1850.190 1441.980 1850.510 1442.040 ;
        RECT 1850.190 1414.440 1850.510 1414.700 ;
        RECT 1850.280 1413.960 1850.420 1414.440 ;
        RECT 1850.650 1413.960 1850.970 1414.020 ;
        RECT 1850.280 1413.820 1850.970 1413.960 ;
        RECT 1850.650 1413.760 1850.970 1413.820 ;
        RECT 1848.810 1400.700 1849.130 1400.760 ;
        RECT 1850.650 1400.700 1850.970 1400.760 ;
        RECT 1848.810 1400.560 1850.970 1400.700 ;
        RECT 1848.810 1400.500 1849.130 1400.560 ;
        RECT 1850.650 1400.500 1850.970 1400.560 ;
        RECT 1848.810 1374.180 1849.130 1374.240 ;
        RECT 1850.650 1374.180 1850.970 1374.240 ;
        RECT 1848.810 1374.040 1850.970 1374.180 ;
        RECT 1848.810 1373.980 1849.130 1374.040 ;
        RECT 1850.650 1373.980 1850.970 1374.040 ;
        RECT 1850.205 1270.140 1850.495 1270.185 ;
        RECT 1850.650 1270.140 1850.970 1270.200 ;
        RECT 1850.205 1270.000 1850.970 1270.140 ;
        RECT 1850.205 1269.955 1850.495 1270.000 ;
        RECT 1850.650 1269.940 1850.970 1270.000 ;
        RECT 1850.190 1242.600 1850.510 1242.660 ;
        RECT 1849.995 1242.460 1850.510 1242.600 ;
        RECT 1850.190 1242.400 1850.510 1242.460 ;
        RECT 1850.190 1241.920 1850.510 1241.980 ;
        RECT 1851.570 1241.920 1851.890 1241.980 ;
        RECT 1850.190 1241.780 1851.890 1241.920 ;
        RECT 1850.190 1241.720 1850.510 1241.780 ;
        RECT 1851.570 1241.720 1851.890 1241.780 ;
        RECT 1848.810 1169.500 1849.130 1169.560 ;
        RECT 1851.570 1169.500 1851.890 1169.560 ;
        RECT 1848.810 1169.360 1851.890 1169.500 ;
        RECT 1848.810 1169.300 1849.130 1169.360 ;
        RECT 1851.570 1169.300 1851.890 1169.360 ;
        RECT 1848.810 1104.220 1849.130 1104.280 ;
        RECT 1849.730 1104.220 1850.050 1104.280 ;
        RECT 1848.810 1104.080 1850.050 1104.220 ;
        RECT 1848.810 1104.020 1849.130 1104.080 ;
        RECT 1849.730 1104.020 1850.050 1104.080 ;
        RECT 1849.730 1062.400 1850.050 1062.460 ;
        RECT 1849.535 1062.260 1850.050 1062.400 ;
        RECT 1849.730 1062.200 1850.050 1062.260 ;
        RECT 1849.730 1014.460 1850.050 1014.520 ;
        RECT 1849.535 1014.320 1850.050 1014.460 ;
        RECT 1849.730 1014.260 1850.050 1014.320 ;
        RECT 1849.730 1007.320 1850.050 1007.380 ;
        RECT 1849.535 1007.180 1850.050 1007.320 ;
        RECT 1849.730 1007.120 1850.050 1007.180 ;
        RECT 1849.730 965.840 1850.050 965.900 ;
        RECT 1849.535 965.700 1850.050 965.840 ;
        RECT 1849.730 965.640 1850.050 965.700 ;
        RECT 1850.190 869.620 1850.510 869.680 ;
        RECT 1850.650 869.620 1850.970 869.680 ;
        RECT 1850.190 869.480 1850.970 869.620 ;
        RECT 1850.190 869.420 1850.510 869.480 ;
        RECT 1850.650 869.420 1850.970 869.480 ;
        RECT 1850.205 821.000 1850.495 821.045 ;
        RECT 1850.650 821.000 1850.970 821.060 ;
        RECT 1850.205 820.860 1850.970 821.000 ;
        RECT 1850.205 820.815 1850.495 820.860 ;
        RECT 1850.650 820.800 1850.970 820.860 ;
        RECT 1850.190 773.060 1850.510 773.120 ;
        RECT 1849.995 772.920 1850.510 773.060 ;
        RECT 1850.190 772.860 1850.510 772.920 ;
        RECT 1850.190 738.180 1850.510 738.440 ;
        RECT 1850.280 738.040 1850.420 738.180 ;
        RECT 1850.650 738.040 1850.970 738.100 ;
        RECT 1850.280 737.900 1850.970 738.040 ;
        RECT 1850.650 737.840 1850.970 737.900 ;
        RECT 1850.650 724.440 1850.970 724.500 ;
        RECT 1851.110 724.440 1851.430 724.500 ;
        RECT 1850.650 724.300 1851.430 724.440 ;
        RECT 1850.650 724.240 1850.970 724.300 ;
        RECT 1851.110 724.240 1851.430 724.300 ;
        RECT 1849.730 627.880 1850.050 627.940 ;
        RECT 1850.650 627.880 1850.970 627.940 ;
        RECT 1849.730 627.740 1850.970 627.880 ;
        RECT 1849.730 627.680 1850.050 627.740 ;
        RECT 1850.650 627.680 1850.970 627.740 ;
        RECT 1849.730 573.140 1850.050 573.200 ;
        RECT 1849.730 573.000 1850.420 573.140 ;
        RECT 1849.730 572.940 1850.050 573.000 ;
        RECT 1850.280 572.860 1850.420 573.000 ;
        RECT 1850.190 572.600 1850.510 572.860 ;
        RECT 1850.190 531.460 1850.510 531.720 ;
        RECT 1850.280 530.980 1850.420 531.460 ;
        RECT 1850.650 530.980 1850.970 531.040 ;
        RECT 1850.280 530.840 1850.970 530.980 ;
        RECT 1850.650 530.780 1850.970 530.840 ;
        RECT 1850.650 517.380 1850.970 517.440 ;
        RECT 1851.570 517.380 1851.890 517.440 ;
        RECT 1850.650 517.240 1851.890 517.380 ;
        RECT 1850.650 517.180 1850.970 517.240 ;
        RECT 1851.570 517.180 1851.890 517.240 ;
        RECT 1850.190 380.020 1850.510 380.080 ;
        RECT 1851.570 380.020 1851.890 380.080 ;
        RECT 1850.190 379.880 1851.890 380.020 ;
        RECT 1850.190 379.820 1850.510 379.880 ;
        RECT 1851.570 379.820 1851.890 379.880 ;
        RECT 1850.190 331.880 1850.510 332.140 ;
        RECT 1850.280 331.460 1850.420 331.880 ;
        RECT 1850.190 331.200 1850.510 331.460 ;
        RECT 1850.190 234.840 1850.510 234.900 ;
        RECT 1850.650 234.840 1850.970 234.900 ;
        RECT 1850.190 234.700 1850.970 234.840 ;
        RECT 1850.190 234.640 1850.510 234.700 ;
        RECT 1850.650 234.640 1850.970 234.700 ;
        RECT 1850.190 179.760 1850.510 179.820 ;
        RECT 1850.650 179.760 1850.970 179.820 ;
        RECT 1850.190 179.620 1850.970 179.760 ;
        RECT 1850.190 179.560 1850.510 179.620 ;
        RECT 1850.650 179.560 1850.970 179.620 ;
        RECT 1850.190 62.460 1850.510 62.520 ;
        RECT 1849.820 62.320 1850.510 62.460 ;
        RECT 1849.820 62.180 1849.960 62.320 ;
        RECT 1850.190 62.260 1850.510 62.320 ;
        RECT 1849.730 61.920 1850.050 62.180 ;
        RECT 1849.730 48.180 1850.050 48.240 ;
        RECT 1849.535 48.040 1850.050 48.180 ;
        RECT 1849.730 47.980 1850.050 48.040 ;
        RECT 1370.410 41.380 1370.730 41.440 ;
        RECT 1849.745 41.380 1850.035 41.425 ;
        RECT 1370.410 41.240 1850.035 41.380 ;
        RECT 1370.410 41.180 1370.730 41.240 ;
        RECT 1849.745 41.195 1850.035 41.240 ;
      LAYER via ;
        RECT 1850.680 1642.240 1850.940 1642.500 ;
        RECT 1851.600 1642.240 1851.860 1642.500 ;
        RECT 1850.220 1497.060 1850.480 1497.320 ;
        RECT 1850.680 1497.060 1850.940 1497.320 ;
        RECT 1850.220 1490.260 1850.480 1490.520 ;
        RECT 1850.220 1441.980 1850.480 1442.240 ;
        RECT 1850.220 1414.440 1850.480 1414.700 ;
        RECT 1850.680 1413.760 1850.940 1414.020 ;
        RECT 1848.840 1400.500 1849.100 1400.760 ;
        RECT 1850.680 1400.500 1850.940 1400.760 ;
        RECT 1848.840 1373.980 1849.100 1374.240 ;
        RECT 1850.680 1373.980 1850.940 1374.240 ;
        RECT 1850.680 1269.940 1850.940 1270.200 ;
        RECT 1850.220 1242.400 1850.480 1242.660 ;
        RECT 1850.220 1241.720 1850.480 1241.980 ;
        RECT 1851.600 1241.720 1851.860 1241.980 ;
        RECT 1848.840 1169.300 1849.100 1169.560 ;
        RECT 1851.600 1169.300 1851.860 1169.560 ;
        RECT 1848.840 1104.020 1849.100 1104.280 ;
        RECT 1849.760 1104.020 1850.020 1104.280 ;
        RECT 1849.760 1062.200 1850.020 1062.460 ;
        RECT 1849.760 1014.260 1850.020 1014.520 ;
        RECT 1849.760 1007.120 1850.020 1007.380 ;
        RECT 1849.760 965.640 1850.020 965.900 ;
        RECT 1850.220 869.420 1850.480 869.680 ;
        RECT 1850.680 869.420 1850.940 869.680 ;
        RECT 1850.680 820.800 1850.940 821.060 ;
        RECT 1850.220 772.860 1850.480 773.120 ;
        RECT 1850.220 738.180 1850.480 738.440 ;
        RECT 1850.680 737.840 1850.940 738.100 ;
        RECT 1850.680 724.240 1850.940 724.500 ;
        RECT 1851.140 724.240 1851.400 724.500 ;
        RECT 1849.760 627.680 1850.020 627.940 ;
        RECT 1850.680 627.680 1850.940 627.940 ;
        RECT 1849.760 572.940 1850.020 573.200 ;
        RECT 1850.220 572.600 1850.480 572.860 ;
        RECT 1850.220 531.460 1850.480 531.720 ;
        RECT 1850.680 530.780 1850.940 531.040 ;
        RECT 1850.680 517.180 1850.940 517.440 ;
        RECT 1851.600 517.180 1851.860 517.440 ;
        RECT 1850.220 379.820 1850.480 380.080 ;
        RECT 1851.600 379.820 1851.860 380.080 ;
        RECT 1850.220 331.880 1850.480 332.140 ;
        RECT 1850.220 331.200 1850.480 331.460 ;
        RECT 1850.220 234.640 1850.480 234.900 ;
        RECT 1850.680 234.640 1850.940 234.900 ;
        RECT 1850.220 179.560 1850.480 179.820 ;
        RECT 1850.680 179.560 1850.940 179.820 ;
        RECT 1850.220 62.260 1850.480 62.520 ;
        RECT 1849.760 61.920 1850.020 62.180 ;
        RECT 1849.760 47.980 1850.020 48.240 ;
        RECT 1370.440 41.180 1370.700 41.440 ;
      LAYER met2 ;
        RECT 1853.820 1701.090 1854.100 1704.000 ;
        RECT 1851.660 1700.950 1854.100 1701.090 ;
        RECT 1851.660 1642.530 1851.800 1700.950 ;
        RECT 1853.820 1700.000 1854.100 1700.950 ;
        RECT 1850.680 1642.210 1850.940 1642.530 ;
        RECT 1851.600 1642.210 1851.860 1642.530 ;
        RECT 1850.740 1497.350 1850.880 1642.210 ;
        RECT 1850.220 1497.030 1850.480 1497.350 ;
        RECT 1850.680 1497.030 1850.940 1497.350 ;
        RECT 1850.280 1490.550 1850.420 1497.030 ;
        RECT 1850.220 1490.230 1850.480 1490.550 ;
        RECT 1850.220 1441.950 1850.480 1442.270 ;
        RECT 1850.280 1414.730 1850.420 1441.950 ;
        RECT 1850.220 1414.410 1850.480 1414.730 ;
        RECT 1850.680 1413.730 1850.940 1414.050 ;
        RECT 1850.740 1400.790 1850.880 1413.730 ;
        RECT 1848.840 1400.470 1849.100 1400.790 ;
        RECT 1850.680 1400.470 1850.940 1400.790 ;
        RECT 1848.900 1374.270 1849.040 1400.470 ;
        RECT 1848.840 1373.950 1849.100 1374.270 ;
        RECT 1850.680 1373.950 1850.940 1374.270 ;
        RECT 1850.740 1338.765 1850.880 1373.950 ;
        RECT 1849.750 1338.395 1850.030 1338.765 ;
        RECT 1850.670 1338.395 1850.950 1338.765 ;
        RECT 1849.820 1290.485 1849.960 1338.395 ;
        RECT 1849.750 1290.115 1850.030 1290.485 ;
        RECT 1850.670 1290.115 1850.950 1290.485 ;
        RECT 1850.740 1270.230 1850.880 1290.115 ;
        RECT 1850.680 1269.910 1850.940 1270.230 ;
        RECT 1850.220 1242.370 1850.480 1242.690 ;
        RECT 1850.280 1242.010 1850.420 1242.370 ;
        RECT 1850.220 1241.690 1850.480 1242.010 ;
        RECT 1851.600 1241.690 1851.860 1242.010 ;
        RECT 1851.660 1169.590 1851.800 1241.690 ;
        RECT 1848.840 1169.270 1849.100 1169.590 ;
        RECT 1851.600 1169.270 1851.860 1169.590 ;
        RECT 1848.900 1104.310 1849.040 1169.270 ;
        RECT 1848.840 1103.990 1849.100 1104.310 ;
        RECT 1849.760 1103.990 1850.020 1104.310 ;
        RECT 1849.820 1062.490 1849.960 1103.990 ;
        RECT 1849.760 1062.170 1850.020 1062.490 ;
        RECT 1849.760 1014.230 1850.020 1014.550 ;
        RECT 1849.820 1007.410 1849.960 1014.230 ;
        RECT 1849.760 1007.090 1850.020 1007.410 ;
        RECT 1849.760 965.610 1850.020 965.930 ;
        RECT 1849.820 931.330 1849.960 965.610 ;
        RECT 1849.820 931.190 1850.880 931.330 ;
        RECT 1850.740 869.710 1850.880 931.190 ;
        RECT 1850.220 869.390 1850.480 869.710 ;
        RECT 1850.680 869.390 1850.940 869.710 ;
        RECT 1850.280 847.010 1850.420 869.390 ;
        RECT 1850.280 846.870 1850.880 847.010 ;
        RECT 1850.740 821.090 1850.880 846.870 ;
        RECT 1850.680 820.770 1850.940 821.090 ;
        RECT 1850.220 772.830 1850.480 773.150 ;
        RECT 1850.280 738.470 1850.420 772.830 ;
        RECT 1850.220 738.150 1850.480 738.470 ;
        RECT 1850.680 737.810 1850.940 738.130 ;
        RECT 1850.740 724.530 1850.880 737.810 ;
        RECT 1850.680 724.210 1850.940 724.530 ;
        RECT 1851.140 724.210 1851.400 724.530 ;
        RECT 1851.200 676.445 1851.340 724.210 ;
        RECT 1850.210 676.075 1850.490 676.445 ;
        RECT 1851.130 676.075 1851.410 676.445 ;
        RECT 1850.280 651.850 1850.420 676.075 ;
        RECT 1850.280 651.710 1851.340 651.850 ;
        RECT 1851.200 640.970 1851.340 651.710 ;
        RECT 1850.740 640.830 1851.340 640.970 ;
        RECT 1850.740 627.970 1850.880 640.830 ;
        RECT 1849.760 627.650 1850.020 627.970 ;
        RECT 1850.680 627.650 1850.940 627.970 ;
        RECT 1849.820 573.230 1849.960 627.650 ;
        RECT 1849.760 572.910 1850.020 573.230 ;
        RECT 1850.220 572.570 1850.480 572.890 ;
        RECT 1850.280 531.750 1850.420 572.570 ;
        RECT 1850.220 531.430 1850.480 531.750 ;
        RECT 1850.680 530.750 1850.940 531.070 ;
        RECT 1850.740 517.470 1850.880 530.750 ;
        RECT 1850.680 517.150 1850.940 517.470 ;
        RECT 1851.600 517.150 1851.860 517.470 ;
        RECT 1851.660 380.110 1851.800 517.150 ;
        RECT 1850.220 379.790 1850.480 380.110 ;
        RECT 1851.600 379.790 1851.860 380.110 ;
        RECT 1850.280 332.170 1850.420 379.790 ;
        RECT 1850.220 331.850 1850.480 332.170 ;
        RECT 1850.220 331.170 1850.480 331.490 ;
        RECT 1850.280 304.370 1850.420 331.170 ;
        RECT 1850.280 304.230 1850.880 304.370 ;
        RECT 1850.740 298.930 1850.880 304.230 ;
        RECT 1850.280 298.790 1850.880 298.930 ;
        RECT 1850.280 234.930 1850.420 298.790 ;
        RECT 1850.220 234.610 1850.480 234.930 ;
        RECT 1850.680 234.610 1850.940 234.930 ;
        RECT 1850.740 179.850 1850.880 234.610 ;
        RECT 1850.220 179.530 1850.480 179.850 ;
        RECT 1850.680 179.530 1850.940 179.850 ;
        RECT 1850.280 62.550 1850.420 179.530 ;
        RECT 1850.220 62.230 1850.480 62.550 ;
        RECT 1849.760 61.890 1850.020 62.210 ;
        RECT 1849.820 48.270 1849.960 61.890 ;
        RECT 1849.760 47.950 1850.020 48.270 ;
        RECT 1370.440 41.150 1370.700 41.470 ;
        RECT 1370.500 2.400 1370.640 41.150 ;
        RECT 1370.290 -4.800 1370.850 2.400 ;
      LAYER via2 ;
        RECT 1849.750 1338.440 1850.030 1338.720 ;
        RECT 1850.670 1338.440 1850.950 1338.720 ;
        RECT 1849.750 1290.160 1850.030 1290.440 ;
        RECT 1850.670 1290.160 1850.950 1290.440 ;
        RECT 1850.210 676.120 1850.490 676.400 ;
        RECT 1851.130 676.120 1851.410 676.400 ;
      LAYER met3 ;
        RECT 1849.725 1338.730 1850.055 1338.745 ;
        RECT 1850.645 1338.730 1850.975 1338.745 ;
        RECT 1849.725 1338.430 1850.975 1338.730 ;
        RECT 1849.725 1338.415 1850.055 1338.430 ;
        RECT 1850.645 1338.415 1850.975 1338.430 ;
        RECT 1849.725 1290.450 1850.055 1290.465 ;
        RECT 1850.645 1290.450 1850.975 1290.465 ;
        RECT 1849.725 1290.150 1850.975 1290.450 ;
        RECT 1849.725 1290.135 1850.055 1290.150 ;
        RECT 1850.645 1290.135 1850.975 1290.150 ;
        RECT 1850.185 676.410 1850.515 676.425 ;
        RECT 1851.105 676.410 1851.435 676.425 ;
        RECT 1850.185 676.110 1851.435 676.410 ;
        RECT 1850.185 676.095 1850.515 676.110 ;
        RECT 1851.105 676.095 1851.435 676.110 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1388.350 37.640 1388.670 37.700 ;
        RECT 1863.530 37.640 1863.850 37.700 ;
        RECT 1388.350 37.500 1863.850 37.640 ;
        RECT 1388.350 37.440 1388.670 37.500 ;
        RECT 1863.530 37.440 1863.850 37.500 ;
      LAYER via ;
        RECT 1388.380 37.440 1388.640 37.700 ;
        RECT 1863.560 37.440 1863.820 37.700 ;
      LAYER met2 ;
        RECT 1863.020 1700.410 1863.300 1704.000 ;
        RECT 1863.020 1700.270 1863.760 1700.410 ;
        RECT 1863.020 1700.000 1863.300 1700.270 ;
        RECT 1863.620 37.730 1863.760 1700.270 ;
        RECT 1388.380 37.410 1388.640 37.730 ;
        RECT 1863.560 37.410 1863.820 37.730 ;
        RECT 1388.440 2.400 1388.580 37.410 ;
        RECT 1388.230 -4.800 1388.790 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1406.290 37.300 1406.610 37.360 ;
        RECT 1870.430 37.300 1870.750 37.360 ;
        RECT 1406.290 37.160 1870.750 37.300 ;
        RECT 1406.290 37.100 1406.610 37.160 ;
        RECT 1870.430 37.100 1870.750 37.160 ;
      LAYER via ;
        RECT 1406.320 37.100 1406.580 37.360 ;
        RECT 1870.460 37.100 1870.720 37.360 ;
      LAYER met2 ;
        RECT 1872.220 1700.410 1872.500 1704.000 ;
        RECT 1870.520 1700.270 1872.500 1700.410 ;
        RECT 1870.520 37.390 1870.660 1700.270 ;
        RECT 1872.220 1700.000 1872.500 1700.270 ;
        RECT 1406.320 37.070 1406.580 37.390 ;
        RECT 1870.460 37.070 1870.720 37.390 ;
        RECT 1406.380 2.400 1406.520 37.070 ;
        RECT 1406.170 -4.800 1406.730 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1877.405 1448.825 1877.575 1490.475 ;
        RECT 1877.865 1242.445 1878.035 1270.155 ;
        RECT 1877.865 1213.885 1878.035 1241.935 ;
        RECT 1877.865 966.025 1878.035 980.475 ;
        RECT 1877.865 737.885 1878.035 772.735 ;
        RECT 1877.865 427.805 1878.035 467.755 ;
        RECT 1877.865 331.585 1878.035 379.355 ;
        RECT 1877.405 282.965 1877.575 331.075 ;
        RECT 1877.865 258.485 1878.035 282.455 ;
      LAYER mcon ;
        RECT 1877.405 1490.305 1877.575 1490.475 ;
        RECT 1877.865 1269.985 1878.035 1270.155 ;
        RECT 1877.865 1241.765 1878.035 1241.935 ;
        RECT 1877.865 980.305 1878.035 980.475 ;
        RECT 1877.865 772.565 1878.035 772.735 ;
        RECT 1877.865 467.585 1878.035 467.755 ;
        RECT 1877.865 379.185 1878.035 379.355 ;
        RECT 1877.405 330.905 1877.575 331.075 ;
        RECT 1877.865 282.285 1878.035 282.455 ;
      LAYER met1 ;
        RECT 1877.790 1594.160 1878.110 1594.220 ;
        RECT 1878.710 1594.160 1879.030 1594.220 ;
        RECT 1877.790 1594.020 1879.030 1594.160 ;
        RECT 1877.790 1593.960 1878.110 1594.020 ;
        RECT 1878.710 1593.960 1879.030 1594.020 ;
        RECT 1877.330 1490.460 1877.650 1490.520 ;
        RECT 1877.135 1490.320 1877.650 1490.460 ;
        RECT 1877.330 1490.260 1877.650 1490.320 ;
        RECT 1877.330 1448.980 1877.650 1449.040 ;
        RECT 1877.135 1448.840 1877.650 1448.980 ;
        RECT 1877.330 1448.780 1877.650 1448.840 ;
        RECT 1877.330 1414.100 1877.650 1414.360 ;
        RECT 1877.420 1413.960 1877.560 1414.100 ;
        RECT 1878.250 1413.960 1878.570 1414.020 ;
        RECT 1877.420 1413.820 1878.570 1413.960 ;
        RECT 1878.250 1413.760 1878.570 1413.820 ;
        RECT 1875.950 1400.700 1876.270 1400.760 ;
        RECT 1878.250 1400.700 1878.570 1400.760 ;
        RECT 1875.950 1400.560 1878.570 1400.700 ;
        RECT 1875.950 1400.500 1876.270 1400.560 ;
        RECT 1878.250 1400.500 1878.570 1400.560 ;
        RECT 1875.950 1345.280 1876.270 1345.340 ;
        RECT 1878.250 1345.280 1878.570 1345.340 ;
        RECT 1875.950 1345.140 1878.570 1345.280 ;
        RECT 1875.950 1345.080 1876.270 1345.140 ;
        RECT 1878.250 1345.080 1878.570 1345.140 ;
        RECT 1877.805 1270.140 1878.095 1270.185 ;
        RECT 1878.250 1270.140 1878.570 1270.200 ;
        RECT 1877.805 1270.000 1878.570 1270.140 ;
        RECT 1877.805 1269.955 1878.095 1270.000 ;
        RECT 1878.250 1269.940 1878.570 1270.000 ;
        RECT 1877.790 1242.600 1878.110 1242.660 ;
        RECT 1877.595 1242.460 1878.110 1242.600 ;
        RECT 1877.790 1242.400 1878.110 1242.460 ;
        RECT 1877.790 1241.920 1878.110 1241.980 ;
        RECT 1877.595 1241.780 1878.110 1241.920 ;
        RECT 1877.790 1241.720 1878.110 1241.780 ;
        RECT 1877.790 1214.040 1878.110 1214.100 ;
        RECT 1877.595 1213.900 1878.110 1214.040 ;
        RECT 1877.790 1213.840 1878.110 1213.900 ;
        RECT 1877.330 1104.220 1877.650 1104.280 ;
        RECT 1877.790 1104.220 1878.110 1104.280 ;
        RECT 1877.330 1104.080 1878.110 1104.220 ;
        RECT 1877.330 1104.020 1877.650 1104.080 ;
        RECT 1877.790 1104.020 1878.110 1104.080 ;
        RECT 1877.330 1103.540 1877.650 1103.600 ;
        RECT 1879.170 1103.540 1879.490 1103.600 ;
        RECT 1877.330 1103.400 1879.490 1103.540 ;
        RECT 1877.330 1103.340 1877.650 1103.400 ;
        RECT 1879.170 1103.340 1879.490 1103.400 ;
        RECT 1877.805 980.460 1878.095 980.505 ;
        RECT 1878.250 980.460 1878.570 980.520 ;
        RECT 1877.805 980.320 1878.570 980.460 ;
        RECT 1877.805 980.275 1878.095 980.320 ;
        RECT 1878.250 980.260 1878.570 980.320 ;
        RECT 1877.790 966.180 1878.110 966.240 ;
        RECT 1877.595 966.040 1878.110 966.180 ;
        RECT 1877.790 965.980 1878.110 966.040 ;
        RECT 1877.790 772.720 1878.110 772.780 ;
        RECT 1877.595 772.580 1878.110 772.720 ;
        RECT 1877.790 772.520 1878.110 772.580 ;
        RECT 1877.790 738.040 1878.110 738.100 ;
        RECT 1877.595 737.900 1878.110 738.040 ;
        RECT 1877.790 737.840 1878.110 737.900 ;
        RECT 1877.790 724.440 1878.110 724.500 ;
        RECT 1878.250 724.440 1878.570 724.500 ;
        RECT 1877.790 724.300 1878.570 724.440 ;
        RECT 1877.790 724.240 1878.110 724.300 ;
        RECT 1878.250 724.240 1878.570 724.300 ;
        RECT 1877.790 467.740 1878.110 467.800 ;
        RECT 1877.595 467.600 1878.110 467.740 ;
        RECT 1877.790 467.540 1878.110 467.600 ;
        RECT 1877.805 427.960 1878.095 428.005 ;
        RECT 1878.250 427.960 1878.570 428.020 ;
        RECT 1877.805 427.820 1878.570 427.960 ;
        RECT 1877.805 427.775 1878.095 427.820 ;
        RECT 1878.250 427.760 1878.570 427.820 ;
        RECT 1877.790 379.340 1878.110 379.400 ;
        RECT 1877.595 379.200 1878.110 379.340 ;
        RECT 1877.790 379.140 1878.110 379.200 ;
        RECT 1877.805 331.740 1878.095 331.785 ;
        RECT 1877.420 331.600 1878.095 331.740 ;
        RECT 1877.420 331.105 1877.560 331.600 ;
        RECT 1877.805 331.555 1878.095 331.600 ;
        RECT 1877.345 330.875 1877.635 331.105 ;
        RECT 1877.345 283.120 1877.635 283.165 ;
        RECT 1877.790 283.120 1878.110 283.180 ;
        RECT 1877.345 282.980 1878.110 283.120 ;
        RECT 1877.345 282.935 1877.635 282.980 ;
        RECT 1877.790 282.920 1878.110 282.980 ;
        RECT 1877.790 282.440 1878.110 282.500 ;
        RECT 1877.595 282.300 1878.110 282.440 ;
        RECT 1877.790 282.240 1878.110 282.300 ;
        RECT 1877.805 258.640 1878.095 258.685 ;
        RECT 1878.250 258.640 1878.570 258.700 ;
        RECT 1877.805 258.500 1878.570 258.640 ;
        RECT 1877.805 258.455 1878.095 258.500 ;
        RECT 1878.250 258.440 1878.570 258.500 ;
        RECT 1877.790 179.420 1878.110 179.480 ;
        RECT 1878.710 179.420 1879.030 179.480 ;
        RECT 1877.790 179.280 1879.030 179.420 ;
        RECT 1877.790 179.220 1878.110 179.280 ;
        RECT 1878.710 179.220 1879.030 179.280 ;
        RECT 1877.330 48.520 1877.650 48.580 ;
        RECT 1878.710 48.520 1879.030 48.580 ;
        RECT 1877.330 48.380 1879.030 48.520 ;
        RECT 1877.330 48.320 1877.650 48.380 ;
        RECT 1878.710 48.320 1879.030 48.380 ;
        RECT 1423.770 36.960 1424.090 37.020 ;
        RECT 1877.330 36.960 1877.650 37.020 ;
        RECT 1423.770 36.820 1877.650 36.960 ;
        RECT 1423.770 36.760 1424.090 36.820 ;
        RECT 1877.330 36.760 1877.650 36.820 ;
      LAYER via ;
        RECT 1877.820 1593.960 1878.080 1594.220 ;
        RECT 1878.740 1593.960 1879.000 1594.220 ;
        RECT 1877.360 1490.260 1877.620 1490.520 ;
        RECT 1877.360 1448.780 1877.620 1449.040 ;
        RECT 1877.360 1414.100 1877.620 1414.360 ;
        RECT 1878.280 1413.760 1878.540 1414.020 ;
        RECT 1875.980 1400.500 1876.240 1400.760 ;
        RECT 1878.280 1400.500 1878.540 1400.760 ;
        RECT 1875.980 1345.080 1876.240 1345.340 ;
        RECT 1878.280 1345.080 1878.540 1345.340 ;
        RECT 1878.280 1269.940 1878.540 1270.200 ;
        RECT 1877.820 1242.400 1878.080 1242.660 ;
        RECT 1877.820 1241.720 1878.080 1241.980 ;
        RECT 1877.820 1213.840 1878.080 1214.100 ;
        RECT 1877.360 1104.020 1877.620 1104.280 ;
        RECT 1877.820 1104.020 1878.080 1104.280 ;
        RECT 1877.360 1103.340 1877.620 1103.600 ;
        RECT 1879.200 1103.340 1879.460 1103.600 ;
        RECT 1878.280 980.260 1878.540 980.520 ;
        RECT 1877.820 965.980 1878.080 966.240 ;
        RECT 1877.820 772.520 1878.080 772.780 ;
        RECT 1877.820 737.840 1878.080 738.100 ;
        RECT 1877.820 724.240 1878.080 724.500 ;
        RECT 1878.280 724.240 1878.540 724.500 ;
        RECT 1877.820 467.540 1878.080 467.800 ;
        RECT 1878.280 427.760 1878.540 428.020 ;
        RECT 1877.820 379.140 1878.080 379.400 ;
        RECT 1877.820 282.920 1878.080 283.180 ;
        RECT 1877.820 282.240 1878.080 282.500 ;
        RECT 1878.280 258.440 1878.540 258.700 ;
        RECT 1877.820 179.220 1878.080 179.480 ;
        RECT 1878.740 179.220 1879.000 179.480 ;
        RECT 1877.360 48.320 1877.620 48.580 ;
        RECT 1878.740 48.320 1879.000 48.580 ;
        RECT 1423.800 36.760 1424.060 37.020 ;
        RECT 1877.360 36.760 1877.620 37.020 ;
      LAYER met2 ;
        RECT 1881.420 1700.410 1881.700 1704.000 ;
        RECT 1879.260 1700.270 1881.700 1700.410 ;
        RECT 1879.260 1641.930 1879.400 1700.270 ;
        RECT 1881.420 1700.000 1881.700 1700.270 ;
        RECT 1878.800 1641.790 1879.400 1641.930 ;
        RECT 1878.800 1594.250 1878.940 1641.790 ;
        RECT 1877.820 1593.930 1878.080 1594.250 ;
        RECT 1878.740 1593.930 1879.000 1594.250 ;
        RECT 1877.880 1593.650 1878.020 1593.930 ;
        RECT 1877.880 1593.510 1878.480 1593.650 ;
        RECT 1878.340 1497.090 1878.480 1593.510 ;
        RECT 1877.420 1496.950 1878.480 1497.090 ;
        RECT 1877.420 1490.550 1877.560 1496.950 ;
        RECT 1877.360 1490.230 1877.620 1490.550 ;
        RECT 1877.360 1448.750 1877.620 1449.070 ;
        RECT 1877.420 1414.390 1877.560 1448.750 ;
        RECT 1877.360 1414.070 1877.620 1414.390 ;
        RECT 1878.280 1413.730 1878.540 1414.050 ;
        RECT 1878.340 1400.790 1878.480 1413.730 ;
        RECT 1875.980 1400.470 1876.240 1400.790 ;
        RECT 1878.280 1400.470 1878.540 1400.790 ;
        RECT 1876.040 1345.370 1876.180 1400.470 ;
        RECT 1875.980 1345.050 1876.240 1345.370 ;
        RECT 1878.280 1345.050 1878.540 1345.370 ;
        RECT 1878.340 1338.765 1878.480 1345.050 ;
        RECT 1877.350 1338.395 1877.630 1338.765 ;
        RECT 1878.270 1338.395 1878.550 1338.765 ;
        RECT 1877.420 1290.485 1877.560 1338.395 ;
        RECT 1877.350 1290.115 1877.630 1290.485 ;
        RECT 1878.270 1290.115 1878.550 1290.485 ;
        RECT 1878.340 1270.230 1878.480 1290.115 ;
        RECT 1878.280 1269.910 1878.540 1270.230 ;
        RECT 1877.820 1242.370 1878.080 1242.690 ;
        RECT 1877.880 1242.010 1878.020 1242.370 ;
        RECT 1877.820 1241.690 1878.080 1242.010 ;
        RECT 1877.820 1213.810 1878.080 1214.130 ;
        RECT 1877.880 1104.310 1878.020 1213.810 ;
        RECT 1877.360 1103.990 1877.620 1104.310 ;
        RECT 1877.820 1103.990 1878.080 1104.310 ;
        RECT 1877.420 1103.630 1877.560 1103.990 ;
        RECT 1877.360 1103.310 1877.620 1103.630 ;
        RECT 1879.200 1103.310 1879.460 1103.630 ;
        RECT 1879.260 1055.885 1879.400 1103.310 ;
        RECT 1878.270 1055.515 1878.550 1055.885 ;
        RECT 1879.190 1055.515 1879.470 1055.885 ;
        RECT 1878.340 980.550 1878.480 1055.515 ;
        RECT 1878.280 980.230 1878.540 980.550 ;
        RECT 1877.820 965.950 1878.080 966.270 ;
        RECT 1877.880 931.330 1878.020 965.950 ;
        RECT 1877.880 931.190 1878.480 931.330 ;
        RECT 1878.340 772.890 1878.480 931.190 ;
        RECT 1877.880 772.810 1878.480 772.890 ;
        RECT 1877.820 772.750 1878.480 772.810 ;
        RECT 1877.820 772.490 1878.080 772.750 ;
        RECT 1877.880 772.335 1878.020 772.490 ;
        RECT 1877.820 737.810 1878.080 738.130 ;
        RECT 1877.880 724.610 1878.020 737.810 ;
        RECT 1877.880 724.530 1878.480 724.610 ;
        RECT 1877.820 724.470 1878.540 724.530 ;
        RECT 1877.820 724.210 1878.080 724.470 ;
        RECT 1878.280 724.210 1878.540 724.470 ;
        RECT 1877.880 641.650 1878.020 724.210 ;
        RECT 1877.880 641.510 1878.480 641.650 ;
        RECT 1878.340 497.490 1878.480 641.510 ;
        RECT 1877.880 497.350 1878.480 497.490 ;
        RECT 1877.880 467.830 1878.020 497.350 ;
        RECT 1877.820 467.510 1878.080 467.830 ;
        RECT 1878.280 427.730 1878.540 428.050 ;
        RECT 1878.340 427.450 1878.480 427.730 ;
        RECT 1877.880 427.310 1878.480 427.450 ;
        RECT 1877.880 400.420 1878.020 427.310 ;
        RECT 1877.880 400.280 1878.940 400.420 ;
        RECT 1878.800 379.850 1878.940 400.280 ;
        RECT 1877.880 379.710 1878.940 379.850 ;
        RECT 1877.880 379.430 1878.020 379.710 ;
        RECT 1877.820 379.110 1878.080 379.430 ;
        RECT 1877.820 282.890 1878.080 283.210 ;
        RECT 1877.880 282.530 1878.020 282.890 ;
        RECT 1877.820 282.210 1878.080 282.530 ;
        RECT 1878.280 258.410 1878.540 258.730 ;
        RECT 1878.340 179.930 1878.480 258.410 ;
        RECT 1877.880 179.790 1878.480 179.930 ;
        RECT 1877.880 179.510 1878.020 179.790 ;
        RECT 1877.820 179.190 1878.080 179.510 ;
        RECT 1878.740 179.190 1879.000 179.510 ;
        RECT 1878.800 48.610 1878.940 179.190 ;
        RECT 1877.360 48.290 1877.620 48.610 ;
        RECT 1878.740 48.290 1879.000 48.610 ;
        RECT 1877.420 37.050 1877.560 48.290 ;
        RECT 1423.800 36.730 1424.060 37.050 ;
        RECT 1877.360 36.730 1877.620 37.050 ;
        RECT 1423.860 2.400 1424.000 36.730 ;
        RECT 1423.650 -4.800 1424.210 2.400 ;
      LAYER via2 ;
        RECT 1877.350 1338.440 1877.630 1338.720 ;
        RECT 1878.270 1338.440 1878.550 1338.720 ;
        RECT 1877.350 1290.160 1877.630 1290.440 ;
        RECT 1878.270 1290.160 1878.550 1290.440 ;
        RECT 1878.270 1055.560 1878.550 1055.840 ;
        RECT 1879.190 1055.560 1879.470 1055.840 ;
      LAYER met3 ;
        RECT 1877.325 1338.730 1877.655 1338.745 ;
        RECT 1878.245 1338.730 1878.575 1338.745 ;
        RECT 1877.325 1338.430 1878.575 1338.730 ;
        RECT 1877.325 1338.415 1877.655 1338.430 ;
        RECT 1878.245 1338.415 1878.575 1338.430 ;
        RECT 1877.325 1290.450 1877.655 1290.465 ;
        RECT 1878.245 1290.450 1878.575 1290.465 ;
        RECT 1877.325 1290.150 1878.575 1290.450 ;
        RECT 1877.325 1290.135 1877.655 1290.150 ;
        RECT 1878.245 1290.135 1878.575 1290.150 ;
        RECT 1878.245 1055.850 1878.575 1055.865 ;
        RECT 1879.165 1055.850 1879.495 1055.865 ;
        RECT 1878.245 1055.550 1879.495 1055.850 ;
        RECT 1878.245 1055.535 1878.575 1055.550 ;
        RECT 1879.165 1055.535 1879.495 1055.550 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1464.710 51.580 1465.030 51.640 ;
        RECT 1891.590 51.580 1891.910 51.640 ;
        RECT 1464.710 51.440 1891.910 51.580 ;
        RECT 1464.710 51.380 1465.030 51.440 ;
        RECT 1891.590 51.380 1891.910 51.440 ;
        RECT 1441.710 16.220 1442.030 16.280 ;
        RECT 1464.710 16.220 1465.030 16.280 ;
        RECT 1441.710 16.080 1465.030 16.220 ;
        RECT 1441.710 16.020 1442.030 16.080 ;
        RECT 1464.710 16.020 1465.030 16.080 ;
      LAYER via ;
        RECT 1464.740 51.380 1465.000 51.640 ;
        RECT 1891.620 51.380 1891.880 51.640 ;
        RECT 1441.740 16.020 1442.000 16.280 ;
        RECT 1464.740 16.020 1465.000 16.280 ;
      LAYER met2 ;
        RECT 1890.620 1700.410 1890.900 1704.000 ;
        RECT 1890.620 1700.270 1891.820 1700.410 ;
        RECT 1890.620 1700.000 1890.900 1700.270 ;
        RECT 1891.680 51.670 1891.820 1700.270 ;
        RECT 1464.740 51.350 1465.000 51.670 ;
        RECT 1891.620 51.350 1891.880 51.670 ;
        RECT 1464.800 16.310 1464.940 51.350 ;
        RECT 1441.740 15.990 1442.000 16.310 ;
        RECT 1464.740 15.990 1465.000 16.310 ;
        RECT 1441.800 2.400 1441.940 15.990 ;
        RECT 1441.590 -4.800 1442.150 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1498.290 52.260 1498.610 52.320 ;
        RECT 1898.030 52.260 1898.350 52.320 ;
        RECT 1498.290 52.120 1898.350 52.260 ;
        RECT 1498.290 52.060 1498.610 52.120 ;
        RECT 1898.030 52.060 1898.350 52.120 ;
        RECT 1459.650 18.260 1459.970 18.320 ;
        RECT 1498.290 18.260 1498.610 18.320 ;
        RECT 1459.650 18.120 1498.610 18.260 ;
        RECT 1459.650 18.060 1459.970 18.120 ;
        RECT 1498.290 18.060 1498.610 18.120 ;
      LAYER via ;
        RECT 1498.320 52.060 1498.580 52.320 ;
        RECT 1898.060 52.060 1898.320 52.320 ;
        RECT 1459.680 18.060 1459.940 18.320 ;
        RECT 1498.320 18.060 1498.580 18.320 ;
      LAYER met2 ;
        RECT 1899.820 1700.410 1900.100 1704.000 ;
        RECT 1898.120 1700.270 1900.100 1700.410 ;
        RECT 1898.120 52.350 1898.260 1700.270 ;
        RECT 1899.820 1700.000 1900.100 1700.270 ;
        RECT 1498.320 52.030 1498.580 52.350 ;
        RECT 1898.060 52.030 1898.320 52.350 ;
        RECT 1498.380 18.350 1498.520 52.030 ;
        RECT 1459.680 18.030 1459.940 18.350 ;
        RECT 1498.320 18.030 1498.580 18.350 ;
        RECT 1459.740 2.400 1459.880 18.030 ;
        RECT 1459.530 -4.800 1460.090 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1905.925 1642.285 1906.095 1655.715 ;
        RECT 1905.465 1352.605 1905.635 1400.375 ;
        RECT 1905.465 1304.325 1905.635 1352.095 ;
        RECT 1905.465 737.885 1905.635 772.735 ;
        RECT 1905.465 676.345 1905.635 724.115 ;
        RECT 1905.925 579.785 1906.095 627.895 ;
        RECT 1905.005 434.945 1905.175 449.055 ;
        RECT 1905.005 379.525 1905.175 427.635 ;
        RECT 1905.465 289.765 1905.635 337.875 ;
      LAYER mcon ;
        RECT 1905.925 1655.545 1906.095 1655.715 ;
        RECT 1905.465 1400.205 1905.635 1400.375 ;
        RECT 1905.465 1351.925 1905.635 1352.095 ;
        RECT 1905.465 772.565 1905.635 772.735 ;
        RECT 1905.465 723.945 1905.635 724.115 ;
        RECT 1905.925 627.725 1906.095 627.895 ;
        RECT 1905.005 448.885 1905.175 449.055 ;
        RECT 1905.005 427.465 1905.175 427.635 ;
        RECT 1905.465 337.705 1905.635 337.875 ;
      LAYER met1 ;
        RECT 1905.850 1655.700 1906.170 1655.760 ;
        RECT 1905.655 1655.560 1906.170 1655.700 ;
        RECT 1905.850 1655.500 1906.170 1655.560 ;
        RECT 1905.390 1642.440 1905.710 1642.500 ;
        RECT 1905.865 1642.440 1906.155 1642.485 ;
        RECT 1905.390 1642.300 1906.155 1642.440 ;
        RECT 1905.390 1642.240 1905.710 1642.300 ;
        RECT 1905.865 1642.255 1906.155 1642.300 ;
        RECT 1905.390 1587.020 1905.710 1587.080 ;
        RECT 1906.770 1587.020 1907.090 1587.080 ;
        RECT 1905.390 1586.880 1907.090 1587.020 ;
        RECT 1905.390 1586.820 1905.710 1586.880 ;
        RECT 1906.770 1586.820 1907.090 1586.880 ;
        RECT 1905.390 1449.320 1905.710 1449.380 ;
        RECT 1906.770 1449.320 1907.090 1449.380 ;
        RECT 1905.390 1449.180 1907.090 1449.320 ;
        RECT 1905.390 1449.120 1905.710 1449.180 ;
        RECT 1906.770 1449.120 1907.090 1449.180 ;
        RECT 1905.390 1414.440 1905.710 1414.700 ;
        RECT 1905.480 1413.960 1905.620 1414.440 ;
        RECT 1905.850 1413.960 1906.170 1414.020 ;
        RECT 1905.480 1413.820 1906.170 1413.960 ;
        RECT 1905.850 1413.760 1906.170 1413.820 ;
        RECT 1905.405 1400.360 1905.695 1400.405 ;
        RECT 1905.850 1400.360 1906.170 1400.420 ;
        RECT 1905.405 1400.220 1906.170 1400.360 ;
        RECT 1905.405 1400.175 1905.695 1400.220 ;
        RECT 1905.850 1400.160 1906.170 1400.220 ;
        RECT 1905.390 1352.760 1905.710 1352.820 ;
        RECT 1905.195 1352.620 1905.710 1352.760 ;
        RECT 1905.390 1352.560 1905.710 1352.620 ;
        RECT 1905.390 1352.080 1905.710 1352.140 ;
        RECT 1905.195 1351.940 1905.710 1352.080 ;
        RECT 1905.390 1351.880 1905.710 1351.940 ;
        RECT 1905.405 1304.480 1905.695 1304.525 ;
        RECT 1905.850 1304.480 1906.170 1304.540 ;
        RECT 1905.405 1304.340 1906.170 1304.480 ;
        RECT 1905.405 1304.295 1905.695 1304.340 ;
        RECT 1905.850 1304.280 1906.170 1304.340 ;
        RECT 1906.310 1256.540 1906.630 1256.600 ;
        RECT 1905.480 1256.400 1906.630 1256.540 ;
        RECT 1905.480 1256.260 1905.620 1256.400 ;
        RECT 1906.310 1256.340 1906.630 1256.400 ;
        RECT 1905.390 1256.000 1905.710 1256.260 ;
        RECT 1905.390 1221.320 1905.710 1221.580 ;
        RECT 1905.480 1220.840 1905.620 1221.320 ;
        RECT 1905.850 1220.840 1906.170 1220.900 ;
        RECT 1905.480 1220.700 1906.170 1220.840 ;
        RECT 1905.850 1220.640 1906.170 1220.700 ;
        RECT 1905.850 1173.240 1906.170 1173.300 ;
        RECT 1905.480 1173.100 1906.170 1173.240 ;
        RECT 1905.480 1172.960 1905.620 1173.100 ;
        RECT 1905.850 1173.040 1906.170 1173.100 ;
        RECT 1905.390 1172.700 1905.710 1172.960 ;
        RECT 1905.390 1124.760 1905.710 1125.020 ;
        RECT 1905.480 1124.280 1905.620 1124.760 ;
        RECT 1905.850 1124.280 1906.170 1124.340 ;
        RECT 1905.480 1124.140 1906.170 1124.280 ;
        RECT 1905.850 1124.080 1906.170 1124.140 ;
        RECT 1905.390 772.720 1905.710 772.780 ;
        RECT 1905.195 772.580 1905.710 772.720 ;
        RECT 1905.390 772.520 1905.710 772.580 ;
        RECT 1905.390 738.040 1905.710 738.100 ;
        RECT 1905.195 737.900 1905.710 738.040 ;
        RECT 1905.390 737.840 1905.710 737.900 ;
        RECT 1905.405 724.100 1905.695 724.145 ;
        RECT 1905.850 724.100 1906.170 724.160 ;
        RECT 1905.405 723.960 1906.170 724.100 ;
        RECT 1905.405 723.915 1905.695 723.960 ;
        RECT 1905.850 723.900 1906.170 723.960 ;
        RECT 1905.390 676.500 1905.710 676.560 ;
        RECT 1905.195 676.360 1905.710 676.500 ;
        RECT 1905.390 676.300 1905.710 676.360 ;
        RECT 1905.850 627.880 1906.170 627.940 ;
        RECT 1905.655 627.740 1906.170 627.880 ;
        RECT 1905.850 627.680 1906.170 627.740 ;
        RECT 1905.850 579.940 1906.170 580.000 ;
        RECT 1905.655 579.800 1906.170 579.940 ;
        RECT 1905.850 579.740 1906.170 579.800 ;
        RECT 1904.945 449.040 1905.235 449.085 ;
        RECT 1905.390 449.040 1905.710 449.100 ;
        RECT 1904.945 448.900 1905.710 449.040 ;
        RECT 1904.945 448.855 1905.235 448.900 ;
        RECT 1905.390 448.840 1905.710 448.900 ;
        RECT 1904.930 435.100 1905.250 435.160 ;
        RECT 1904.735 434.960 1905.250 435.100 ;
        RECT 1904.930 434.900 1905.250 434.960 ;
        RECT 1904.930 427.620 1905.250 427.680 ;
        RECT 1904.735 427.480 1905.250 427.620 ;
        RECT 1904.930 427.420 1905.250 427.480 ;
        RECT 1904.945 379.680 1905.235 379.725 ;
        RECT 1905.390 379.680 1905.710 379.740 ;
        RECT 1904.945 379.540 1905.710 379.680 ;
        RECT 1904.945 379.495 1905.235 379.540 ;
        RECT 1905.390 379.480 1905.710 379.540 ;
        RECT 1905.390 337.860 1905.710 337.920 ;
        RECT 1905.195 337.720 1905.710 337.860 ;
        RECT 1905.390 337.660 1905.710 337.720 ;
        RECT 1905.390 289.920 1905.710 289.980 ;
        RECT 1905.195 289.780 1905.710 289.920 ;
        RECT 1905.390 289.720 1905.710 289.780 ;
        RECT 1904.930 241.300 1905.250 241.360 ;
        RECT 1905.850 241.300 1906.170 241.360 ;
        RECT 1904.930 241.160 1906.170 241.300 ;
        RECT 1904.930 241.100 1905.250 241.160 ;
        RECT 1905.850 241.100 1906.170 241.160 ;
        RECT 1905.390 145.080 1905.710 145.140 ;
        RECT 1905.850 145.080 1906.170 145.140 ;
        RECT 1905.390 144.940 1906.170 145.080 ;
        RECT 1905.390 144.880 1905.710 144.940 ;
        RECT 1905.850 144.880 1906.170 144.940 ;
        RECT 1904.010 111.080 1904.330 111.140 ;
        RECT 1905.850 111.080 1906.170 111.140 ;
        RECT 1904.010 110.940 1906.170 111.080 ;
        RECT 1904.010 110.880 1904.330 110.940 ;
        RECT 1905.850 110.880 1906.170 110.940 ;
        RECT 1593.970 33.560 1594.290 33.620 ;
        RECT 1904.010 33.560 1904.330 33.620 ;
        RECT 1593.970 33.420 1904.330 33.560 ;
        RECT 1593.970 33.360 1594.290 33.420 ;
        RECT 1904.010 33.360 1904.330 33.420 ;
        RECT 1477.590 16.900 1477.910 16.960 ;
        RECT 1593.970 16.900 1594.290 16.960 ;
        RECT 1477.590 16.760 1594.290 16.900 ;
        RECT 1477.590 16.700 1477.910 16.760 ;
        RECT 1593.970 16.700 1594.290 16.760 ;
      LAYER via ;
        RECT 1905.880 1655.500 1906.140 1655.760 ;
        RECT 1905.420 1642.240 1905.680 1642.500 ;
        RECT 1905.420 1586.820 1905.680 1587.080 ;
        RECT 1906.800 1586.820 1907.060 1587.080 ;
        RECT 1905.420 1449.120 1905.680 1449.380 ;
        RECT 1906.800 1449.120 1907.060 1449.380 ;
        RECT 1905.420 1414.440 1905.680 1414.700 ;
        RECT 1905.880 1413.760 1906.140 1414.020 ;
        RECT 1905.880 1400.160 1906.140 1400.420 ;
        RECT 1905.420 1352.560 1905.680 1352.820 ;
        RECT 1905.420 1351.880 1905.680 1352.140 ;
        RECT 1905.880 1304.280 1906.140 1304.540 ;
        RECT 1906.340 1256.340 1906.600 1256.600 ;
        RECT 1905.420 1256.000 1905.680 1256.260 ;
        RECT 1905.420 1221.320 1905.680 1221.580 ;
        RECT 1905.880 1220.640 1906.140 1220.900 ;
        RECT 1905.880 1173.040 1906.140 1173.300 ;
        RECT 1905.420 1172.700 1905.680 1172.960 ;
        RECT 1905.420 1124.760 1905.680 1125.020 ;
        RECT 1905.880 1124.080 1906.140 1124.340 ;
        RECT 1905.420 772.520 1905.680 772.780 ;
        RECT 1905.420 737.840 1905.680 738.100 ;
        RECT 1905.880 723.900 1906.140 724.160 ;
        RECT 1905.420 676.300 1905.680 676.560 ;
        RECT 1905.880 627.680 1906.140 627.940 ;
        RECT 1905.880 579.740 1906.140 580.000 ;
        RECT 1905.420 448.840 1905.680 449.100 ;
        RECT 1904.960 434.900 1905.220 435.160 ;
        RECT 1904.960 427.420 1905.220 427.680 ;
        RECT 1905.420 379.480 1905.680 379.740 ;
        RECT 1905.420 337.660 1905.680 337.920 ;
        RECT 1905.420 289.720 1905.680 289.980 ;
        RECT 1904.960 241.100 1905.220 241.360 ;
        RECT 1905.880 241.100 1906.140 241.360 ;
        RECT 1905.420 144.880 1905.680 145.140 ;
        RECT 1905.880 144.880 1906.140 145.140 ;
        RECT 1904.040 110.880 1904.300 111.140 ;
        RECT 1905.880 110.880 1906.140 111.140 ;
        RECT 1594.000 33.360 1594.260 33.620 ;
        RECT 1904.040 33.360 1904.300 33.620 ;
        RECT 1477.620 16.700 1477.880 16.960 ;
        RECT 1594.000 16.700 1594.260 16.960 ;
      LAYER met2 ;
        RECT 1909.020 1701.090 1909.300 1704.000 ;
        RECT 1906.400 1700.950 1909.300 1701.090 ;
        RECT 1906.400 1690.210 1906.540 1700.950 ;
        RECT 1909.020 1700.000 1909.300 1700.950 ;
        RECT 1905.940 1690.070 1906.540 1690.210 ;
        RECT 1905.940 1655.790 1906.080 1690.070 ;
        RECT 1905.880 1655.470 1906.140 1655.790 ;
        RECT 1905.420 1642.440 1905.680 1642.530 ;
        RECT 1905.420 1642.300 1906.080 1642.440 ;
        RECT 1905.420 1642.210 1905.680 1642.300 ;
        RECT 1905.940 1595.125 1906.080 1642.300 ;
        RECT 1905.870 1594.755 1906.150 1595.125 ;
        RECT 1905.410 1594.075 1905.690 1594.445 ;
        RECT 1905.480 1587.110 1905.620 1594.075 ;
        RECT 1905.420 1586.790 1905.680 1587.110 ;
        RECT 1906.800 1586.790 1907.060 1587.110 ;
        RECT 1906.860 1449.410 1907.000 1586.790 ;
        RECT 1905.420 1449.090 1905.680 1449.410 ;
        RECT 1906.800 1449.090 1907.060 1449.410 ;
        RECT 1905.480 1414.730 1905.620 1449.090 ;
        RECT 1905.420 1414.410 1905.680 1414.730 ;
        RECT 1905.880 1413.730 1906.140 1414.050 ;
        RECT 1905.940 1400.450 1906.080 1413.730 ;
        RECT 1905.880 1400.130 1906.140 1400.450 ;
        RECT 1905.420 1352.530 1905.680 1352.850 ;
        RECT 1905.480 1352.170 1905.620 1352.530 ;
        RECT 1905.420 1351.850 1905.680 1352.170 ;
        RECT 1905.880 1304.250 1906.140 1304.570 ;
        RECT 1905.940 1303.970 1906.080 1304.250 ;
        RECT 1905.940 1303.830 1906.540 1303.970 ;
        RECT 1906.400 1256.630 1906.540 1303.830 ;
        RECT 1906.340 1256.310 1906.600 1256.630 ;
        RECT 1905.420 1255.970 1905.680 1256.290 ;
        RECT 1905.480 1221.610 1905.620 1255.970 ;
        RECT 1905.420 1221.290 1905.680 1221.610 ;
        RECT 1905.880 1220.610 1906.140 1220.930 ;
        RECT 1905.940 1207.410 1906.080 1220.610 ;
        RECT 1905.480 1207.270 1906.080 1207.410 ;
        RECT 1905.480 1200.610 1905.620 1207.270 ;
        RECT 1905.480 1200.470 1906.080 1200.610 ;
        RECT 1905.940 1173.330 1906.080 1200.470 ;
        RECT 1905.880 1173.010 1906.140 1173.330 ;
        RECT 1905.420 1172.670 1905.680 1172.990 ;
        RECT 1905.480 1125.050 1905.620 1172.670 ;
        RECT 1905.420 1124.730 1905.680 1125.050 ;
        RECT 1905.880 1124.050 1906.140 1124.370 ;
        RECT 1905.940 1110.850 1906.080 1124.050 ;
        RECT 1905.480 1110.710 1906.080 1110.850 ;
        RECT 1905.480 1104.165 1905.620 1110.710 ;
        RECT 1904.030 1103.795 1904.310 1104.165 ;
        RECT 1905.410 1103.795 1905.690 1104.165 ;
        RECT 1904.100 1055.885 1904.240 1103.795 ;
        RECT 1904.030 1055.515 1904.310 1055.885 ;
        RECT 1904.950 1055.515 1905.230 1055.885 ;
        RECT 1905.020 1027.890 1905.160 1055.515 ;
        RECT 1905.020 1027.750 1906.080 1027.890 ;
        RECT 1905.940 1014.290 1906.080 1027.750 ;
        RECT 1905.480 1014.150 1906.080 1014.290 ;
        RECT 1905.480 931.330 1905.620 1014.150 ;
        RECT 1905.480 931.190 1906.080 931.330 ;
        RECT 1905.940 772.890 1906.080 931.190 ;
        RECT 1905.480 772.810 1906.080 772.890 ;
        RECT 1905.420 772.750 1906.080 772.810 ;
        RECT 1905.420 772.490 1905.680 772.750 ;
        RECT 1905.480 772.335 1905.620 772.490 ;
        RECT 1905.420 737.810 1905.680 738.130 ;
        RECT 1905.480 724.610 1905.620 737.810 ;
        RECT 1905.480 724.470 1906.080 724.610 ;
        RECT 1905.940 724.190 1906.080 724.470 ;
        RECT 1905.880 723.870 1906.140 724.190 ;
        RECT 1905.420 676.270 1905.680 676.590 ;
        RECT 1905.480 641.650 1905.620 676.270 ;
        RECT 1905.480 641.510 1906.080 641.650 ;
        RECT 1905.940 627.970 1906.080 641.510 ;
        RECT 1905.880 627.650 1906.140 627.970 ;
        RECT 1905.880 579.710 1906.140 580.030 ;
        RECT 1905.940 497.490 1906.080 579.710 ;
        RECT 1905.480 497.350 1906.080 497.490 ;
        RECT 1905.480 449.130 1905.620 497.350 ;
        RECT 1905.420 448.810 1905.680 449.130 ;
        RECT 1904.960 434.870 1905.220 435.190 ;
        RECT 1905.020 427.710 1905.160 434.870 ;
        RECT 1904.960 427.390 1905.220 427.710 ;
        RECT 1905.420 379.450 1905.680 379.770 ;
        RECT 1905.480 337.950 1905.620 379.450 ;
        RECT 1905.420 337.630 1905.680 337.950 ;
        RECT 1905.420 289.690 1905.680 290.010 ;
        RECT 1905.480 265.610 1905.620 289.690 ;
        RECT 1905.480 265.470 1906.540 265.610 ;
        RECT 1906.400 254.730 1906.540 265.470 ;
        RECT 1905.940 254.590 1906.540 254.730 ;
        RECT 1905.940 241.390 1906.080 254.590 ;
        RECT 1904.960 241.070 1905.220 241.390 ;
        RECT 1905.880 241.070 1906.140 241.390 ;
        RECT 1905.020 206.450 1905.160 241.070 ;
        RECT 1905.020 206.310 1905.620 206.450 ;
        RECT 1905.480 145.170 1905.620 206.310 ;
        RECT 1905.420 144.850 1905.680 145.170 ;
        RECT 1905.880 144.850 1906.140 145.170 ;
        RECT 1905.940 111.170 1906.080 144.850 ;
        RECT 1904.040 110.850 1904.300 111.170 ;
        RECT 1905.880 110.850 1906.140 111.170 ;
        RECT 1904.100 33.650 1904.240 110.850 ;
        RECT 1594.000 33.330 1594.260 33.650 ;
        RECT 1904.040 33.330 1904.300 33.650 ;
        RECT 1594.060 16.990 1594.200 33.330 ;
        RECT 1477.620 16.670 1477.880 16.990 ;
        RECT 1594.000 16.670 1594.260 16.990 ;
        RECT 1477.680 2.400 1477.820 16.670 ;
        RECT 1477.470 -4.800 1478.030 2.400 ;
      LAYER via2 ;
        RECT 1905.870 1594.800 1906.150 1595.080 ;
        RECT 1905.410 1594.120 1905.690 1594.400 ;
        RECT 1904.030 1103.840 1904.310 1104.120 ;
        RECT 1905.410 1103.840 1905.690 1104.120 ;
        RECT 1904.030 1055.560 1904.310 1055.840 ;
        RECT 1904.950 1055.560 1905.230 1055.840 ;
      LAYER met3 ;
        RECT 1905.845 1595.090 1906.175 1595.105 ;
        RECT 1904.710 1594.790 1906.175 1595.090 ;
        RECT 1904.710 1594.410 1905.010 1594.790 ;
        RECT 1905.845 1594.775 1906.175 1594.790 ;
        RECT 1905.385 1594.410 1905.715 1594.425 ;
        RECT 1904.710 1594.110 1905.715 1594.410 ;
        RECT 1905.385 1594.095 1905.715 1594.110 ;
        RECT 1904.005 1104.130 1904.335 1104.145 ;
        RECT 1905.385 1104.130 1905.715 1104.145 ;
        RECT 1904.005 1103.830 1905.715 1104.130 ;
        RECT 1904.005 1103.815 1904.335 1103.830 ;
        RECT 1905.385 1103.815 1905.715 1103.830 ;
        RECT 1904.005 1055.850 1904.335 1055.865 ;
        RECT 1904.925 1055.850 1905.255 1055.865 ;
        RECT 1904.005 1055.550 1905.255 1055.850 ;
        RECT 1904.005 1055.535 1904.335 1055.550 ;
        RECT 1904.925 1055.535 1905.255 1055.550 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1504.730 51.920 1505.050 51.980 ;
        RECT 1918.730 51.920 1919.050 51.980 ;
        RECT 1504.730 51.780 1919.050 51.920 ;
        RECT 1504.730 51.720 1505.050 51.780 ;
        RECT 1918.730 51.720 1919.050 51.780 ;
        RECT 1495.530 18.600 1495.850 18.660 ;
        RECT 1504.730 18.600 1505.050 18.660 ;
        RECT 1495.530 18.460 1505.050 18.600 ;
        RECT 1495.530 18.400 1495.850 18.460 ;
        RECT 1504.730 18.400 1505.050 18.460 ;
      LAYER via ;
        RECT 1504.760 51.720 1505.020 51.980 ;
        RECT 1918.760 51.720 1919.020 51.980 ;
        RECT 1495.560 18.400 1495.820 18.660 ;
        RECT 1504.760 18.400 1505.020 18.660 ;
      LAYER met2 ;
        RECT 1918.220 1700.410 1918.500 1704.000 ;
        RECT 1918.220 1700.270 1918.960 1700.410 ;
        RECT 1918.220 1700.000 1918.500 1700.270 ;
        RECT 1918.820 52.010 1918.960 1700.270 ;
        RECT 1504.760 51.690 1505.020 52.010 ;
        RECT 1918.760 51.690 1919.020 52.010 ;
        RECT 1504.820 18.690 1504.960 51.690 ;
        RECT 1495.560 18.370 1495.820 18.690 ;
        RECT 1504.760 18.370 1505.020 18.690 ;
        RECT 1495.620 2.400 1495.760 18.370 ;
        RECT 1495.410 -4.800 1495.970 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1600.870 33.220 1601.190 33.280 ;
        RECT 1925.630 33.220 1925.950 33.280 ;
        RECT 1600.870 33.080 1925.950 33.220 ;
        RECT 1600.870 33.020 1601.190 33.080 ;
        RECT 1925.630 33.020 1925.950 33.080 ;
        RECT 1513.010 16.220 1513.330 16.280 ;
        RECT 1600.870 16.220 1601.190 16.280 ;
        RECT 1513.010 16.080 1601.190 16.220 ;
        RECT 1513.010 16.020 1513.330 16.080 ;
        RECT 1600.870 16.020 1601.190 16.080 ;
      LAYER via ;
        RECT 1600.900 33.020 1601.160 33.280 ;
        RECT 1925.660 33.020 1925.920 33.280 ;
        RECT 1513.040 16.020 1513.300 16.280 ;
        RECT 1600.900 16.020 1601.160 16.280 ;
      LAYER met2 ;
        RECT 1927.420 1700.410 1927.700 1704.000 ;
        RECT 1925.720 1700.270 1927.700 1700.410 ;
        RECT 1925.720 33.310 1925.860 1700.270 ;
        RECT 1927.420 1700.000 1927.700 1700.270 ;
        RECT 1600.900 32.990 1601.160 33.310 ;
        RECT 1925.660 32.990 1925.920 33.310 ;
        RECT 1600.960 16.310 1601.100 32.990 ;
        RECT 1513.040 15.990 1513.300 16.310 ;
        RECT 1600.900 15.990 1601.160 16.310 ;
        RECT 1513.100 2.400 1513.240 15.990 ;
        RECT 1512.890 -4.800 1513.450 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 709.850 36.280 710.170 36.340 ;
        RECT 1512.550 36.280 1512.870 36.340 ;
        RECT 709.850 36.140 1512.870 36.280 ;
        RECT 709.850 36.080 710.170 36.140 ;
        RECT 1512.550 36.080 1512.870 36.140 ;
      LAYER via ;
        RECT 709.880 36.080 710.140 36.340 ;
        RECT 1512.580 36.080 1512.840 36.340 ;
      LAYER met2 ;
        RECT 1513.880 1700.410 1514.160 1704.000 ;
        RECT 1512.640 1700.270 1514.160 1700.410 ;
        RECT 1512.640 36.370 1512.780 1700.270 ;
        RECT 1513.880 1700.000 1514.160 1700.270 ;
        RECT 709.880 36.050 710.140 36.370 ;
        RECT 1512.580 36.050 1512.840 36.370 ;
        RECT 709.940 17.410 710.080 36.050 ;
        RECT 709.940 17.270 710.540 17.410 ;
        RECT 710.400 2.400 710.540 17.270 ;
        RECT 710.190 -4.800 710.750 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1933.525 1545.725 1933.695 1593.835 ;
        RECT 1933.065 1393.745 1933.235 1435.395 ;
        RECT 1933.065 1345.805 1933.235 1366.375 ;
        RECT 1932.605 1297.185 1932.775 1321.495 ;
        RECT 1933.065 931.345 1933.235 993.395 ;
        RECT 1933.065 614.465 1933.235 669.375 ;
        RECT 1934.445 517.565 1934.615 607.155 ;
      LAYER mcon ;
        RECT 1933.525 1593.665 1933.695 1593.835 ;
        RECT 1933.065 1435.225 1933.235 1435.395 ;
        RECT 1933.065 1366.205 1933.235 1366.375 ;
        RECT 1932.605 1321.325 1932.775 1321.495 ;
        RECT 1933.065 993.225 1933.235 993.395 ;
        RECT 1933.065 669.205 1933.235 669.375 ;
        RECT 1934.445 606.985 1934.615 607.155 ;
      LAYER met1 ;
        RECT 1933.450 1642.440 1933.770 1642.500 ;
        RECT 1934.370 1642.440 1934.690 1642.500 ;
        RECT 1933.450 1642.300 1934.690 1642.440 ;
        RECT 1933.450 1642.240 1933.770 1642.300 ;
        RECT 1934.370 1642.240 1934.690 1642.300 ;
        RECT 1933.450 1593.820 1933.770 1593.880 ;
        RECT 1933.255 1593.680 1933.770 1593.820 ;
        RECT 1933.450 1593.620 1933.770 1593.680 ;
        RECT 1933.450 1545.880 1933.770 1545.940 ;
        RECT 1933.255 1545.740 1933.770 1545.880 ;
        RECT 1933.450 1545.680 1933.770 1545.740 ;
        RECT 1932.990 1435.380 1933.310 1435.440 ;
        RECT 1932.795 1435.240 1933.310 1435.380 ;
        RECT 1932.990 1435.180 1933.310 1435.240 ;
        RECT 1933.005 1393.900 1933.295 1393.945 ;
        RECT 1933.450 1393.900 1933.770 1393.960 ;
        RECT 1933.005 1393.760 1933.770 1393.900 ;
        RECT 1933.005 1393.715 1933.295 1393.760 ;
        RECT 1933.450 1393.700 1933.770 1393.760 ;
        RECT 1932.990 1366.360 1933.310 1366.420 ;
        RECT 1932.795 1366.220 1933.310 1366.360 ;
        RECT 1932.990 1366.160 1933.310 1366.220 ;
        RECT 1932.990 1345.960 1933.310 1346.020 ;
        RECT 1932.795 1345.820 1933.310 1345.960 ;
        RECT 1932.990 1345.760 1933.310 1345.820 ;
        RECT 1932.545 1321.480 1932.835 1321.525 ;
        RECT 1932.990 1321.480 1933.310 1321.540 ;
        RECT 1932.545 1321.340 1933.310 1321.480 ;
        RECT 1932.545 1321.295 1932.835 1321.340 ;
        RECT 1932.990 1321.280 1933.310 1321.340 ;
        RECT 1932.530 1297.340 1932.850 1297.400 ;
        RECT 1932.335 1297.200 1932.850 1297.340 ;
        RECT 1932.530 1297.140 1932.850 1297.200 ;
        RECT 1932.530 1255.860 1932.850 1255.920 ;
        RECT 1934.370 1255.860 1934.690 1255.920 ;
        RECT 1932.530 1255.720 1934.690 1255.860 ;
        RECT 1932.530 1255.660 1932.850 1255.720 ;
        RECT 1934.370 1255.660 1934.690 1255.720 ;
        RECT 1932.990 1159.300 1933.310 1159.360 ;
        RECT 1934.370 1159.300 1934.690 1159.360 ;
        RECT 1932.990 1159.160 1934.690 1159.300 ;
        RECT 1932.990 1159.100 1933.310 1159.160 ;
        RECT 1934.370 1159.100 1934.690 1159.160 ;
        RECT 1932.990 1062.740 1933.310 1062.800 ;
        RECT 1934.370 1062.740 1934.690 1062.800 ;
        RECT 1932.990 1062.600 1934.690 1062.740 ;
        RECT 1932.990 1062.540 1933.310 1062.600 ;
        RECT 1934.370 1062.540 1934.690 1062.600 ;
        RECT 1932.990 1048.800 1933.310 1048.860 ;
        RECT 1933.910 1048.800 1934.230 1048.860 ;
        RECT 1932.990 1048.660 1934.230 1048.800 ;
        RECT 1932.990 1048.600 1933.310 1048.660 ;
        RECT 1933.910 1048.600 1934.230 1048.660 ;
        RECT 1932.990 1000.520 1933.310 1000.580 ;
        RECT 1934.370 1000.520 1934.690 1000.580 ;
        RECT 1932.990 1000.380 1934.690 1000.520 ;
        RECT 1932.990 1000.320 1933.310 1000.380 ;
        RECT 1934.370 1000.320 1934.690 1000.380 ;
        RECT 1932.990 993.380 1933.310 993.440 ;
        RECT 1932.795 993.240 1933.310 993.380 ;
        RECT 1932.990 993.180 1933.310 993.240 ;
        RECT 1932.990 931.500 1933.310 931.560 ;
        RECT 1932.795 931.360 1933.310 931.500 ;
        RECT 1932.990 931.300 1933.310 931.360 ;
        RECT 1933.450 883.700 1933.770 883.960 ;
        RECT 1933.540 883.280 1933.680 883.700 ;
        RECT 1933.450 883.020 1933.770 883.280 ;
        RECT 1933.450 821.000 1933.770 821.060 ;
        RECT 1933.910 821.000 1934.230 821.060 ;
        RECT 1933.450 820.860 1934.230 821.000 ;
        RECT 1933.450 820.800 1933.770 820.860 ;
        RECT 1933.910 820.800 1934.230 820.860 ;
        RECT 1932.990 772.720 1933.310 772.780 ;
        RECT 1933.910 772.720 1934.230 772.780 ;
        RECT 1932.990 772.580 1934.230 772.720 ;
        RECT 1932.990 772.520 1933.310 772.580 ;
        RECT 1933.910 772.520 1934.230 772.580 ;
        RECT 1932.990 669.360 1933.310 669.420 ;
        RECT 1932.795 669.220 1933.310 669.360 ;
        RECT 1932.990 669.160 1933.310 669.220 ;
        RECT 1933.005 614.620 1933.295 614.665 ;
        RECT 1933.450 614.620 1933.770 614.680 ;
        RECT 1933.005 614.480 1933.770 614.620 ;
        RECT 1933.005 614.435 1933.295 614.480 ;
        RECT 1933.450 614.420 1933.770 614.480 ;
        RECT 1932.990 607.140 1933.310 607.200 ;
        RECT 1934.385 607.140 1934.675 607.185 ;
        RECT 1932.990 607.000 1934.675 607.140 ;
        RECT 1932.990 606.940 1933.310 607.000 ;
        RECT 1934.385 606.955 1934.675 607.000 ;
        RECT 1934.370 517.720 1934.690 517.780 ;
        RECT 1934.370 517.580 1934.885 517.720 ;
        RECT 1934.370 517.520 1934.690 517.580 ;
        RECT 1933.910 469.780 1934.230 469.840 ;
        RECT 1933.910 469.640 1934.600 469.780 ;
        RECT 1933.910 469.580 1934.230 469.640 ;
        RECT 1934.460 469.500 1934.600 469.640 ;
        RECT 1934.370 469.240 1934.690 469.500 ;
        RECT 1932.990 386.960 1933.310 387.220 ;
        RECT 1933.080 386.540 1933.220 386.960 ;
        RECT 1932.990 386.280 1933.310 386.540 ;
        RECT 1932.990 307.260 1933.310 307.320 ;
        RECT 1933.910 307.260 1934.230 307.320 ;
        RECT 1932.990 307.120 1934.230 307.260 ;
        RECT 1932.990 307.060 1933.310 307.120 ;
        RECT 1933.910 307.060 1934.230 307.120 ;
        RECT 1933.450 241.300 1933.770 241.360 ;
        RECT 1933.910 241.300 1934.230 241.360 ;
        RECT 1933.450 241.160 1934.230 241.300 ;
        RECT 1933.450 241.100 1933.770 241.160 ;
        RECT 1933.910 241.100 1934.230 241.160 ;
        RECT 1933.910 145.420 1934.230 145.480 ;
        RECT 1933.540 145.280 1934.230 145.420 ;
        RECT 1933.540 145.140 1933.680 145.280 ;
        RECT 1933.910 145.220 1934.230 145.280 ;
        RECT 1933.450 144.880 1933.770 145.140 ;
        RECT 1628.010 33.900 1628.330 33.960 ;
        RECT 1932.530 33.900 1932.850 33.960 ;
        RECT 1628.010 33.760 1932.850 33.900 ;
        RECT 1628.010 33.700 1628.330 33.760 ;
        RECT 1932.530 33.700 1932.850 33.760 ;
        RECT 1530.950 16.560 1531.270 16.620 ;
        RECT 1628.010 16.560 1628.330 16.620 ;
        RECT 1530.950 16.420 1628.330 16.560 ;
        RECT 1530.950 16.360 1531.270 16.420 ;
        RECT 1628.010 16.360 1628.330 16.420 ;
      LAYER via ;
        RECT 1933.480 1642.240 1933.740 1642.500 ;
        RECT 1934.400 1642.240 1934.660 1642.500 ;
        RECT 1933.480 1593.620 1933.740 1593.880 ;
        RECT 1933.480 1545.680 1933.740 1545.940 ;
        RECT 1933.020 1435.180 1933.280 1435.440 ;
        RECT 1933.480 1393.700 1933.740 1393.960 ;
        RECT 1933.020 1366.160 1933.280 1366.420 ;
        RECT 1933.020 1345.760 1933.280 1346.020 ;
        RECT 1933.020 1321.280 1933.280 1321.540 ;
        RECT 1932.560 1297.140 1932.820 1297.400 ;
        RECT 1932.560 1255.660 1932.820 1255.920 ;
        RECT 1934.400 1255.660 1934.660 1255.920 ;
        RECT 1933.020 1159.100 1933.280 1159.360 ;
        RECT 1934.400 1159.100 1934.660 1159.360 ;
        RECT 1933.020 1062.540 1933.280 1062.800 ;
        RECT 1934.400 1062.540 1934.660 1062.800 ;
        RECT 1933.020 1048.600 1933.280 1048.860 ;
        RECT 1933.940 1048.600 1934.200 1048.860 ;
        RECT 1933.020 1000.320 1933.280 1000.580 ;
        RECT 1934.400 1000.320 1934.660 1000.580 ;
        RECT 1933.020 993.180 1933.280 993.440 ;
        RECT 1933.020 931.300 1933.280 931.560 ;
        RECT 1933.480 883.700 1933.740 883.960 ;
        RECT 1933.480 883.020 1933.740 883.280 ;
        RECT 1933.480 820.800 1933.740 821.060 ;
        RECT 1933.940 820.800 1934.200 821.060 ;
        RECT 1933.020 772.520 1933.280 772.780 ;
        RECT 1933.940 772.520 1934.200 772.780 ;
        RECT 1933.020 669.160 1933.280 669.420 ;
        RECT 1933.480 614.420 1933.740 614.680 ;
        RECT 1933.020 606.940 1933.280 607.200 ;
        RECT 1934.400 517.520 1934.660 517.780 ;
        RECT 1933.940 469.580 1934.200 469.840 ;
        RECT 1934.400 469.240 1934.660 469.500 ;
        RECT 1933.020 386.960 1933.280 387.220 ;
        RECT 1933.020 386.280 1933.280 386.540 ;
        RECT 1933.020 307.060 1933.280 307.320 ;
        RECT 1933.940 307.060 1934.200 307.320 ;
        RECT 1933.480 241.100 1933.740 241.360 ;
        RECT 1933.940 241.100 1934.200 241.360 ;
        RECT 1933.940 145.220 1934.200 145.480 ;
        RECT 1933.480 144.880 1933.740 145.140 ;
        RECT 1628.040 33.700 1628.300 33.960 ;
        RECT 1932.560 33.700 1932.820 33.960 ;
        RECT 1530.980 16.360 1531.240 16.620 ;
        RECT 1628.040 16.360 1628.300 16.620 ;
      LAYER met2 ;
        RECT 1936.620 1700.410 1936.900 1704.000 ;
        RECT 1934.460 1700.270 1936.900 1700.410 ;
        RECT 1934.460 1642.530 1934.600 1700.270 ;
        RECT 1936.620 1700.000 1936.900 1700.270 ;
        RECT 1933.480 1642.210 1933.740 1642.530 ;
        RECT 1934.400 1642.210 1934.660 1642.530 ;
        RECT 1933.540 1593.910 1933.680 1642.210 ;
        RECT 1933.480 1593.590 1933.740 1593.910 ;
        RECT 1933.480 1545.650 1933.740 1545.970 ;
        RECT 1933.540 1463.090 1933.680 1545.650 ;
        RECT 1933.080 1462.950 1933.680 1463.090 ;
        RECT 1933.080 1435.470 1933.220 1462.950 ;
        RECT 1933.020 1435.150 1933.280 1435.470 ;
        RECT 1933.540 1393.990 1933.680 1394.145 ;
        RECT 1933.480 1393.730 1933.740 1393.990 ;
        RECT 1933.080 1393.670 1933.740 1393.730 ;
        RECT 1933.080 1393.590 1933.680 1393.670 ;
        RECT 1933.080 1366.450 1933.220 1393.590 ;
        RECT 1933.020 1366.130 1933.280 1366.450 ;
        RECT 1933.020 1345.730 1933.280 1346.050 ;
        RECT 1933.080 1321.570 1933.220 1345.730 ;
        RECT 1933.020 1321.250 1933.280 1321.570 ;
        RECT 1932.560 1297.110 1932.820 1297.430 ;
        RECT 1932.620 1255.950 1932.760 1297.110 ;
        RECT 1932.560 1255.630 1932.820 1255.950 ;
        RECT 1934.400 1255.630 1934.660 1255.950 ;
        RECT 1934.460 1159.390 1934.600 1255.630 ;
        RECT 1933.020 1159.245 1933.280 1159.390 ;
        RECT 1934.400 1159.245 1934.660 1159.390 ;
        RECT 1933.010 1158.875 1933.290 1159.245 ;
        RECT 1934.390 1158.875 1934.670 1159.245 ;
        RECT 1934.460 1062.830 1934.600 1158.875 ;
        RECT 1933.020 1062.510 1933.280 1062.830 ;
        RECT 1934.400 1062.510 1934.660 1062.830 ;
        RECT 1933.080 1048.890 1933.220 1062.510 ;
        RECT 1933.020 1048.570 1933.280 1048.890 ;
        RECT 1933.940 1048.570 1934.200 1048.890 ;
        RECT 1934.000 1000.690 1934.140 1048.570 ;
        RECT 1934.000 1000.610 1934.600 1000.690 ;
        RECT 1933.020 1000.290 1933.280 1000.610 ;
        RECT 1934.000 1000.550 1934.660 1000.610 ;
        RECT 1934.400 1000.290 1934.660 1000.550 ;
        RECT 1933.080 993.470 1933.220 1000.290 ;
        RECT 1933.020 993.150 1933.280 993.470 ;
        RECT 1933.020 931.270 1933.280 931.590 ;
        RECT 1933.080 904.130 1933.220 931.270 ;
        RECT 1933.080 903.990 1933.680 904.130 ;
        RECT 1933.540 883.990 1933.680 903.990 ;
        RECT 1933.480 883.670 1933.740 883.990 ;
        RECT 1933.480 882.990 1933.740 883.310 ;
        RECT 1933.540 821.090 1933.680 882.990 ;
        RECT 1933.480 820.770 1933.740 821.090 ;
        RECT 1933.940 820.770 1934.200 821.090 ;
        RECT 1934.000 773.005 1934.140 820.770 ;
        RECT 1933.010 772.635 1933.290 773.005 ;
        RECT 1933.930 772.635 1934.210 773.005 ;
        RECT 1933.020 772.490 1933.280 772.635 ;
        RECT 1933.940 772.490 1934.200 772.635 ;
        RECT 1934.000 677.125 1934.140 772.490 ;
        RECT 1933.930 676.755 1934.210 677.125 ;
        RECT 1933.010 676.075 1933.290 676.445 ;
        RECT 1933.080 669.450 1933.220 676.075 ;
        RECT 1933.020 669.130 1933.280 669.450 ;
        RECT 1933.480 614.450 1933.740 614.710 ;
        RECT 1933.080 614.390 1933.740 614.450 ;
        RECT 1933.080 614.310 1933.680 614.390 ;
        RECT 1933.080 607.230 1933.220 614.310 ;
        RECT 1933.020 606.910 1933.280 607.230 ;
        RECT 1934.400 517.490 1934.660 517.810 ;
        RECT 1934.460 517.210 1934.600 517.490 ;
        RECT 1934.000 517.070 1934.600 517.210 ;
        RECT 1934.000 469.870 1934.140 517.070 ;
        RECT 1933.940 469.550 1934.200 469.870 ;
        RECT 1934.400 469.210 1934.660 469.530 ;
        RECT 1934.460 434.250 1934.600 469.210 ;
        RECT 1933.080 434.110 1934.600 434.250 ;
        RECT 1933.080 387.250 1933.220 434.110 ;
        RECT 1933.020 386.930 1933.280 387.250 ;
        RECT 1933.020 386.250 1933.280 386.570 ;
        RECT 1933.080 307.350 1933.220 386.250 ;
        RECT 1933.020 307.030 1933.280 307.350 ;
        RECT 1933.940 307.030 1934.200 307.350 ;
        RECT 1934.000 241.810 1934.140 307.030 ;
        RECT 1933.540 241.670 1934.140 241.810 ;
        RECT 1933.540 241.390 1933.680 241.670 ;
        RECT 1933.480 241.070 1933.740 241.390 ;
        RECT 1933.940 241.070 1934.200 241.390 ;
        RECT 1934.000 145.510 1934.140 241.070 ;
        RECT 1933.940 145.190 1934.200 145.510 ;
        RECT 1933.480 144.850 1933.740 145.170 ;
        RECT 1933.540 110.570 1933.680 144.850 ;
        RECT 1933.540 110.430 1934.140 110.570 ;
        RECT 1934.000 109.890 1934.140 110.430 ;
        RECT 1933.080 109.750 1934.140 109.890 ;
        RECT 1933.080 73.170 1933.220 109.750 ;
        RECT 1933.080 73.030 1933.680 73.170 ;
        RECT 1933.540 71.810 1933.680 73.030 ;
        RECT 1932.620 71.670 1933.680 71.810 ;
        RECT 1932.620 33.990 1932.760 71.670 ;
        RECT 1628.040 33.670 1628.300 33.990 ;
        RECT 1932.560 33.670 1932.820 33.990 ;
        RECT 1628.100 16.650 1628.240 33.670 ;
        RECT 1530.980 16.330 1531.240 16.650 ;
        RECT 1628.040 16.330 1628.300 16.650 ;
        RECT 1531.040 2.400 1531.180 16.330 ;
        RECT 1530.830 -4.800 1531.390 2.400 ;
      LAYER via2 ;
        RECT 1933.010 1158.920 1933.290 1159.200 ;
        RECT 1934.390 1158.920 1934.670 1159.200 ;
        RECT 1933.010 772.680 1933.290 772.960 ;
        RECT 1933.930 772.680 1934.210 772.960 ;
        RECT 1933.930 676.800 1934.210 677.080 ;
        RECT 1933.010 676.120 1933.290 676.400 ;
      LAYER met3 ;
        RECT 1932.985 1159.210 1933.315 1159.225 ;
        RECT 1934.365 1159.210 1934.695 1159.225 ;
        RECT 1932.985 1158.910 1934.695 1159.210 ;
        RECT 1932.985 1158.895 1933.315 1158.910 ;
        RECT 1934.365 1158.895 1934.695 1158.910 ;
        RECT 1932.985 772.970 1933.315 772.985 ;
        RECT 1933.905 772.970 1934.235 772.985 ;
        RECT 1932.985 772.670 1934.235 772.970 ;
        RECT 1932.985 772.655 1933.315 772.670 ;
        RECT 1933.905 772.655 1934.235 772.670 ;
        RECT 1933.905 677.090 1934.235 677.105 ;
        RECT 1932.310 676.790 1934.235 677.090 ;
        RECT 1932.310 676.410 1932.610 676.790 ;
        RECT 1933.905 676.775 1934.235 676.790 ;
        RECT 1932.985 676.410 1933.315 676.425 ;
        RECT 1932.310 676.110 1933.315 676.410 ;
        RECT 1932.985 676.095 1933.315 676.110 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1617.890 45.120 1618.210 45.180 ;
        RECT 1946.330 45.120 1946.650 45.180 ;
        RECT 1617.890 44.980 1946.650 45.120 ;
        RECT 1617.890 44.920 1618.210 44.980 ;
        RECT 1946.330 44.920 1946.650 44.980 ;
        RECT 1548.890 15.880 1549.210 15.940 ;
        RECT 1617.890 15.880 1618.210 15.940 ;
        RECT 1548.890 15.740 1618.210 15.880 ;
        RECT 1548.890 15.680 1549.210 15.740 ;
        RECT 1617.890 15.680 1618.210 15.740 ;
      LAYER via ;
        RECT 1617.920 44.920 1618.180 45.180 ;
        RECT 1946.360 44.920 1946.620 45.180 ;
        RECT 1548.920 15.680 1549.180 15.940 ;
        RECT 1617.920 15.680 1618.180 15.940 ;
      LAYER met2 ;
        RECT 1945.820 1700.410 1946.100 1704.000 ;
        RECT 1945.820 1700.270 1946.560 1700.410 ;
        RECT 1945.820 1700.000 1946.100 1700.270 ;
        RECT 1946.420 45.210 1946.560 1700.270 ;
        RECT 1617.920 44.890 1618.180 45.210 ;
        RECT 1946.360 44.890 1946.620 45.210 ;
        RECT 1617.980 15.970 1618.120 44.890 ;
        RECT 1548.920 15.650 1549.180 15.970 ;
        RECT 1617.920 15.650 1618.180 15.970 ;
        RECT 1548.980 2.400 1549.120 15.650 ;
        RECT 1548.770 -4.800 1549.330 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1627.550 45.800 1627.870 45.860 ;
        RECT 1953.230 45.800 1953.550 45.860 ;
        RECT 1627.550 45.660 1953.550 45.800 ;
        RECT 1627.550 45.600 1627.870 45.660 ;
        RECT 1953.230 45.600 1953.550 45.660 ;
        RECT 1566.830 15.540 1567.150 15.600 ;
        RECT 1627.550 15.540 1627.870 15.600 ;
        RECT 1566.830 15.400 1627.870 15.540 ;
        RECT 1566.830 15.340 1567.150 15.400 ;
        RECT 1627.550 15.340 1627.870 15.400 ;
      LAYER via ;
        RECT 1627.580 45.600 1627.840 45.860 ;
        RECT 1953.260 45.600 1953.520 45.860 ;
        RECT 1566.860 15.340 1567.120 15.600 ;
        RECT 1627.580 15.340 1627.840 15.600 ;
      LAYER met2 ;
        RECT 1955.020 1700.410 1955.300 1704.000 ;
        RECT 1953.320 1700.270 1955.300 1700.410 ;
        RECT 1953.320 45.890 1953.460 1700.270 ;
        RECT 1955.020 1700.000 1955.300 1700.270 ;
        RECT 1627.580 45.570 1627.840 45.890 ;
        RECT 1953.260 45.570 1953.520 45.890 ;
        RECT 1627.640 15.630 1627.780 45.570 ;
        RECT 1566.860 15.310 1567.120 15.630 ;
        RECT 1627.580 15.310 1627.840 15.630 ;
        RECT 1566.920 2.400 1567.060 15.310 ;
        RECT 1566.710 -4.800 1567.270 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1961.585 1594.005 1961.755 1642.115 ;
        RECT 1960.205 1297.185 1960.375 1321.495 ;
        RECT 1960.665 737.885 1960.835 772.735 ;
        RECT 1960.665 179.605 1960.835 241.315 ;
        RECT 1961.125 83.045 1961.295 131.155 ;
      LAYER mcon ;
        RECT 1961.585 1641.945 1961.755 1642.115 ;
        RECT 1960.205 1321.325 1960.375 1321.495 ;
        RECT 1960.665 772.565 1960.835 772.735 ;
        RECT 1960.665 241.145 1960.835 241.315 ;
        RECT 1961.125 130.985 1961.295 131.155 ;
      LAYER met1 ;
        RECT 1961.510 1642.100 1961.830 1642.160 ;
        RECT 1961.315 1641.960 1961.830 1642.100 ;
        RECT 1961.510 1641.900 1961.830 1641.960 ;
        RECT 1961.525 1594.160 1961.815 1594.205 ;
        RECT 1961.970 1594.160 1962.290 1594.220 ;
        RECT 1961.525 1594.020 1962.290 1594.160 ;
        RECT 1961.525 1593.975 1961.815 1594.020 ;
        RECT 1961.970 1593.960 1962.290 1594.020 ;
        RECT 1960.130 1554.720 1960.450 1554.780 ;
        RECT 1962.430 1554.720 1962.750 1554.780 ;
        RECT 1960.130 1554.580 1962.750 1554.720 ;
        RECT 1960.130 1554.520 1960.450 1554.580 ;
        RECT 1962.430 1554.520 1962.750 1554.580 ;
        RECT 1961.050 1462.920 1961.370 1462.980 ;
        RECT 1960.680 1462.780 1961.370 1462.920 ;
        RECT 1960.680 1462.640 1960.820 1462.780 ;
        RECT 1961.050 1462.720 1961.370 1462.780 ;
        RECT 1960.590 1462.380 1960.910 1462.640 ;
        RECT 1960.145 1321.480 1960.435 1321.525 ;
        RECT 1961.050 1321.480 1961.370 1321.540 ;
        RECT 1960.145 1321.340 1961.370 1321.480 ;
        RECT 1960.145 1321.295 1960.435 1321.340 ;
        RECT 1961.050 1321.280 1961.370 1321.340 ;
        RECT 1960.130 1297.340 1960.450 1297.400 ;
        RECT 1959.935 1297.200 1960.450 1297.340 ;
        RECT 1960.130 1297.140 1960.450 1297.200 ;
        RECT 1960.130 1207.580 1960.450 1207.640 ;
        RECT 1960.590 1207.580 1960.910 1207.640 ;
        RECT 1960.130 1207.440 1960.910 1207.580 ;
        RECT 1960.130 1207.380 1960.450 1207.440 ;
        RECT 1960.590 1207.380 1960.910 1207.440 ;
        RECT 1960.590 1111.020 1960.910 1111.080 ;
        RECT 1961.510 1111.020 1961.830 1111.080 ;
        RECT 1960.590 1110.880 1961.830 1111.020 ;
        RECT 1960.590 1110.820 1960.910 1110.880 ;
        RECT 1961.510 1110.820 1961.830 1110.880 ;
        RECT 1960.590 966.180 1960.910 966.240 ;
        RECT 1961.050 966.180 1961.370 966.240 ;
        RECT 1960.590 966.040 1961.370 966.180 ;
        RECT 1960.590 965.980 1960.910 966.040 ;
        RECT 1961.050 965.980 1961.370 966.040 ;
        RECT 1960.590 772.720 1960.910 772.780 ;
        RECT 1960.395 772.580 1960.910 772.720 ;
        RECT 1960.590 772.520 1960.910 772.580 ;
        RECT 1960.590 738.040 1960.910 738.100 ;
        RECT 1960.395 737.900 1960.910 738.040 ;
        RECT 1960.590 737.840 1960.910 737.900 ;
        RECT 1960.130 531.320 1960.450 531.380 ;
        RECT 1961.510 531.320 1961.830 531.380 ;
        RECT 1960.130 531.180 1961.830 531.320 ;
        RECT 1960.130 531.120 1960.450 531.180 ;
        RECT 1961.510 531.120 1961.830 531.180 ;
        RECT 1961.050 386.820 1961.370 386.880 ;
        RECT 1960.680 386.680 1961.370 386.820 ;
        RECT 1960.680 386.540 1960.820 386.680 ;
        RECT 1961.050 386.620 1961.370 386.680 ;
        RECT 1960.590 386.280 1960.910 386.540 ;
        RECT 1961.050 255.580 1961.370 255.640 ;
        RECT 1960.680 255.440 1961.370 255.580 ;
        RECT 1960.680 255.300 1960.820 255.440 ;
        RECT 1961.050 255.380 1961.370 255.440 ;
        RECT 1960.590 255.040 1960.910 255.300 ;
        RECT 1960.590 241.300 1960.910 241.360 ;
        RECT 1960.395 241.160 1960.910 241.300 ;
        RECT 1960.590 241.100 1960.910 241.160 ;
        RECT 1960.605 179.760 1960.895 179.805 ;
        RECT 1961.050 179.760 1961.370 179.820 ;
        RECT 1960.605 179.620 1961.370 179.760 ;
        RECT 1960.605 179.575 1960.895 179.620 ;
        RECT 1961.050 179.560 1961.370 179.620 ;
        RECT 1961.050 131.140 1961.370 131.200 ;
        RECT 1960.855 131.000 1961.370 131.140 ;
        RECT 1961.050 130.940 1961.370 131.000 ;
        RECT 1961.050 83.200 1961.370 83.260 ;
        RECT 1960.855 83.060 1961.370 83.200 ;
        RECT 1961.050 83.000 1961.370 83.060 ;
        RECT 1960.130 73.340 1960.450 73.400 ;
        RECT 1961.050 73.340 1961.370 73.400 ;
        RECT 1960.130 73.200 1961.370 73.340 ;
        RECT 1960.130 73.140 1960.450 73.200 ;
        RECT 1961.050 73.140 1961.370 73.200 ;
        RECT 1635.370 46.140 1635.690 46.200 ;
        RECT 1960.130 46.140 1960.450 46.200 ;
        RECT 1635.370 46.000 1960.450 46.140 ;
        RECT 1635.370 45.940 1635.690 46.000 ;
        RECT 1960.130 45.940 1960.450 46.000 ;
        RECT 1584.770 19.280 1585.090 19.340 ;
        RECT 1635.370 19.280 1635.690 19.340 ;
        RECT 1584.770 19.140 1635.690 19.280 ;
        RECT 1584.770 19.080 1585.090 19.140 ;
        RECT 1635.370 19.080 1635.690 19.140 ;
      LAYER via ;
        RECT 1961.540 1641.900 1961.800 1642.160 ;
        RECT 1962.000 1593.960 1962.260 1594.220 ;
        RECT 1960.160 1554.520 1960.420 1554.780 ;
        RECT 1962.460 1554.520 1962.720 1554.780 ;
        RECT 1961.080 1462.720 1961.340 1462.980 ;
        RECT 1960.620 1462.380 1960.880 1462.640 ;
        RECT 1961.080 1321.280 1961.340 1321.540 ;
        RECT 1960.160 1297.140 1960.420 1297.400 ;
        RECT 1960.160 1207.380 1960.420 1207.640 ;
        RECT 1960.620 1207.380 1960.880 1207.640 ;
        RECT 1960.620 1110.820 1960.880 1111.080 ;
        RECT 1961.540 1110.820 1961.800 1111.080 ;
        RECT 1960.620 965.980 1960.880 966.240 ;
        RECT 1961.080 965.980 1961.340 966.240 ;
        RECT 1960.620 772.520 1960.880 772.780 ;
        RECT 1960.620 737.840 1960.880 738.100 ;
        RECT 1960.160 531.120 1960.420 531.380 ;
        RECT 1961.540 531.120 1961.800 531.380 ;
        RECT 1961.080 386.620 1961.340 386.880 ;
        RECT 1960.620 386.280 1960.880 386.540 ;
        RECT 1961.080 255.380 1961.340 255.640 ;
        RECT 1960.620 255.040 1960.880 255.300 ;
        RECT 1960.620 241.100 1960.880 241.360 ;
        RECT 1961.080 179.560 1961.340 179.820 ;
        RECT 1961.080 130.940 1961.340 131.200 ;
        RECT 1961.080 83.000 1961.340 83.260 ;
        RECT 1960.160 73.140 1960.420 73.400 ;
        RECT 1961.080 73.140 1961.340 73.400 ;
        RECT 1635.400 45.940 1635.660 46.200 ;
        RECT 1960.160 45.940 1960.420 46.200 ;
        RECT 1584.800 19.080 1585.060 19.340 ;
        RECT 1635.400 19.080 1635.660 19.340 ;
      LAYER met2 ;
        RECT 1964.220 1701.090 1964.500 1704.000 ;
        RECT 1961.600 1700.950 1964.500 1701.090 ;
        RECT 1961.600 1690.210 1961.740 1700.950 ;
        RECT 1964.220 1700.000 1964.500 1700.950 ;
        RECT 1961.600 1690.070 1962.200 1690.210 ;
        RECT 1962.060 1642.610 1962.200 1690.070 ;
        RECT 1961.600 1642.470 1962.200 1642.610 ;
        RECT 1961.600 1642.190 1961.740 1642.470 ;
        RECT 1961.540 1641.870 1961.800 1642.190 ;
        RECT 1962.000 1593.930 1962.260 1594.250 ;
        RECT 1962.060 1593.650 1962.200 1593.930 ;
        RECT 1962.060 1593.510 1962.660 1593.650 ;
        RECT 1962.520 1554.810 1962.660 1593.510 ;
        RECT 1960.160 1554.490 1960.420 1554.810 ;
        RECT 1962.460 1554.490 1962.720 1554.810 ;
        RECT 1960.220 1490.970 1960.360 1554.490 ;
        RECT 1960.220 1490.830 1960.820 1490.970 ;
        RECT 1960.680 1483.490 1960.820 1490.830 ;
        RECT 1960.680 1483.350 1961.280 1483.490 ;
        RECT 1961.140 1463.010 1961.280 1483.350 ;
        RECT 1961.080 1462.690 1961.340 1463.010 ;
        RECT 1960.620 1462.350 1960.880 1462.670 ;
        RECT 1960.680 1393.845 1960.820 1462.350 ;
        RECT 1960.610 1393.475 1960.890 1393.845 ;
        RECT 1961.070 1392.795 1961.350 1393.165 ;
        RECT 1961.140 1321.570 1961.280 1392.795 ;
        RECT 1961.080 1321.250 1961.340 1321.570 ;
        RECT 1960.160 1297.110 1960.420 1297.430 ;
        RECT 1960.220 1207.670 1960.360 1297.110 ;
        RECT 1960.160 1207.350 1960.420 1207.670 ;
        RECT 1960.620 1207.525 1960.880 1207.670 ;
        RECT 1960.610 1207.155 1960.890 1207.525 ;
        RECT 1961.530 1207.155 1961.810 1207.525 ;
        RECT 1961.600 1200.725 1961.740 1207.155 ;
        RECT 1961.530 1200.355 1961.810 1200.725 ;
        RECT 1962.450 1200.355 1962.730 1200.725 ;
        RECT 1962.520 1157.770 1962.660 1200.355 ;
        RECT 1961.600 1157.630 1962.660 1157.770 ;
        RECT 1961.600 1111.110 1961.740 1157.630 ;
        RECT 1960.620 1110.965 1960.880 1111.110 ;
        RECT 1960.610 1110.595 1960.890 1110.965 ;
        RECT 1961.540 1110.790 1961.800 1111.110 ;
        RECT 1961.070 1109.915 1961.350 1110.285 ;
        RECT 1961.140 1014.290 1961.280 1109.915 ;
        RECT 1960.680 1014.150 1961.280 1014.290 ;
        RECT 1960.680 966.270 1960.820 1014.150 ;
        RECT 1960.620 965.950 1960.880 966.270 ;
        RECT 1961.080 965.950 1961.340 966.270 ;
        RECT 1961.140 883.730 1961.280 965.950 ;
        RECT 1960.680 883.590 1961.280 883.730 ;
        RECT 1960.680 773.685 1960.820 883.590 ;
        RECT 1960.610 773.315 1960.890 773.685 ;
        RECT 1960.610 772.635 1960.890 773.005 ;
        RECT 1960.620 772.490 1960.880 772.635 ;
        RECT 1960.620 737.810 1960.880 738.130 ;
        RECT 1960.680 724.610 1960.820 737.810 ;
        RECT 1960.680 724.470 1961.280 724.610 ;
        RECT 1961.140 691.405 1961.280 724.470 ;
        RECT 1961.070 691.035 1961.350 691.405 ;
        RECT 1960.610 676.075 1960.890 676.445 ;
        RECT 1960.680 628.050 1960.820 676.075 ;
        RECT 1960.680 627.910 1961.280 628.050 ;
        RECT 1961.140 596.770 1961.280 627.910 ;
        RECT 1960.680 596.630 1961.280 596.770 ;
        RECT 1960.680 593.370 1960.820 596.630 ;
        RECT 1960.680 593.230 1961.280 593.370 ;
        RECT 1961.140 592.010 1961.280 593.230 ;
        RECT 1960.680 591.870 1961.280 592.010 ;
        RECT 1960.680 545.090 1960.820 591.870 ;
        RECT 1960.680 544.950 1961.740 545.090 ;
        RECT 1961.600 531.410 1961.740 544.950 ;
        RECT 1960.160 531.090 1960.420 531.410 ;
        RECT 1961.540 531.090 1961.800 531.410 ;
        RECT 1960.220 483.325 1960.360 531.090 ;
        RECT 1960.150 482.955 1960.430 483.325 ;
        RECT 1961.070 482.955 1961.350 483.325 ;
        RECT 1961.140 386.910 1961.280 482.955 ;
        RECT 1961.080 386.590 1961.340 386.910 ;
        RECT 1960.620 386.250 1960.880 386.570 ;
        RECT 1960.680 351.290 1960.820 386.250 ;
        RECT 1960.680 351.150 1961.280 351.290 ;
        RECT 1961.140 255.670 1961.280 351.150 ;
        RECT 1961.080 255.350 1961.340 255.670 ;
        RECT 1960.620 255.010 1960.880 255.330 ;
        RECT 1960.680 241.390 1960.820 255.010 ;
        RECT 1960.620 241.070 1960.880 241.390 ;
        RECT 1961.080 179.530 1961.340 179.850 ;
        RECT 1961.140 131.230 1961.280 179.530 ;
        RECT 1961.080 130.910 1961.340 131.230 ;
        RECT 1961.080 82.970 1961.340 83.290 ;
        RECT 1961.140 73.430 1961.280 82.970 ;
        RECT 1960.160 73.110 1960.420 73.430 ;
        RECT 1961.080 73.110 1961.340 73.430 ;
        RECT 1960.220 46.230 1960.360 73.110 ;
        RECT 1635.400 45.910 1635.660 46.230 ;
        RECT 1960.160 45.910 1960.420 46.230 ;
        RECT 1635.460 19.370 1635.600 45.910 ;
        RECT 1584.800 19.050 1585.060 19.370 ;
        RECT 1635.400 19.050 1635.660 19.370 ;
        RECT 1584.860 2.400 1585.000 19.050 ;
        RECT 1584.650 -4.800 1585.210 2.400 ;
      LAYER via2 ;
        RECT 1960.610 1393.520 1960.890 1393.800 ;
        RECT 1961.070 1392.840 1961.350 1393.120 ;
        RECT 1960.610 1207.200 1960.890 1207.480 ;
        RECT 1961.530 1207.200 1961.810 1207.480 ;
        RECT 1961.530 1200.400 1961.810 1200.680 ;
        RECT 1962.450 1200.400 1962.730 1200.680 ;
        RECT 1960.610 1110.640 1960.890 1110.920 ;
        RECT 1961.070 1109.960 1961.350 1110.240 ;
        RECT 1960.610 773.360 1960.890 773.640 ;
        RECT 1960.610 772.680 1960.890 772.960 ;
        RECT 1961.070 691.080 1961.350 691.360 ;
        RECT 1960.610 676.120 1960.890 676.400 ;
        RECT 1960.150 483.000 1960.430 483.280 ;
        RECT 1961.070 483.000 1961.350 483.280 ;
      LAYER met3 ;
        RECT 1960.585 1393.810 1960.915 1393.825 ;
        RECT 1959.910 1393.510 1960.915 1393.810 ;
        RECT 1959.910 1393.130 1960.210 1393.510 ;
        RECT 1960.585 1393.495 1960.915 1393.510 ;
        RECT 1961.045 1393.130 1961.375 1393.145 ;
        RECT 1959.910 1392.830 1961.375 1393.130 ;
        RECT 1961.045 1392.815 1961.375 1392.830 ;
        RECT 1960.585 1207.490 1960.915 1207.505 ;
        RECT 1961.505 1207.490 1961.835 1207.505 ;
        RECT 1960.585 1207.190 1961.835 1207.490 ;
        RECT 1960.585 1207.175 1960.915 1207.190 ;
        RECT 1961.505 1207.175 1961.835 1207.190 ;
        RECT 1961.505 1200.690 1961.835 1200.705 ;
        RECT 1962.425 1200.690 1962.755 1200.705 ;
        RECT 1961.505 1200.390 1962.755 1200.690 ;
        RECT 1961.505 1200.375 1961.835 1200.390 ;
        RECT 1962.425 1200.375 1962.755 1200.390 ;
        RECT 1960.585 1110.930 1960.915 1110.945 ;
        RECT 1960.585 1110.615 1961.130 1110.930 ;
        RECT 1960.830 1110.265 1961.130 1110.615 ;
        RECT 1960.830 1109.950 1961.375 1110.265 ;
        RECT 1961.045 1109.935 1961.375 1109.950 ;
        RECT 1960.585 773.650 1960.915 773.665 ;
        RECT 1960.585 773.335 1961.130 773.650 ;
        RECT 1960.830 772.985 1961.130 773.335 ;
        RECT 1960.585 772.670 1961.130 772.985 ;
        RECT 1960.585 772.655 1960.915 772.670 ;
        RECT 1961.045 691.380 1961.375 691.385 ;
        RECT 1960.790 691.370 1961.375 691.380 ;
        RECT 1960.590 691.070 1961.375 691.370 ;
        RECT 1960.790 691.060 1961.375 691.070 ;
        RECT 1961.045 691.055 1961.375 691.060 ;
        RECT 1960.585 676.420 1960.915 676.425 ;
        RECT 1960.585 676.410 1961.170 676.420 ;
        RECT 1960.360 676.110 1961.170 676.410 ;
        RECT 1960.585 676.100 1961.170 676.110 ;
        RECT 1960.585 676.095 1960.915 676.100 ;
        RECT 1960.125 483.290 1960.455 483.305 ;
        RECT 1961.045 483.290 1961.375 483.305 ;
        RECT 1960.125 482.990 1961.375 483.290 ;
        RECT 1960.125 482.975 1960.455 482.990 ;
        RECT 1961.045 482.975 1961.375 482.990 ;
      LAYER via3 ;
        RECT 1960.820 691.060 1961.140 691.380 ;
        RECT 1960.820 676.100 1961.140 676.420 ;
      LAYER met4 ;
        RECT 1960.815 691.055 1961.145 691.385 ;
        RECT 1960.830 676.425 1961.130 691.055 ;
        RECT 1960.815 676.095 1961.145 676.425 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1642.730 45.460 1643.050 45.520 ;
        RECT 1973.930 45.460 1974.250 45.520 ;
        RECT 1642.730 45.320 1974.250 45.460 ;
        RECT 1642.730 45.260 1643.050 45.320 ;
        RECT 1973.930 45.260 1974.250 45.320 ;
        RECT 1602.250 15.200 1602.570 15.260 ;
        RECT 1642.730 15.200 1643.050 15.260 ;
        RECT 1602.250 15.060 1643.050 15.200 ;
        RECT 1602.250 15.000 1602.570 15.060 ;
        RECT 1642.730 15.000 1643.050 15.060 ;
      LAYER via ;
        RECT 1642.760 45.260 1643.020 45.520 ;
        RECT 1973.960 45.260 1974.220 45.520 ;
        RECT 1602.280 15.000 1602.540 15.260 ;
        RECT 1642.760 15.000 1643.020 15.260 ;
      LAYER met2 ;
        RECT 1973.420 1700.410 1973.700 1704.000 ;
        RECT 1973.420 1700.270 1974.160 1700.410 ;
        RECT 1973.420 1700.000 1973.700 1700.270 ;
        RECT 1974.020 45.550 1974.160 1700.270 ;
        RECT 1642.760 45.230 1643.020 45.550 ;
        RECT 1973.960 45.230 1974.220 45.550 ;
        RECT 1642.820 15.290 1642.960 45.230 ;
        RECT 1602.280 14.970 1602.540 15.290 ;
        RECT 1642.760 14.970 1643.020 15.290 ;
        RECT 1602.340 2.400 1602.480 14.970 ;
        RECT 1602.130 -4.800 1602.690 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1732.430 36.280 1732.750 36.340 ;
        RECT 1980.830 36.280 1981.150 36.340 ;
        RECT 1732.430 36.140 1981.150 36.280 ;
        RECT 1732.430 36.080 1732.750 36.140 ;
        RECT 1980.830 36.080 1981.150 36.140 ;
        RECT 1620.190 16.900 1620.510 16.960 ;
        RECT 1732.430 16.900 1732.750 16.960 ;
        RECT 1620.190 16.760 1732.750 16.900 ;
        RECT 1620.190 16.700 1620.510 16.760 ;
        RECT 1732.430 16.700 1732.750 16.760 ;
      LAYER via ;
        RECT 1732.460 36.080 1732.720 36.340 ;
        RECT 1980.860 36.080 1981.120 36.340 ;
        RECT 1620.220 16.700 1620.480 16.960 ;
        RECT 1732.460 16.700 1732.720 16.960 ;
      LAYER met2 ;
        RECT 1982.620 1700.410 1982.900 1704.000 ;
        RECT 1980.920 1700.270 1982.900 1700.410 ;
        RECT 1980.920 36.370 1981.060 1700.270 ;
        RECT 1982.620 1700.000 1982.900 1700.270 ;
        RECT 1732.460 36.050 1732.720 36.370 ;
        RECT 1980.860 36.050 1981.120 36.370 ;
        RECT 1732.520 16.990 1732.660 36.050 ;
        RECT 1620.220 16.670 1620.480 16.990 ;
        RECT 1732.460 16.670 1732.720 16.990 ;
        RECT 1620.280 2.400 1620.420 16.670 ;
        RECT 1620.070 -4.800 1620.630 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1989.185 1594.005 1989.355 1642.115 ;
        RECT 1988.725 1442.025 1988.895 1490.475 ;
        RECT 1988.265 1345.465 1988.435 1392.895 ;
        RECT 1987.805 1248.905 1987.975 1269.815 ;
        RECT 1987.805 1200.625 1987.975 1224.935 ;
        RECT 1988.725 869.465 1988.895 883.235 ;
        RECT 1988.725 772.905 1988.895 821.015 ;
        RECT 1988.725 717.825 1988.895 724.795 ;
        RECT 1988.265 524.705 1988.435 572.475 ;
        RECT 1988.725 234.685 1988.895 282.795 ;
        RECT 1987.805 48.365 1987.975 96.475 ;
        RECT 1675.925 15.725 1676.095 16.575 ;
      LAYER mcon ;
        RECT 1989.185 1641.945 1989.355 1642.115 ;
        RECT 1988.725 1490.305 1988.895 1490.475 ;
        RECT 1988.265 1392.725 1988.435 1392.895 ;
        RECT 1987.805 1269.645 1987.975 1269.815 ;
        RECT 1987.805 1224.765 1987.975 1224.935 ;
        RECT 1988.725 883.065 1988.895 883.235 ;
        RECT 1988.725 820.845 1988.895 821.015 ;
        RECT 1988.725 724.625 1988.895 724.795 ;
        RECT 1988.265 572.305 1988.435 572.475 ;
        RECT 1988.725 282.625 1988.895 282.795 ;
        RECT 1987.805 96.305 1987.975 96.475 ;
        RECT 1675.925 16.405 1676.095 16.575 ;
      LAYER met1 ;
        RECT 1989.110 1642.100 1989.430 1642.160 ;
        RECT 1988.915 1641.960 1989.430 1642.100 ;
        RECT 1989.110 1641.900 1989.430 1641.960 ;
        RECT 1989.125 1594.160 1989.415 1594.205 ;
        RECT 1989.570 1594.160 1989.890 1594.220 ;
        RECT 1989.125 1594.020 1989.890 1594.160 ;
        RECT 1989.125 1593.975 1989.415 1594.020 ;
        RECT 1989.570 1593.960 1989.890 1594.020 ;
        RECT 1987.730 1559.480 1988.050 1559.540 ;
        RECT 1989.570 1559.480 1989.890 1559.540 ;
        RECT 1987.730 1559.340 1989.890 1559.480 ;
        RECT 1987.730 1559.280 1988.050 1559.340 ;
        RECT 1989.570 1559.280 1989.890 1559.340 ;
        RECT 1988.650 1490.460 1988.970 1490.520 ;
        RECT 1988.455 1490.320 1988.970 1490.460 ;
        RECT 1988.650 1490.260 1988.970 1490.320 ;
        RECT 1988.650 1442.180 1988.970 1442.240 ;
        RECT 1988.455 1442.040 1988.970 1442.180 ;
        RECT 1988.650 1441.980 1988.970 1442.040 ;
        RECT 1988.190 1393.900 1988.510 1393.960 ;
        RECT 1988.650 1393.900 1988.970 1393.960 ;
        RECT 1988.190 1393.760 1988.970 1393.900 ;
        RECT 1988.190 1393.700 1988.510 1393.760 ;
        RECT 1988.650 1393.700 1988.970 1393.760 ;
        RECT 1988.190 1392.880 1988.510 1392.940 ;
        RECT 1987.995 1392.740 1988.510 1392.880 ;
        RECT 1988.190 1392.680 1988.510 1392.740 ;
        RECT 1988.205 1345.620 1988.495 1345.665 ;
        RECT 1989.570 1345.620 1989.890 1345.680 ;
        RECT 1988.205 1345.480 1989.890 1345.620 ;
        RECT 1988.205 1345.435 1988.495 1345.480 ;
        RECT 1989.570 1345.420 1989.890 1345.480 ;
        RECT 1988.190 1304.480 1988.510 1304.540 ;
        RECT 1989.570 1304.480 1989.890 1304.540 ;
        RECT 1988.190 1304.340 1989.890 1304.480 ;
        RECT 1988.190 1304.280 1988.510 1304.340 ;
        RECT 1989.570 1304.280 1989.890 1304.340 ;
        RECT 1987.745 1269.800 1988.035 1269.845 ;
        RECT 1988.650 1269.800 1988.970 1269.860 ;
        RECT 1987.745 1269.660 1988.970 1269.800 ;
        RECT 1987.745 1269.615 1988.035 1269.660 ;
        RECT 1988.650 1269.600 1988.970 1269.660 ;
        RECT 1987.730 1249.060 1988.050 1249.120 ;
        RECT 1987.535 1248.920 1988.050 1249.060 ;
        RECT 1987.730 1248.860 1988.050 1248.920 ;
        RECT 1987.730 1224.920 1988.050 1224.980 ;
        RECT 1987.535 1224.780 1988.050 1224.920 ;
        RECT 1987.730 1224.720 1988.050 1224.780 ;
        RECT 1987.745 1200.780 1988.035 1200.825 ;
        RECT 1988.190 1200.780 1988.510 1200.840 ;
        RECT 1987.745 1200.640 1988.510 1200.780 ;
        RECT 1987.745 1200.595 1988.035 1200.640 ;
        RECT 1988.190 1200.580 1988.510 1200.640 ;
        RECT 1988.190 1173.380 1988.510 1173.640 ;
        RECT 1988.280 1172.960 1988.420 1173.380 ;
        RECT 1988.190 1172.700 1988.510 1172.960 ;
        RECT 1988.650 966.180 1988.970 966.240 ;
        RECT 1989.570 966.180 1989.890 966.240 ;
        RECT 1988.650 966.040 1989.890 966.180 ;
        RECT 1988.650 965.980 1988.970 966.040 ;
        RECT 1989.570 965.980 1989.890 966.040 ;
        RECT 1988.650 883.220 1988.970 883.280 ;
        RECT 1988.455 883.080 1988.970 883.220 ;
        RECT 1988.650 883.020 1988.970 883.080 ;
        RECT 1988.650 869.620 1988.970 869.680 ;
        RECT 1988.455 869.480 1988.970 869.620 ;
        RECT 1988.650 869.420 1988.970 869.480 ;
        RECT 1988.650 821.000 1988.970 821.060 ;
        RECT 1988.455 820.860 1988.970 821.000 ;
        RECT 1988.650 820.800 1988.970 820.860 ;
        RECT 1988.650 773.060 1988.970 773.120 ;
        RECT 1988.455 772.920 1988.970 773.060 ;
        RECT 1988.650 772.860 1988.970 772.920 ;
        RECT 1988.650 724.780 1988.970 724.840 ;
        RECT 1988.455 724.640 1988.970 724.780 ;
        RECT 1988.650 724.580 1988.970 724.640 ;
        RECT 1988.650 717.980 1988.970 718.040 ;
        RECT 1988.650 717.840 1989.165 717.980 ;
        RECT 1988.650 717.780 1988.970 717.840 ;
        RECT 1988.650 621.080 1988.970 621.140 ;
        RECT 1989.570 621.080 1989.890 621.140 ;
        RECT 1988.650 620.940 1989.890 621.080 ;
        RECT 1988.650 620.880 1988.970 620.940 ;
        RECT 1989.570 620.880 1989.890 620.940 ;
        RECT 1988.205 572.460 1988.495 572.505 ;
        RECT 1988.650 572.460 1988.970 572.520 ;
        RECT 1988.205 572.320 1988.970 572.460 ;
        RECT 1988.205 572.275 1988.495 572.320 ;
        RECT 1988.650 572.260 1988.970 572.320 ;
        RECT 1988.190 524.860 1988.510 524.920 ;
        RECT 1987.995 524.720 1988.510 524.860 ;
        RECT 1988.190 524.660 1988.510 524.720 ;
        RECT 1988.190 523.980 1988.510 524.240 ;
        RECT 1988.280 523.840 1988.420 523.980 ;
        RECT 1989.110 523.840 1989.430 523.900 ;
        RECT 1988.280 523.700 1989.430 523.840 ;
        RECT 1989.110 523.640 1989.430 523.700 ;
        RECT 1988.665 282.780 1988.955 282.825 ;
        RECT 1989.110 282.780 1989.430 282.840 ;
        RECT 1988.665 282.640 1989.430 282.780 ;
        RECT 1988.665 282.595 1988.955 282.640 ;
        RECT 1989.110 282.580 1989.430 282.640 ;
        RECT 1988.650 234.840 1988.970 234.900 ;
        RECT 1988.455 234.700 1988.970 234.840 ;
        RECT 1988.650 234.640 1988.970 234.700 ;
        RECT 1987.745 96.460 1988.035 96.505 ;
        RECT 1988.190 96.460 1988.510 96.520 ;
        RECT 1987.745 96.320 1988.510 96.460 ;
        RECT 1987.745 96.275 1988.035 96.320 ;
        RECT 1988.190 96.260 1988.510 96.320 ;
        RECT 1987.730 48.520 1988.050 48.580 ;
        RECT 1987.535 48.380 1988.050 48.520 ;
        RECT 1987.730 48.320 1988.050 48.380 ;
        RECT 1739.790 36.620 1740.110 36.680 ;
        RECT 1987.730 36.620 1988.050 36.680 ;
        RECT 1739.790 36.480 1988.050 36.620 ;
        RECT 1739.790 36.420 1740.110 36.480 ;
        RECT 1987.730 36.420 1988.050 36.480 ;
        RECT 1675.865 16.560 1676.155 16.605 ;
        RECT 1739.790 16.560 1740.110 16.620 ;
        RECT 1675.865 16.420 1740.110 16.560 ;
        RECT 1675.865 16.375 1676.155 16.420 ;
        RECT 1739.790 16.360 1740.110 16.420 ;
        RECT 1638.130 15.880 1638.450 15.940 ;
        RECT 1675.865 15.880 1676.155 15.925 ;
        RECT 1638.130 15.740 1676.155 15.880 ;
        RECT 1638.130 15.680 1638.450 15.740 ;
        RECT 1675.865 15.695 1676.155 15.740 ;
      LAYER via ;
        RECT 1989.140 1641.900 1989.400 1642.160 ;
        RECT 1989.600 1593.960 1989.860 1594.220 ;
        RECT 1987.760 1559.280 1988.020 1559.540 ;
        RECT 1989.600 1559.280 1989.860 1559.540 ;
        RECT 1988.680 1490.260 1988.940 1490.520 ;
        RECT 1988.680 1441.980 1988.940 1442.240 ;
        RECT 1988.220 1393.700 1988.480 1393.960 ;
        RECT 1988.680 1393.700 1988.940 1393.960 ;
        RECT 1988.220 1392.680 1988.480 1392.940 ;
        RECT 1989.600 1345.420 1989.860 1345.680 ;
        RECT 1988.220 1304.280 1988.480 1304.540 ;
        RECT 1989.600 1304.280 1989.860 1304.540 ;
        RECT 1988.680 1269.600 1988.940 1269.860 ;
        RECT 1987.760 1248.860 1988.020 1249.120 ;
        RECT 1987.760 1224.720 1988.020 1224.980 ;
        RECT 1988.220 1200.580 1988.480 1200.840 ;
        RECT 1988.220 1173.380 1988.480 1173.640 ;
        RECT 1988.220 1172.700 1988.480 1172.960 ;
        RECT 1988.680 965.980 1988.940 966.240 ;
        RECT 1989.600 965.980 1989.860 966.240 ;
        RECT 1988.680 883.020 1988.940 883.280 ;
        RECT 1988.680 869.420 1988.940 869.680 ;
        RECT 1988.680 820.800 1988.940 821.060 ;
        RECT 1988.680 772.860 1988.940 773.120 ;
        RECT 1988.680 724.580 1988.940 724.840 ;
        RECT 1988.680 717.780 1988.940 718.040 ;
        RECT 1988.680 620.880 1988.940 621.140 ;
        RECT 1989.600 620.880 1989.860 621.140 ;
        RECT 1988.680 572.260 1988.940 572.520 ;
        RECT 1988.220 524.660 1988.480 524.920 ;
        RECT 1988.220 523.980 1988.480 524.240 ;
        RECT 1989.140 523.640 1989.400 523.900 ;
        RECT 1989.140 282.580 1989.400 282.840 ;
        RECT 1988.680 234.640 1988.940 234.900 ;
        RECT 1988.220 96.260 1988.480 96.520 ;
        RECT 1987.760 48.320 1988.020 48.580 ;
        RECT 1739.820 36.420 1740.080 36.680 ;
        RECT 1987.760 36.420 1988.020 36.680 ;
        RECT 1739.820 16.360 1740.080 16.620 ;
        RECT 1638.160 15.680 1638.420 15.940 ;
      LAYER met2 ;
        RECT 1991.820 1701.090 1992.100 1704.000 ;
        RECT 1989.200 1700.950 1992.100 1701.090 ;
        RECT 1989.200 1642.190 1989.340 1700.950 ;
        RECT 1991.820 1700.000 1992.100 1700.950 ;
        RECT 1989.140 1641.870 1989.400 1642.190 ;
        RECT 1989.600 1593.930 1989.860 1594.250 ;
        RECT 1989.660 1559.570 1989.800 1593.930 ;
        RECT 1987.760 1559.250 1988.020 1559.570 ;
        RECT 1989.600 1559.250 1989.860 1559.570 ;
        RECT 1987.820 1510.690 1987.960 1559.250 ;
        RECT 1987.820 1510.550 1988.420 1510.690 ;
        RECT 1988.280 1497.090 1988.420 1510.550 ;
        RECT 1988.280 1496.950 1988.880 1497.090 ;
        RECT 1988.740 1490.550 1988.880 1496.950 ;
        RECT 1988.680 1490.230 1988.940 1490.550 ;
        RECT 1988.680 1441.950 1988.940 1442.270 ;
        RECT 1988.740 1393.990 1988.880 1441.950 ;
        RECT 1988.220 1393.670 1988.480 1393.990 ;
        RECT 1988.680 1393.670 1988.940 1393.990 ;
        RECT 1988.280 1392.970 1988.420 1393.670 ;
        RECT 1988.220 1392.650 1988.480 1392.970 ;
        RECT 1989.600 1345.390 1989.860 1345.710 ;
        RECT 1989.660 1304.570 1989.800 1345.390 ;
        RECT 1988.220 1304.250 1988.480 1304.570 ;
        RECT 1989.600 1304.250 1989.860 1304.570 ;
        RECT 1988.280 1297.170 1988.420 1304.250 ;
        RECT 1988.280 1297.030 1988.880 1297.170 ;
        RECT 1988.740 1269.890 1988.880 1297.030 ;
        RECT 1988.680 1269.570 1988.940 1269.890 ;
        RECT 1987.760 1248.830 1988.020 1249.150 ;
        RECT 1987.820 1225.010 1987.960 1248.830 ;
        RECT 1987.760 1224.690 1988.020 1225.010 ;
        RECT 1988.220 1200.550 1988.480 1200.870 ;
        RECT 1988.280 1173.670 1988.420 1200.550 ;
        RECT 1988.220 1173.350 1988.480 1173.670 ;
        RECT 1988.220 1172.670 1988.480 1172.990 ;
        RECT 1988.280 1135.330 1988.420 1172.670 ;
        RECT 1987.820 1135.190 1988.420 1135.330 ;
        RECT 1987.820 1076.340 1987.960 1135.190 ;
        RECT 1987.820 1076.200 1988.880 1076.340 ;
        RECT 1988.740 1014.290 1988.880 1076.200 ;
        RECT 1988.740 1014.150 1989.800 1014.290 ;
        RECT 1989.660 966.270 1989.800 1014.150 ;
        RECT 1988.680 965.950 1988.940 966.270 ;
        RECT 1989.600 965.950 1989.860 966.270 ;
        RECT 1988.740 883.310 1988.880 965.950 ;
        RECT 1988.680 882.990 1988.940 883.310 ;
        RECT 1988.680 869.390 1988.940 869.710 ;
        RECT 1988.740 821.090 1988.880 869.390 ;
        RECT 1988.680 820.770 1988.940 821.090 ;
        RECT 1988.680 772.830 1988.940 773.150 ;
        RECT 1988.740 724.870 1988.880 772.830 ;
        RECT 1988.680 724.550 1988.940 724.870 ;
        RECT 1988.680 717.750 1988.940 718.070 ;
        RECT 1988.740 621.170 1988.880 717.750 ;
        RECT 1988.680 620.850 1988.940 621.170 ;
        RECT 1989.600 620.850 1989.860 621.170 ;
        RECT 1989.660 579.885 1989.800 620.850 ;
        RECT 1988.670 579.515 1988.950 579.885 ;
        RECT 1989.590 579.515 1989.870 579.885 ;
        RECT 1988.740 572.550 1988.880 579.515 ;
        RECT 1988.680 572.230 1988.940 572.550 ;
        RECT 1988.220 524.630 1988.480 524.950 ;
        RECT 1988.280 524.270 1988.420 524.630 ;
        RECT 1988.220 523.950 1988.480 524.270 ;
        RECT 1989.140 523.610 1989.400 523.930 ;
        RECT 1989.200 496.810 1989.340 523.610 ;
        RECT 1988.740 496.670 1989.340 496.810 ;
        RECT 1988.740 400.930 1988.880 496.670 ;
        RECT 1988.280 400.790 1988.880 400.930 ;
        RECT 1988.280 400.250 1988.420 400.790 ;
        RECT 1988.280 400.110 1988.880 400.250 ;
        RECT 1988.740 283.290 1988.880 400.110 ;
        RECT 1988.740 283.150 1989.340 283.290 ;
        RECT 1989.200 282.870 1989.340 283.150 ;
        RECT 1989.140 282.550 1989.400 282.870 ;
        RECT 1988.680 234.610 1988.940 234.930 ;
        RECT 1988.740 110.570 1988.880 234.610 ;
        RECT 1988.280 110.430 1988.880 110.570 ;
        RECT 1988.280 96.550 1988.420 110.430 ;
        RECT 1988.220 96.230 1988.480 96.550 ;
        RECT 1987.760 48.290 1988.020 48.610 ;
        RECT 1987.820 36.710 1987.960 48.290 ;
        RECT 1739.820 36.390 1740.080 36.710 ;
        RECT 1987.760 36.390 1988.020 36.710 ;
        RECT 1739.880 16.650 1740.020 36.390 ;
        RECT 1739.820 16.330 1740.080 16.650 ;
        RECT 1638.160 15.650 1638.420 15.970 ;
        RECT 1638.220 2.400 1638.360 15.650 ;
        RECT 1638.010 -4.800 1638.570 2.400 ;
      LAYER via2 ;
        RECT 1988.670 579.560 1988.950 579.840 ;
        RECT 1989.590 579.560 1989.870 579.840 ;
      LAYER met3 ;
        RECT 1988.645 579.850 1988.975 579.865 ;
        RECT 1989.565 579.850 1989.895 579.865 ;
        RECT 1988.645 579.550 1989.895 579.850 ;
        RECT 1988.645 579.535 1988.975 579.550 ;
        RECT 1989.565 579.535 1989.895 579.550 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1662.510 1690.380 1662.830 1690.440 ;
        RECT 2001.070 1690.380 2001.390 1690.440 ;
        RECT 1662.510 1690.240 2001.390 1690.380 ;
        RECT 1662.510 1690.180 1662.830 1690.240 ;
        RECT 2001.070 1690.180 2001.390 1690.240 ;
        RECT 1656.070 20.640 1656.390 20.700 ;
        RECT 1662.510 20.640 1662.830 20.700 ;
        RECT 1656.070 20.500 1662.830 20.640 ;
        RECT 1656.070 20.440 1656.390 20.500 ;
        RECT 1662.510 20.440 1662.830 20.500 ;
      LAYER via ;
        RECT 1662.540 1690.180 1662.800 1690.440 ;
        RECT 2001.100 1690.180 2001.360 1690.440 ;
        RECT 1656.100 20.440 1656.360 20.700 ;
        RECT 1662.540 20.440 1662.800 20.700 ;
      LAYER met2 ;
        RECT 2001.020 1700.000 2001.300 1704.000 ;
        RECT 2001.160 1690.470 2001.300 1700.000 ;
        RECT 1662.540 1690.150 1662.800 1690.470 ;
        RECT 2001.100 1690.150 2001.360 1690.470 ;
        RECT 1662.600 20.730 1662.740 1690.150 ;
        RECT 1656.100 20.410 1656.360 20.730 ;
        RECT 1662.540 20.410 1662.800 20.730 ;
        RECT 1656.160 2.400 1656.300 20.410 ;
        RECT 1655.950 -4.800 1656.510 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1673.550 44.780 1673.870 44.840 ;
        RECT 2008.430 44.780 2008.750 44.840 ;
        RECT 1673.550 44.640 2008.750 44.780 ;
        RECT 1673.550 44.580 1673.870 44.640 ;
        RECT 2008.430 44.580 2008.750 44.640 ;
      LAYER via ;
        RECT 1673.580 44.580 1673.840 44.840 ;
        RECT 2008.460 44.580 2008.720 44.840 ;
      LAYER met2 ;
        RECT 2010.220 1700.410 2010.500 1704.000 ;
        RECT 2008.520 1700.270 2010.500 1700.410 ;
        RECT 2008.520 44.870 2008.660 1700.270 ;
        RECT 2010.220 1700.000 2010.500 1700.270 ;
        RECT 1673.580 44.550 1673.840 44.870 ;
        RECT 2008.460 44.550 2008.720 44.870 ;
        RECT 1673.640 2.400 1673.780 44.550 ;
        RECT 1673.430 -4.800 1673.990 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1738.945 1684.785 1739.115 1685.975 ;
        RECT 1786.785 1684.785 1786.955 1686.655 ;
        RECT 1835.545 1683.425 1835.715 1686.655 ;
        RECT 1897.185 1683.765 1897.355 1686.655 ;
        RECT 1932.145 1686.485 1932.315 1687.675 ;
        RECT 1945.025 1687.505 1945.195 1689.375 ;
        RECT 1993.785 1686.485 1993.955 1689.715 ;
      LAYER mcon ;
        RECT 1993.785 1689.545 1993.955 1689.715 ;
        RECT 1945.025 1689.205 1945.195 1689.375 ;
        RECT 1932.145 1687.505 1932.315 1687.675 ;
        RECT 1786.785 1686.485 1786.955 1686.655 ;
        RECT 1738.945 1685.805 1739.115 1685.975 ;
        RECT 1835.545 1686.485 1835.715 1686.655 ;
        RECT 1897.185 1686.485 1897.355 1686.655 ;
      LAYER met1 ;
        RECT 1993.725 1689.700 1994.015 1689.745 ;
        RECT 1949.180 1689.560 1994.015 1689.700 ;
        RECT 1944.965 1689.360 1945.255 1689.405 ;
        RECT 1949.180 1689.360 1949.320 1689.560 ;
        RECT 1993.725 1689.515 1994.015 1689.560 ;
        RECT 1944.965 1689.220 1949.320 1689.360 ;
        RECT 1944.965 1689.175 1945.255 1689.220 ;
        RECT 1932.085 1687.660 1932.375 1687.705 ;
        RECT 1944.965 1687.660 1945.255 1687.705 ;
        RECT 1932.085 1687.520 1945.255 1687.660 ;
        RECT 1932.085 1687.475 1932.375 1687.520 ;
        RECT 1944.965 1687.475 1945.255 1687.520 ;
        RECT 1786.725 1686.640 1787.015 1686.685 ;
        RECT 1835.485 1686.640 1835.775 1686.685 ;
        RECT 1786.725 1686.500 1835.775 1686.640 ;
        RECT 1786.725 1686.455 1787.015 1686.500 ;
        RECT 1835.485 1686.455 1835.775 1686.500 ;
        RECT 1897.125 1686.640 1897.415 1686.685 ;
        RECT 1932.085 1686.640 1932.375 1686.685 ;
        RECT 1897.125 1686.500 1932.375 1686.640 ;
        RECT 1897.125 1686.455 1897.415 1686.500 ;
        RECT 1932.085 1686.455 1932.375 1686.500 ;
        RECT 1993.725 1686.640 1994.015 1686.685 ;
        RECT 2019.470 1686.640 2019.790 1686.700 ;
        RECT 1993.725 1686.500 2019.790 1686.640 ;
        RECT 1993.725 1686.455 1994.015 1686.500 ;
        RECT 2019.470 1686.440 2019.790 1686.500 ;
        RECT 1697.010 1686.300 1697.330 1686.360 ;
        RECT 1697.010 1686.160 1728.520 1686.300 ;
        RECT 1697.010 1686.100 1697.330 1686.160 ;
        RECT 1728.380 1685.960 1728.520 1686.160 ;
        RECT 1738.885 1685.960 1739.175 1686.005 ;
        RECT 1728.380 1685.820 1739.175 1685.960 ;
        RECT 1738.885 1685.775 1739.175 1685.820 ;
        RECT 1738.885 1684.940 1739.175 1684.985 ;
        RECT 1786.725 1684.940 1787.015 1684.985 ;
        RECT 1738.885 1684.800 1787.015 1684.940 ;
        RECT 1738.885 1684.755 1739.175 1684.800 ;
        RECT 1786.725 1684.755 1787.015 1684.800 ;
        RECT 1897.125 1683.920 1897.415 1683.965 ;
        RECT 1885.700 1683.780 1897.415 1683.920 ;
        RECT 1835.485 1683.580 1835.775 1683.625 ;
        RECT 1885.700 1683.580 1885.840 1683.780 ;
        RECT 1897.125 1683.735 1897.415 1683.780 ;
        RECT 1835.485 1683.440 1885.840 1683.580 ;
        RECT 1835.485 1683.395 1835.775 1683.440 ;
        RECT 1691.490 15.200 1691.810 15.260 ;
        RECT 1697.010 15.200 1697.330 15.260 ;
        RECT 1691.490 15.060 1697.330 15.200 ;
        RECT 1691.490 15.000 1691.810 15.060 ;
        RECT 1697.010 15.000 1697.330 15.060 ;
      LAYER via ;
        RECT 2019.500 1686.440 2019.760 1686.700 ;
        RECT 1697.040 1686.100 1697.300 1686.360 ;
        RECT 1691.520 15.000 1691.780 15.260 ;
        RECT 1697.040 15.000 1697.300 15.260 ;
      LAYER met2 ;
        RECT 2019.420 1700.000 2019.700 1704.000 ;
        RECT 2019.560 1686.730 2019.700 1700.000 ;
        RECT 2019.500 1686.410 2019.760 1686.730 ;
        RECT 1697.040 1686.070 1697.300 1686.390 ;
        RECT 1697.100 15.290 1697.240 1686.070 ;
        RECT 1691.520 14.970 1691.780 15.290 ;
        RECT 1697.040 14.970 1697.300 15.290 ;
        RECT 1691.580 2.400 1691.720 14.970 ;
        RECT 1691.370 -4.800 1691.930 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1518.070 1678.140 1518.390 1678.200 ;
        RECT 1521.750 1678.140 1522.070 1678.200 ;
        RECT 1518.070 1678.000 1522.070 1678.140 ;
        RECT 1518.070 1677.940 1518.390 1678.000 ;
        RECT 1521.750 1677.940 1522.070 1678.000 ;
        RECT 731.010 66.540 731.330 66.600 ;
        RECT 1518.070 66.540 1518.390 66.600 ;
        RECT 731.010 66.400 1518.390 66.540 ;
        RECT 731.010 66.340 731.330 66.400 ;
        RECT 1518.070 66.340 1518.390 66.400 ;
      LAYER via ;
        RECT 1518.100 1677.940 1518.360 1678.200 ;
        RECT 1521.780 1677.940 1522.040 1678.200 ;
        RECT 731.040 66.340 731.300 66.600 ;
        RECT 1518.100 66.340 1518.360 66.600 ;
      LAYER met2 ;
        RECT 1523.080 1700.410 1523.360 1704.000 ;
        RECT 1521.840 1700.270 1523.360 1700.410 ;
        RECT 1521.840 1678.230 1521.980 1700.270 ;
        RECT 1523.080 1700.000 1523.360 1700.270 ;
        RECT 1518.100 1677.910 1518.360 1678.230 ;
        RECT 1521.780 1677.910 1522.040 1678.230 ;
        RECT 1518.160 66.630 1518.300 1677.910 ;
        RECT 731.040 66.310 731.300 66.630 ;
        RECT 1518.100 66.310 1518.360 66.630 ;
        RECT 731.100 16.730 731.240 66.310 ;
        RECT 728.340 16.590 731.240 16.730 ;
        RECT 728.340 2.400 728.480 16.590 ;
        RECT 728.130 -4.800 728.690 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1759.110 37.980 1759.430 38.040 ;
        RECT 2029.130 37.980 2029.450 38.040 ;
        RECT 1759.110 37.840 2029.450 37.980 ;
        RECT 1759.110 37.780 1759.430 37.840 ;
        RECT 2029.130 37.780 2029.450 37.840 ;
        RECT 1709.430 14.860 1709.750 14.920 ;
        RECT 1759.110 14.860 1759.430 14.920 ;
        RECT 1709.430 14.720 1759.430 14.860 ;
        RECT 1709.430 14.660 1709.750 14.720 ;
        RECT 1759.110 14.660 1759.430 14.720 ;
      LAYER via ;
        RECT 1759.140 37.780 1759.400 38.040 ;
        RECT 2029.160 37.780 2029.420 38.040 ;
        RECT 1709.460 14.660 1709.720 14.920 ;
        RECT 1759.140 14.660 1759.400 14.920 ;
      LAYER met2 ;
        RECT 2028.620 1700.410 2028.900 1704.000 ;
        RECT 2028.620 1700.270 2029.360 1700.410 ;
        RECT 2028.620 1700.000 2028.900 1700.270 ;
        RECT 2029.220 38.070 2029.360 1700.270 ;
        RECT 1759.140 37.750 1759.400 38.070 ;
        RECT 2029.160 37.750 2029.420 38.070 ;
        RECT 1759.200 14.950 1759.340 37.750 ;
        RECT 1709.460 14.630 1709.720 14.950 ;
        RECT 1759.140 14.630 1759.400 14.950 ;
        RECT 1709.520 2.400 1709.660 14.630 ;
        RECT 1709.310 -4.800 1709.870 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1731.510 1686.300 1731.830 1686.360 ;
        RECT 2037.410 1686.300 2037.730 1686.360 ;
        RECT 1731.510 1686.160 2037.730 1686.300 ;
        RECT 1731.510 1686.100 1731.830 1686.160 ;
        RECT 2037.410 1686.100 2037.730 1686.160 ;
        RECT 1731.050 380.020 1731.370 380.080 ;
        RECT 1731.050 379.880 1731.740 380.020 ;
        RECT 1731.050 379.820 1731.370 379.880 ;
        RECT 1731.600 379.740 1731.740 379.880 ;
        RECT 1731.510 379.480 1731.830 379.740 ;
        RECT 1727.370 3.640 1727.690 3.700 ;
        RECT 1731.510 3.640 1731.830 3.700 ;
        RECT 1727.370 3.500 1731.830 3.640 ;
        RECT 1727.370 3.440 1727.690 3.500 ;
        RECT 1731.510 3.440 1731.830 3.500 ;
      LAYER via ;
        RECT 1731.540 1686.100 1731.800 1686.360 ;
        RECT 2037.440 1686.100 2037.700 1686.360 ;
        RECT 1731.080 379.820 1731.340 380.080 ;
        RECT 1731.540 379.480 1731.800 379.740 ;
        RECT 1727.400 3.440 1727.660 3.700 ;
        RECT 1731.540 3.440 1731.800 3.700 ;
      LAYER met2 ;
        RECT 2037.360 1700.000 2037.640 1704.000 ;
        RECT 2037.500 1686.390 2037.640 1700.000 ;
        RECT 1731.540 1686.070 1731.800 1686.390 ;
        RECT 2037.440 1686.070 2037.700 1686.390 ;
        RECT 1731.600 382.570 1731.740 1686.070 ;
        RECT 1731.140 382.430 1731.740 382.570 ;
        RECT 1731.140 380.110 1731.280 382.430 ;
        RECT 1731.080 379.790 1731.340 380.110 ;
        RECT 1731.540 379.450 1731.800 379.770 ;
        RECT 1731.600 3.730 1731.740 379.450 ;
        RECT 1727.400 3.410 1727.660 3.730 ;
        RECT 1731.540 3.410 1731.800 3.730 ;
        RECT 1727.460 2.400 1727.600 3.410 ;
        RECT 1727.250 -4.800 1727.810 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2043.925 1510.365 2044.095 1579.895 ;
        RECT 2043.465 1393.745 2043.635 1441.855 ;
        RECT 2043.925 1062.585 2044.095 1076.695 ;
        RECT 2043.465 524.365 2043.635 572.475 ;
        RECT 2043.925 448.205 2044.095 500.395 ;
        RECT 2043.465 379.865 2043.635 427.635 ;
        RECT 2043.465 331.245 2043.635 379.355 ;
      LAYER mcon ;
        RECT 2043.925 1579.725 2044.095 1579.895 ;
        RECT 2043.465 1441.685 2043.635 1441.855 ;
        RECT 2043.925 1076.525 2044.095 1076.695 ;
        RECT 2043.465 572.305 2043.635 572.475 ;
        RECT 2043.925 500.225 2044.095 500.395 ;
        RECT 2043.465 427.465 2043.635 427.635 ;
        RECT 2043.465 379.185 2043.635 379.355 ;
      LAYER met1 ;
        RECT 2043.390 1607.900 2043.710 1608.160 ;
        RECT 2043.480 1607.420 2043.620 1607.900 ;
        RECT 2043.850 1607.420 2044.170 1607.480 ;
        RECT 2043.480 1607.280 2044.170 1607.420 ;
        RECT 2043.850 1607.220 2044.170 1607.280 ;
        RECT 2043.850 1579.880 2044.170 1579.940 ;
        RECT 2043.655 1579.740 2044.170 1579.880 ;
        RECT 2043.850 1579.680 2044.170 1579.740 ;
        RECT 2043.850 1510.520 2044.170 1510.580 ;
        RECT 2043.655 1510.380 2044.170 1510.520 ;
        RECT 2043.850 1510.320 2044.170 1510.380 ;
        RECT 2043.850 1463.260 2044.170 1463.320 ;
        RECT 2043.480 1463.120 2044.170 1463.260 ;
        RECT 2043.480 1462.640 2043.620 1463.120 ;
        RECT 2043.850 1463.060 2044.170 1463.120 ;
        RECT 2043.390 1462.380 2043.710 1462.640 ;
        RECT 2043.390 1441.840 2043.710 1441.900 ;
        RECT 2043.195 1441.700 2043.710 1441.840 ;
        RECT 2043.390 1441.640 2043.710 1441.700 ;
        RECT 2043.405 1393.900 2043.695 1393.945 ;
        RECT 2043.850 1393.900 2044.170 1393.960 ;
        RECT 2043.405 1393.760 2044.170 1393.900 ;
        RECT 2043.405 1393.715 2043.695 1393.760 ;
        RECT 2043.850 1393.700 2044.170 1393.760 ;
        RECT 2043.850 1366.700 2044.170 1366.760 ;
        RECT 2043.480 1366.560 2044.170 1366.700 ;
        RECT 2043.480 1366.080 2043.620 1366.560 ;
        RECT 2043.850 1366.500 2044.170 1366.560 ;
        RECT 2043.390 1365.820 2043.710 1366.080 ;
        RECT 2043.390 1317.880 2043.710 1318.140 ;
        RECT 2043.480 1317.400 2043.620 1317.880 ;
        RECT 2043.850 1317.400 2044.170 1317.460 ;
        RECT 2043.480 1317.260 2044.170 1317.400 ;
        RECT 2043.850 1317.200 2044.170 1317.260 ;
        RECT 2043.850 1290.200 2044.170 1290.260 ;
        RECT 2044.770 1290.200 2045.090 1290.260 ;
        RECT 2043.850 1290.060 2045.090 1290.200 ;
        RECT 2043.850 1290.000 2044.170 1290.060 ;
        RECT 2044.770 1290.000 2045.090 1290.060 ;
        RECT 2043.390 1124.620 2043.710 1124.680 ;
        RECT 2044.310 1124.620 2044.630 1124.680 ;
        RECT 2043.390 1124.480 2044.630 1124.620 ;
        RECT 2043.390 1124.420 2043.710 1124.480 ;
        RECT 2044.310 1124.420 2044.630 1124.480 ;
        RECT 2043.850 1076.680 2044.170 1076.740 ;
        RECT 2043.655 1076.540 2044.170 1076.680 ;
        RECT 2043.850 1076.480 2044.170 1076.540 ;
        RECT 2043.850 1062.740 2044.170 1062.800 ;
        RECT 2043.655 1062.600 2044.170 1062.740 ;
        RECT 2043.850 1062.540 2044.170 1062.600 ;
        RECT 2043.850 966.180 2044.170 966.240 ;
        RECT 2044.770 966.180 2045.090 966.240 ;
        RECT 2043.850 966.040 2045.090 966.180 ;
        RECT 2043.850 965.980 2044.170 966.040 ;
        RECT 2044.770 965.980 2045.090 966.040 ;
        RECT 2043.850 869.620 2044.170 869.680 ;
        RECT 2044.770 869.620 2045.090 869.680 ;
        RECT 2043.850 869.480 2045.090 869.620 ;
        RECT 2043.850 869.420 2044.170 869.480 ;
        RECT 2044.770 869.420 2045.090 869.480 ;
        RECT 2042.010 821.000 2042.330 821.060 ;
        RECT 2042.930 821.000 2043.250 821.060 ;
        RECT 2042.010 820.860 2043.250 821.000 ;
        RECT 2042.010 820.800 2042.330 820.860 ;
        RECT 2042.930 820.800 2043.250 820.860 ;
        RECT 2044.310 700.300 2044.630 700.360 ;
        RECT 2045.230 700.300 2045.550 700.360 ;
        RECT 2044.310 700.160 2045.550 700.300 ;
        RECT 2044.310 700.100 2044.630 700.160 ;
        RECT 2045.230 700.100 2045.550 700.160 ;
        RECT 2042.930 573.140 2043.250 573.200 ;
        RECT 2043.850 573.140 2044.170 573.200 ;
        RECT 2042.930 573.000 2044.170 573.140 ;
        RECT 2042.930 572.940 2043.250 573.000 ;
        RECT 2043.850 572.940 2044.170 573.000 ;
        RECT 2043.405 572.460 2043.695 572.505 ;
        RECT 2043.850 572.460 2044.170 572.520 ;
        RECT 2043.405 572.320 2044.170 572.460 ;
        RECT 2043.405 572.275 2043.695 572.320 ;
        RECT 2043.850 572.260 2044.170 572.320 ;
        RECT 2043.390 524.520 2043.710 524.580 ;
        RECT 2043.195 524.380 2043.710 524.520 ;
        RECT 2043.390 524.320 2043.710 524.380 ;
        RECT 2043.850 500.380 2044.170 500.440 ;
        RECT 2043.655 500.240 2044.170 500.380 ;
        RECT 2043.850 500.180 2044.170 500.240 ;
        RECT 2043.850 448.360 2044.170 448.420 ;
        RECT 2043.655 448.220 2044.170 448.360 ;
        RECT 2043.850 448.160 2044.170 448.220 ;
        RECT 2043.405 427.620 2043.695 427.665 ;
        RECT 2044.310 427.620 2044.630 427.680 ;
        RECT 2043.405 427.480 2044.630 427.620 ;
        RECT 2043.405 427.435 2043.695 427.480 ;
        RECT 2044.310 427.420 2044.630 427.480 ;
        RECT 2043.390 380.020 2043.710 380.080 ;
        RECT 2043.195 379.880 2043.710 380.020 ;
        RECT 2043.390 379.820 2043.710 379.880 ;
        RECT 2043.390 379.340 2043.710 379.400 ;
        RECT 2043.195 379.200 2043.710 379.340 ;
        RECT 2043.390 379.140 2043.710 379.200 ;
        RECT 2043.405 331.400 2043.695 331.445 ;
        RECT 2043.850 331.400 2044.170 331.460 ;
        RECT 2043.405 331.260 2044.170 331.400 ;
        RECT 2043.405 331.215 2043.695 331.260 ;
        RECT 2043.850 331.200 2044.170 331.260 ;
        RECT 2043.390 255.580 2043.710 255.640 ;
        RECT 2043.390 255.440 2044.080 255.580 ;
        RECT 2043.390 255.380 2043.710 255.440 ;
        RECT 2043.940 255.300 2044.080 255.440 ;
        RECT 2043.850 255.040 2044.170 255.300 ;
        RECT 2043.390 227.700 2043.710 227.760 ;
        RECT 2043.850 227.700 2044.170 227.760 ;
        RECT 2043.390 227.560 2044.170 227.700 ;
        RECT 2043.390 227.500 2043.710 227.560 ;
        RECT 2043.850 227.500 2044.170 227.560 ;
        RECT 2043.850 159.020 2044.170 159.080 ;
        RECT 2043.480 158.880 2044.170 159.020 ;
        RECT 2043.480 158.740 2043.620 158.880 ;
        RECT 2043.850 158.820 2044.170 158.880 ;
        RECT 2043.390 158.480 2043.710 158.740 ;
        RECT 1745.310 34.240 1745.630 34.300 ;
        RECT 2043.850 34.240 2044.170 34.300 ;
        RECT 1745.310 34.100 2044.170 34.240 ;
        RECT 1745.310 34.040 1745.630 34.100 ;
        RECT 2043.850 34.040 2044.170 34.100 ;
      LAYER via ;
        RECT 2043.420 1607.900 2043.680 1608.160 ;
        RECT 2043.880 1607.220 2044.140 1607.480 ;
        RECT 2043.880 1579.680 2044.140 1579.940 ;
        RECT 2043.880 1510.320 2044.140 1510.580 ;
        RECT 2043.880 1463.060 2044.140 1463.320 ;
        RECT 2043.420 1462.380 2043.680 1462.640 ;
        RECT 2043.420 1441.640 2043.680 1441.900 ;
        RECT 2043.880 1393.700 2044.140 1393.960 ;
        RECT 2043.880 1366.500 2044.140 1366.760 ;
        RECT 2043.420 1365.820 2043.680 1366.080 ;
        RECT 2043.420 1317.880 2043.680 1318.140 ;
        RECT 2043.880 1317.200 2044.140 1317.460 ;
        RECT 2043.880 1290.000 2044.140 1290.260 ;
        RECT 2044.800 1290.000 2045.060 1290.260 ;
        RECT 2043.420 1124.420 2043.680 1124.680 ;
        RECT 2044.340 1124.420 2044.600 1124.680 ;
        RECT 2043.880 1076.480 2044.140 1076.740 ;
        RECT 2043.880 1062.540 2044.140 1062.800 ;
        RECT 2043.880 965.980 2044.140 966.240 ;
        RECT 2044.800 965.980 2045.060 966.240 ;
        RECT 2043.880 869.420 2044.140 869.680 ;
        RECT 2044.800 869.420 2045.060 869.680 ;
        RECT 2042.040 820.800 2042.300 821.060 ;
        RECT 2042.960 820.800 2043.220 821.060 ;
        RECT 2044.340 700.100 2044.600 700.360 ;
        RECT 2045.260 700.100 2045.520 700.360 ;
        RECT 2042.960 572.940 2043.220 573.200 ;
        RECT 2043.880 572.940 2044.140 573.200 ;
        RECT 2043.880 572.260 2044.140 572.520 ;
        RECT 2043.420 524.320 2043.680 524.580 ;
        RECT 2043.880 500.180 2044.140 500.440 ;
        RECT 2043.880 448.160 2044.140 448.420 ;
        RECT 2044.340 427.420 2044.600 427.680 ;
        RECT 2043.420 379.820 2043.680 380.080 ;
        RECT 2043.420 379.140 2043.680 379.400 ;
        RECT 2043.880 331.200 2044.140 331.460 ;
        RECT 2043.420 255.380 2043.680 255.640 ;
        RECT 2043.880 255.040 2044.140 255.300 ;
        RECT 2043.420 227.500 2043.680 227.760 ;
        RECT 2043.880 227.500 2044.140 227.760 ;
        RECT 2043.880 158.820 2044.140 159.080 ;
        RECT 2043.420 158.480 2043.680 158.740 ;
        RECT 1745.340 34.040 1745.600 34.300 ;
        RECT 2043.880 34.040 2044.140 34.300 ;
      LAYER met2 ;
        RECT 2046.560 1701.090 2046.840 1704.000 ;
        RECT 2044.400 1700.950 2046.840 1701.090 ;
        RECT 2044.400 1656.210 2044.540 1700.950 ;
        RECT 2046.560 1700.000 2046.840 1700.950 ;
        RECT 2043.480 1656.070 2044.540 1656.210 ;
        RECT 2043.480 1608.190 2043.620 1656.070 ;
        RECT 2043.420 1607.870 2043.680 1608.190 ;
        RECT 2043.880 1607.190 2044.140 1607.510 ;
        RECT 2043.940 1579.970 2044.080 1607.190 ;
        RECT 2043.880 1579.650 2044.140 1579.970 ;
        RECT 2043.880 1510.290 2044.140 1510.610 ;
        RECT 2043.940 1463.350 2044.080 1510.290 ;
        RECT 2043.880 1463.030 2044.140 1463.350 ;
        RECT 2043.420 1462.350 2043.680 1462.670 ;
        RECT 2043.480 1441.930 2043.620 1462.350 ;
        RECT 2043.420 1441.610 2043.680 1441.930 ;
        RECT 2043.880 1393.670 2044.140 1393.990 ;
        RECT 2043.940 1366.790 2044.080 1393.670 ;
        RECT 2043.880 1366.470 2044.140 1366.790 ;
        RECT 2043.420 1365.790 2043.680 1366.110 ;
        RECT 2043.480 1318.170 2043.620 1365.790 ;
        RECT 2043.420 1317.850 2043.680 1318.170 ;
        RECT 2043.880 1317.170 2044.140 1317.490 ;
        RECT 2043.940 1290.290 2044.080 1317.170 ;
        RECT 2043.880 1289.970 2044.140 1290.290 ;
        RECT 2044.800 1289.970 2045.060 1290.290 ;
        RECT 2044.860 1242.205 2045.000 1289.970 ;
        RECT 2043.870 1241.835 2044.150 1242.205 ;
        RECT 2044.790 1241.835 2045.070 1242.205 ;
        RECT 2043.940 1145.530 2044.080 1241.835 ;
        RECT 2043.480 1145.390 2044.080 1145.530 ;
        RECT 2043.480 1124.710 2043.620 1145.390 ;
        RECT 2043.420 1124.390 2043.680 1124.710 ;
        RECT 2044.340 1124.390 2044.600 1124.710 ;
        RECT 2044.400 1110.850 2044.540 1124.390 ;
        RECT 2043.940 1110.710 2044.540 1110.850 ;
        RECT 2043.940 1076.770 2044.080 1110.710 ;
        RECT 2043.880 1076.450 2044.140 1076.770 ;
        RECT 2043.880 1062.510 2044.140 1062.830 ;
        RECT 2043.940 1027.890 2044.080 1062.510 ;
        RECT 2043.480 1027.750 2044.080 1027.890 ;
        RECT 2043.480 1014.405 2043.620 1027.750 ;
        RECT 2043.410 1014.035 2043.690 1014.405 ;
        RECT 2044.790 1014.035 2045.070 1014.405 ;
        RECT 2044.860 966.270 2045.000 1014.035 ;
        RECT 2043.880 965.950 2044.140 966.270 ;
        RECT 2044.800 965.950 2045.060 966.270 ;
        RECT 2043.940 931.330 2044.080 965.950 ;
        RECT 2043.480 931.190 2044.080 931.330 ;
        RECT 2043.480 917.845 2043.620 931.190 ;
        RECT 2043.410 917.475 2043.690 917.845 ;
        RECT 2044.790 917.475 2045.070 917.845 ;
        RECT 2044.860 869.710 2045.000 917.475 ;
        RECT 2043.880 869.390 2044.140 869.710 ;
        RECT 2044.800 869.390 2045.060 869.710 ;
        RECT 2043.940 834.770 2044.080 869.390 ;
        RECT 2043.020 834.630 2044.080 834.770 ;
        RECT 2043.020 821.090 2043.160 834.630 ;
        RECT 2042.040 820.770 2042.300 821.090 ;
        RECT 2042.960 820.770 2043.220 821.090 ;
        RECT 2042.100 773.005 2042.240 820.770 ;
        RECT 2042.030 772.635 2042.310 773.005 ;
        RECT 2043.410 772.635 2043.690 773.005 ;
        RECT 2043.480 738.210 2043.620 772.635 ;
        RECT 2043.480 738.070 2044.540 738.210 ;
        RECT 2044.400 700.390 2044.540 738.070 ;
        RECT 2044.340 700.070 2044.600 700.390 ;
        RECT 2045.260 700.070 2045.520 700.390 ;
        RECT 2045.320 676.445 2045.460 700.070 ;
        RECT 2044.330 676.075 2044.610 676.445 ;
        RECT 2045.250 676.075 2045.530 676.445 ;
        RECT 2044.400 628.845 2044.540 676.075 ;
        RECT 2044.330 628.475 2044.610 628.845 ;
        RECT 2043.410 627.795 2043.690 628.165 ;
        RECT 2043.480 596.770 2043.620 627.795 ;
        RECT 2043.020 596.630 2043.620 596.770 ;
        RECT 2043.020 573.230 2043.160 596.630 ;
        RECT 2042.960 572.910 2043.220 573.230 ;
        RECT 2043.880 572.910 2044.140 573.230 ;
        RECT 2043.940 572.550 2044.080 572.910 ;
        RECT 2043.880 572.230 2044.140 572.550 ;
        RECT 2043.420 524.290 2043.680 524.610 ;
        RECT 2043.480 524.010 2043.620 524.290 ;
        RECT 2043.480 523.870 2044.080 524.010 ;
        RECT 2043.940 500.470 2044.080 523.870 ;
        RECT 2043.880 500.150 2044.140 500.470 ;
        RECT 2043.880 448.130 2044.140 448.450 ;
        RECT 2043.940 434.930 2044.080 448.130 ;
        RECT 2043.940 434.790 2044.540 434.930 ;
        RECT 2044.400 427.710 2044.540 434.790 ;
        RECT 2044.340 427.390 2044.600 427.710 ;
        RECT 2043.420 379.790 2043.680 380.110 ;
        RECT 2043.480 379.430 2043.620 379.790 ;
        RECT 2043.420 379.110 2043.680 379.430 ;
        RECT 2043.880 331.170 2044.140 331.490 ;
        RECT 2043.940 330.890 2044.080 331.170 ;
        RECT 2043.480 330.750 2044.080 330.890 ;
        RECT 2043.480 303.690 2043.620 330.750 ;
        RECT 2043.480 303.550 2044.080 303.690 ;
        RECT 2043.940 283.290 2044.080 303.550 ;
        RECT 2043.480 283.150 2044.080 283.290 ;
        RECT 2043.480 255.670 2043.620 283.150 ;
        RECT 2043.420 255.350 2043.680 255.670 ;
        RECT 2043.880 255.010 2044.140 255.330 ;
        RECT 2043.940 235.010 2044.080 255.010 ;
        RECT 2043.480 234.870 2044.080 235.010 ;
        RECT 2043.480 227.790 2043.620 234.870 ;
        RECT 2043.420 227.470 2043.680 227.790 ;
        RECT 2043.880 227.470 2044.140 227.790 ;
        RECT 2043.940 159.110 2044.080 227.470 ;
        RECT 2043.880 158.790 2044.140 159.110 ;
        RECT 2043.420 158.450 2043.680 158.770 ;
        RECT 2043.480 137.885 2043.620 158.450 ;
        RECT 2043.410 137.515 2043.690 137.885 ;
        RECT 2043.870 136.835 2044.150 137.205 ;
        RECT 2043.940 34.330 2044.080 136.835 ;
        RECT 1745.340 34.010 1745.600 34.330 ;
        RECT 2043.880 34.010 2044.140 34.330 ;
        RECT 1745.400 2.400 1745.540 34.010 ;
        RECT 1745.190 -4.800 1745.750 2.400 ;
      LAYER via2 ;
        RECT 2043.870 1241.880 2044.150 1242.160 ;
        RECT 2044.790 1241.880 2045.070 1242.160 ;
        RECT 2043.410 1014.080 2043.690 1014.360 ;
        RECT 2044.790 1014.080 2045.070 1014.360 ;
        RECT 2043.410 917.520 2043.690 917.800 ;
        RECT 2044.790 917.520 2045.070 917.800 ;
        RECT 2042.030 772.680 2042.310 772.960 ;
        RECT 2043.410 772.680 2043.690 772.960 ;
        RECT 2044.330 676.120 2044.610 676.400 ;
        RECT 2045.250 676.120 2045.530 676.400 ;
        RECT 2044.330 628.520 2044.610 628.800 ;
        RECT 2043.410 627.840 2043.690 628.120 ;
        RECT 2043.410 137.560 2043.690 137.840 ;
        RECT 2043.870 136.880 2044.150 137.160 ;
      LAYER met3 ;
        RECT 2043.845 1242.170 2044.175 1242.185 ;
        RECT 2044.765 1242.170 2045.095 1242.185 ;
        RECT 2043.845 1241.870 2045.095 1242.170 ;
        RECT 2043.845 1241.855 2044.175 1241.870 ;
        RECT 2044.765 1241.855 2045.095 1241.870 ;
        RECT 2043.385 1014.370 2043.715 1014.385 ;
        RECT 2044.765 1014.370 2045.095 1014.385 ;
        RECT 2043.385 1014.070 2045.095 1014.370 ;
        RECT 2043.385 1014.055 2043.715 1014.070 ;
        RECT 2044.765 1014.055 2045.095 1014.070 ;
        RECT 2043.385 917.810 2043.715 917.825 ;
        RECT 2044.765 917.810 2045.095 917.825 ;
        RECT 2043.385 917.510 2045.095 917.810 ;
        RECT 2043.385 917.495 2043.715 917.510 ;
        RECT 2044.765 917.495 2045.095 917.510 ;
        RECT 2042.005 772.970 2042.335 772.985 ;
        RECT 2043.385 772.970 2043.715 772.985 ;
        RECT 2042.005 772.670 2043.715 772.970 ;
        RECT 2042.005 772.655 2042.335 772.670 ;
        RECT 2043.385 772.655 2043.715 772.670 ;
        RECT 2044.305 676.410 2044.635 676.425 ;
        RECT 2045.225 676.410 2045.555 676.425 ;
        RECT 2044.305 676.110 2045.555 676.410 ;
        RECT 2044.305 676.095 2044.635 676.110 ;
        RECT 2045.225 676.095 2045.555 676.110 ;
        RECT 2044.305 628.810 2044.635 628.825 ;
        RECT 2042.710 628.510 2044.635 628.810 ;
        RECT 2042.710 628.130 2043.010 628.510 ;
        RECT 2044.305 628.495 2044.635 628.510 ;
        RECT 2043.385 628.130 2043.715 628.145 ;
        RECT 2042.710 627.830 2043.715 628.130 ;
        RECT 2043.385 627.815 2043.715 627.830 ;
        RECT 2043.385 137.850 2043.715 137.865 ;
        RECT 2042.710 137.550 2043.715 137.850 ;
        RECT 2042.710 137.170 2043.010 137.550 ;
        RECT 2043.385 137.535 2043.715 137.550 ;
        RECT 2043.845 137.170 2044.175 137.185 ;
        RECT 2042.710 136.870 2044.175 137.170 ;
        RECT 2043.845 136.855 2044.175 136.870 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1994.245 1685.805 1994.415 1689.375 ;
        RECT 2020.005 1686.485 2020.175 1689.375 ;
      LAYER mcon ;
        RECT 1994.245 1689.205 1994.415 1689.375 ;
        RECT 2020.005 1689.205 2020.175 1689.375 ;
      LAYER met1 ;
        RECT 1994.185 1689.360 1994.475 1689.405 ;
        RECT 2019.945 1689.360 2020.235 1689.405 ;
        RECT 1994.185 1689.220 2020.235 1689.360 ;
        RECT 1994.185 1689.175 1994.475 1689.220 ;
        RECT 2019.945 1689.175 2020.235 1689.220 ;
        RECT 2019.945 1686.640 2020.235 1686.685 ;
        RECT 2055.810 1686.640 2056.130 1686.700 ;
        RECT 2019.945 1686.500 2056.130 1686.640 ;
        RECT 2019.945 1686.455 2020.235 1686.500 ;
        RECT 2055.810 1686.440 2056.130 1686.500 ;
        RECT 1994.185 1685.960 1994.475 1686.005 ;
        RECT 1773.000 1685.820 1994.475 1685.960 ;
        RECT 1766.010 1685.620 1766.330 1685.680 ;
        RECT 1773.000 1685.620 1773.140 1685.820 ;
        RECT 1994.185 1685.775 1994.475 1685.820 ;
        RECT 1766.010 1685.480 1773.140 1685.620 ;
        RECT 1766.010 1685.420 1766.330 1685.480 ;
        RECT 1762.790 18.600 1763.110 18.660 ;
        RECT 1766.010 18.600 1766.330 18.660 ;
        RECT 1762.790 18.460 1766.330 18.600 ;
        RECT 1762.790 18.400 1763.110 18.460 ;
        RECT 1766.010 18.400 1766.330 18.460 ;
      LAYER via ;
        RECT 2055.840 1686.440 2056.100 1686.700 ;
        RECT 1766.040 1685.420 1766.300 1685.680 ;
        RECT 1762.820 18.400 1763.080 18.660 ;
        RECT 1766.040 18.400 1766.300 18.660 ;
      LAYER met2 ;
        RECT 2055.760 1700.000 2056.040 1704.000 ;
        RECT 2055.900 1686.730 2056.040 1700.000 ;
        RECT 2055.840 1686.410 2056.100 1686.730 ;
        RECT 1766.040 1685.390 1766.300 1685.710 ;
        RECT 1766.100 18.690 1766.240 1685.390 ;
        RECT 1762.820 18.370 1763.080 18.690 ;
        RECT 1766.040 18.370 1766.300 18.690 ;
        RECT 1762.880 2.400 1763.020 18.370 ;
        RECT 1762.670 -4.800 1763.230 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2052.590 1683.920 2052.910 1683.980 ;
        RECT 2065.010 1683.920 2065.330 1683.980 ;
        RECT 2052.590 1683.780 2065.330 1683.920 ;
        RECT 2052.590 1683.720 2052.910 1683.780 ;
        RECT 2065.010 1683.720 2065.330 1683.780 ;
      LAYER via ;
        RECT 2052.620 1683.720 2052.880 1683.980 ;
        RECT 2065.040 1683.720 2065.300 1683.980 ;
      LAYER met2 ;
        RECT 2064.960 1700.000 2065.240 1704.000 ;
        RECT 2065.100 1684.010 2065.240 1700.000 ;
        RECT 2052.620 1683.690 2052.880 1684.010 ;
        RECT 2065.040 1683.690 2065.300 1684.010 ;
        RECT 2052.680 16.845 2052.820 1683.690 ;
        RECT 1780.750 16.475 1781.030 16.845 ;
        RECT 2052.610 16.475 2052.890 16.845 ;
        RECT 1780.820 2.400 1780.960 16.475 ;
        RECT 1780.610 -4.800 1781.170 2.400 ;
      LAYER via2 ;
        RECT 1780.750 16.520 1781.030 16.800 ;
        RECT 2052.610 16.520 2052.890 16.800 ;
      LAYER met3 ;
        RECT 1780.725 16.810 1781.055 16.825 ;
        RECT 2052.585 16.810 2052.915 16.825 ;
        RECT 1780.725 16.510 2052.915 16.810 ;
        RECT 1780.725 16.495 1781.055 16.510 ;
        RECT 2052.585 16.495 2052.915 16.510 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1800.510 1685.280 1800.830 1685.340 ;
        RECT 2074.210 1685.280 2074.530 1685.340 ;
        RECT 1800.510 1685.140 2074.530 1685.280 ;
        RECT 1800.510 1685.080 1800.830 1685.140 ;
        RECT 2074.210 1685.080 2074.530 1685.140 ;
      LAYER via ;
        RECT 1800.540 1685.080 1800.800 1685.340 ;
        RECT 2074.240 1685.080 2074.500 1685.340 ;
      LAYER met2 ;
        RECT 2074.160 1700.000 2074.440 1704.000 ;
        RECT 2074.300 1685.370 2074.440 1700.000 ;
        RECT 1800.540 1685.050 1800.800 1685.370 ;
        RECT 2074.240 1685.050 2074.500 1685.370 ;
        RECT 1800.600 3.130 1800.740 1685.050 ;
        RECT 1798.760 2.990 1800.740 3.130 ;
        RECT 1798.760 2.400 1798.900 2.990 ;
        RECT 1798.550 -4.800 1799.110 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1857.625 14.705 1857.795 17.255 ;
        RECT 2042.545 15.555 2042.715 16.235 ;
        RECT 2042.545 15.385 2044.095 15.555 ;
      LAYER mcon ;
        RECT 1857.625 17.085 1857.795 17.255 ;
        RECT 2042.545 16.065 2042.715 16.235 ;
        RECT 2043.925 15.385 2044.095 15.555 ;
      LAYER met1 ;
        RECT 2053.050 1684.260 2053.370 1684.320 ;
        RECT 2082.030 1684.260 2082.350 1684.320 ;
        RECT 2053.050 1684.120 2082.350 1684.260 ;
        RECT 2053.050 1684.060 2053.370 1684.120 ;
        RECT 2082.030 1684.060 2082.350 1684.120 ;
        RECT 1857.565 17.240 1857.855 17.285 ;
        RECT 1857.565 17.100 2018.780 17.240 ;
        RECT 1857.565 17.055 1857.855 17.100 ;
        RECT 2018.640 16.900 2018.780 17.100 ;
        RECT 2018.640 16.760 2019.240 16.900 ;
        RECT 2019.100 16.220 2019.240 16.760 ;
        RECT 2042.485 16.220 2042.775 16.265 ;
        RECT 2019.100 16.080 2042.775 16.220 ;
        RECT 2042.485 16.035 2042.775 16.080 ;
        RECT 2043.865 15.540 2044.155 15.585 ;
        RECT 2053.050 15.540 2053.370 15.600 ;
        RECT 2043.865 15.400 2053.370 15.540 ;
        RECT 2043.865 15.355 2044.155 15.400 ;
        RECT 2053.050 15.340 2053.370 15.400 ;
        RECT 1816.610 14.860 1816.930 14.920 ;
        RECT 1857.565 14.860 1857.855 14.905 ;
        RECT 1816.610 14.720 1857.855 14.860 ;
        RECT 1816.610 14.660 1816.930 14.720 ;
        RECT 1857.565 14.675 1857.855 14.720 ;
      LAYER via ;
        RECT 2053.080 1684.060 2053.340 1684.320 ;
        RECT 2082.060 1684.060 2082.320 1684.320 ;
        RECT 2053.080 15.340 2053.340 15.600 ;
        RECT 1816.640 14.660 1816.900 14.920 ;
      LAYER met2 ;
        RECT 2083.360 1700.410 2083.640 1704.000 ;
        RECT 2082.120 1700.270 2083.640 1700.410 ;
        RECT 2082.120 1684.350 2082.260 1700.270 ;
        RECT 2083.360 1700.000 2083.640 1700.270 ;
        RECT 2053.080 1684.030 2053.340 1684.350 ;
        RECT 2082.060 1684.030 2082.320 1684.350 ;
        RECT 2053.140 15.630 2053.280 1684.030 ;
        RECT 2053.080 15.310 2053.340 15.630 ;
        RECT 1816.640 14.630 1816.900 14.950 ;
        RECT 1816.700 2.400 1816.840 14.630 ;
        RECT 1816.490 -4.800 1817.050 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1834.550 1688.340 1834.870 1688.400 ;
        RECT 2092.610 1688.340 2092.930 1688.400 ;
        RECT 1834.550 1688.200 2092.930 1688.340 ;
        RECT 1834.550 1688.140 1834.870 1688.200 ;
        RECT 2092.610 1688.140 2092.930 1688.200 ;
      LAYER via ;
        RECT 1834.580 1688.140 1834.840 1688.400 ;
        RECT 2092.640 1688.140 2092.900 1688.400 ;
      LAYER met2 ;
        RECT 2092.560 1700.000 2092.840 1704.000 ;
        RECT 2092.700 1688.430 2092.840 1700.000 ;
        RECT 1834.580 1688.110 1834.840 1688.430 ;
        RECT 2092.640 1688.110 2092.900 1688.430 ;
        RECT 1834.640 2.400 1834.780 1688.110 ;
        RECT 1834.430 -4.800 1834.990 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2018.165 15.385 2018.335 16.235 ;
      LAYER mcon ;
        RECT 2018.165 16.065 2018.335 16.235 ;
      LAYER met1 ;
        RECT 2101.810 1689.700 2102.130 1689.760 ;
        RECT 2077.980 1689.560 2102.130 1689.700 ;
        RECT 2066.390 1689.360 2066.710 1689.420 ;
        RECT 2077.980 1689.360 2078.120 1689.560 ;
        RECT 2101.810 1689.500 2102.130 1689.560 ;
        RECT 2066.390 1689.220 2078.120 1689.360 ;
        RECT 2066.390 1689.160 2066.710 1689.220 ;
        RECT 1852.030 16.220 1852.350 16.280 ;
        RECT 2018.105 16.220 2018.395 16.265 ;
        RECT 1852.030 16.080 2018.395 16.220 ;
        RECT 1852.030 16.020 1852.350 16.080 ;
        RECT 2018.105 16.035 2018.395 16.080 ;
        RECT 2018.105 15.540 2018.395 15.585 ;
        RECT 2018.105 15.400 2043.620 15.540 ;
        RECT 2018.105 15.355 2018.395 15.400 ;
        RECT 2043.480 15.200 2043.620 15.400 ;
        RECT 2066.390 15.200 2066.710 15.260 ;
        RECT 2043.480 15.060 2066.710 15.200 ;
        RECT 2066.390 15.000 2066.710 15.060 ;
      LAYER via ;
        RECT 2066.420 1689.160 2066.680 1689.420 ;
        RECT 2101.840 1689.500 2102.100 1689.760 ;
        RECT 1852.060 16.020 1852.320 16.280 ;
        RECT 2066.420 15.000 2066.680 15.260 ;
      LAYER met2 ;
        RECT 2101.760 1700.000 2102.040 1704.000 ;
        RECT 2101.900 1689.790 2102.040 1700.000 ;
        RECT 2101.840 1689.470 2102.100 1689.790 ;
        RECT 2066.420 1689.130 2066.680 1689.450 ;
        RECT 1852.060 15.990 1852.320 16.310 ;
        RECT 1852.120 2.400 1852.260 15.990 ;
        RECT 2066.480 15.290 2066.620 1689.130 ;
        RECT 2066.420 14.970 2066.680 15.290 ;
        RECT 1851.910 -4.800 1852.470 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1876.410 1687.320 1876.730 1687.380 ;
        RECT 2111.010 1687.320 2111.330 1687.380 ;
        RECT 1876.410 1687.180 2111.330 1687.320 ;
        RECT 1876.410 1687.120 1876.730 1687.180 ;
        RECT 2111.010 1687.120 2111.330 1687.180 ;
        RECT 1869.970 9.760 1870.290 9.820 ;
        RECT 1876.410 9.760 1876.730 9.820 ;
        RECT 1869.970 9.620 1876.730 9.760 ;
        RECT 1869.970 9.560 1870.290 9.620 ;
        RECT 1876.410 9.560 1876.730 9.620 ;
      LAYER via ;
        RECT 1876.440 1687.120 1876.700 1687.380 ;
        RECT 2111.040 1687.120 2111.300 1687.380 ;
        RECT 1870.000 9.560 1870.260 9.820 ;
        RECT 1876.440 9.560 1876.700 9.820 ;
      LAYER met2 ;
        RECT 2110.960 1700.000 2111.240 1704.000 ;
        RECT 2111.100 1687.410 2111.240 1700.000 ;
        RECT 1876.440 1687.090 1876.700 1687.410 ;
        RECT 2111.040 1687.090 2111.300 1687.410 ;
        RECT 1876.500 9.850 1876.640 1687.090 ;
        RECT 1870.000 9.530 1870.260 9.850 ;
        RECT 1876.440 9.530 1876.700 9.850 ;
        RECT 1870.060 2.400 1870.200 9.530 ;
        RECT 1869.850 -4.800 1870.410 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 751.710 67.560 752.030 67.620 ;
        RECT 1532.330 67.560 1532.650 67.620 ;
        RECT 751.710 67.420 1532.650 67.560 ;
        RECT 751.710 67.360 752.030 67.420 ;
        RECT 1532.330 67.360 1532.650 67.420 ;
      LAYER via ;
        RECT 751.740 67.360 752.000 67.620 ;
        RECT 1532.360 67.360 1532.620 67.620 ;
      LAYER met2 ;
        RECT 1532.280 1700.000 1532.560 1704.000 ;
        RECT 1532.420 67.650 1532.560 1700.000 ;
        RECT 751.740 67.330 752.000 67.650 ;
        RECT 1532.360 67.330 1532.620 67.650 ;
        RECT 751.800 16.730 751.940 67.330 ;
        RECT 746.280 16.590 751.940 16.730 ;
        RECT 746.280 2.400 746.420 16.590 ;
        RECT 746.070 -4.800 746.630 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2067.310 1686.300 2067.630 1686.360 ;
        RECT 2067.310 1686.160 2105.720 1686.300 ;
        RECT 2067.310 1686.100 2067.630 1686.160 ;
        RECT 2105.580 1685.960 2105.720 1686.160 ;
        RECT 2120.210 1685.960 2120.530 1686.020 ;
        RECT 2105.580 1685.820 2120.530 1685.960 ;
        RECT 2120.210 1685.760 2120.530 1685.820 ;
        RECT 1887.910 14.860 1888.230 14.920 ;
        RECT 2067.310 14.860 2067.630 14.920 ;
        RECT 1887.910 14.720 2067.630 14.860 ;
        RECT 1887.910 14.660 1888.230 14.720 ;
        RECT 2067.310 14.660 2067.630 14.720 ;
      LAYER via ;
        RECT 2067.340 1686.100 2067.600 1686.360 ;
        RECT 2120.240 1685.760 2120.500 1686.020 ;
        RECT 1887.940 14.660 1888.200 14.920 ;
        RECT 2067.340 14.660 2067.600 14.920 ;
      LAYER met2 ;
        RECT 2120.160 1700.000 2120.440 1704.000 ;
        RECT 2067.340 1686.070 2067.600 1686.390 ;
        RECT 2067.400 14.950 2067.540 1686.070 ;
        RECT 2120.300 1686.050 2120.440 1700.000 ;
        RECT 2120.240 1685.730 2120.500 1686.050 ;
        RECT 1887.940 14.630 1888.200 14.950 ;
        RECT 2067.340 14.630 2067.600 14.950 ;
        RECT 1888.000 2.400 1888.140 14.630 ;
        RECT 1887.790 -4.800 1888.350 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2121.590 1683.920 2121.910 1683.980 ;
        RECT 2129.410 1683.920 2129.730 1683.980 ;
        RECT 2121.590 1683.780 2129.730 1683.920 ;
        RECT 2121.590 1683.720 2121.910 1683.780 ;
        RECT 2129.410 1683.720 2129.730 1683.780 ;
        RECT 2121.590 16.900 2121.910 16.960 ;
        RECT 2110.640 16.760 2121.910 16.900 ;
        RECT 2110.640 16.220 2110.780 16.760 ;
        RECT 2121.590 16.700 2121.910 16.760 ;
        RECT 2106.040 16.080 2110.780 16.220 ;
        RECT 1905.850 15.880 1906.170 15.940 ;
        RECT 2106.040 15.880 2106.180 16.080 ;
        RECT 1905.850 15.740 2106.180 15.880 ;
        RECT 1905.850 15.680 1906.170 15.740 ;
      LAYER via ;
        RECT 2121.620 1683.720 2121.880 1683.980 ;
        RECT 2129.440 1683.720 2129.700 1683.980 ;
        RECT 2121.620 16.700 2121.880 16.960 ;
        RECT 1905.880 15.680 1906.140 15.940 ;
      LAYER met2 ;
        RECT 2129.360 1700.000 2129.640 1704.000 ;
        RECT 2129.500 1684.010 2129.640 1700.000 ;
        RECT 2121.620 1683.690 2121.880 1684.010 ;
        RECT 2129.440 1683.690 2129.700 1684.010 ;
        RECT 2121.680 16.990 2121.820 1683.690 ;
        RECT 2121.620 16.670 2121.880 16.990 ;
        RECT 1905.880 15.650 1906.140 15.970 ;
        RECT 1905.940 2.400 1906.080 15.650 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2105.105 1684.105 2105.275 1685.975 ;
        RECT 2044.385 15.385 2053.755 15.555 ;
        RECT 2044.385 15.215 2044.555 15.385 ;
        RECT 2042.545 15.045 2044.555 15.215 ;
        RECT 2042.545 14.365 2042.715 15.045 ;
      LAYER mcon ;
        RECT 2105.105 1685.805 2105.275 1685.975 ;
        RECT 2053.585 15.385 2053.755 15.555 ;
      LAYER met1 ;
        RECT 2088.010 1685.960 2088.330 1686.020 ;
        RECT 2105.045 1685.960 2105.335 1686.005 ;
        RECT 2088.010 1685.820 2105.335 1685.960 ;
        RECT 2088.010 1685.760 2088.330 1685.820 ;
        RECT 2105.045 1685.775 2105.335 1685.820 ;
        RECT 2105.045 1684.260 2105.335 1684.305 ;
        RECT 2138.610 1684.260 2138.930 1684.320 ;
        RECT 2105.045 1684.120 2138.930 1684.260 ;
        RECT 2105.045 1684.075 2105.335 1684.120 ;
        RECT 2138.610 1684.060 2138.930 1684.120 ;
        RECT 2083.870 16.560 2084.190 16.620 ;
        RECT 2087.090 16.560 2087.410 16.620 ;
        RECT 2083.870 16.420 2087.410 16.560 ;
        RECT 2083.870 16.360 2084.190 16.420 ;
        RECT 2087.090 16.360 2087.410 16.420 ;
        RECT 2053.525 15.540 2053.815 15.585 ;
        RECT 2083.870 15.540 2084.190 15.600 ;
        RECT 2053.525 15.400 2084.190 15.540 ;
        RECT 2053.525 15.355 2053.815 15.400 ;
        RECT 2083.870 15.340 2084.190 15.400 ;
        RECT 1923.330 14.520 1923.650 14.580 ;
        RECT 2042.485 14.520 2042.775 14.565 ;
        RECT 1923.330 14.380 2042.775 14.520 ;
        RECT 1923.330 14.320 1923.650 14.380 ;
        RECT 2042.485 14.335 2042.775 14.380 ;
      LAYER via ;
        RECT 2088.040 1685.760 2088.300 1686.020 ;
        RECT 2138.640 1684.060 2138.900 1684.320 ;
        RECT 2083.900 16.360 2084.160 16.620 ;
        RECT 2087.120 16.360 2087.380 16.620 ;
        RECT 2083.900 15.340 2084.160 15.600 ;
        RECT 1923.360 14.320 1923.620 14.580 ;
      LAYER met2 ;
        RECT 2138.560 1700.000 2138.840 1704.000 ;
        RECT 2088.040 1685.730 2088.300 1686.050 ;
        RECT 2088.100 1671.170 2088.240 1685.730 ;
        RECT 2138.700 1684.350 2138.840 1700.000 ;
        RECT 2138.640 1684.030 2138.900 1684.350 ;
        RECT 2087.180 1671.030 2088.240 1671.170 ;
        RECT 2087.180 16.650 2087.320 1671.030 ;
        RECT 2083.900 16.330 2084.160 16.650 ;
        RECT 2087.120 16.330 2087.380 16.650 ;
        RECT 2083.960 15.630 2084.100 16.330 ;
        RECT 2083.900 15.310 2084.160 15.630 ;
        RECT 1923.360 14.290 1923.620 14.610 ;
        RECT 1923.420 2.400 1923.560 14.290 ;
        RECT 1923.210 -4.800 1923.770 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1945.410 1687.660 1945.730 1687.720 ;
        RECT 1945.410 1687.520 2114.920 1687.660 ;
        RECT 1945.410 1687.460 1945.730 1687.520 ;
        RECT 2114.780 1686.980 2114.920 1687.520 ;
        RECT 2147.810 1686.980 2148.130 1687.040 ;
        RECT 2114.780 1686.840 2148.130 1686.980 ;
        RECT 2147.810 1686.780 2148.130 1686.840 ;
        RECT 1941.270 18.260 1941.590 18.320 ;
        RECT 1945.410 18.260 1945.730 18.320 ;
        RECT 1941.270 18.120 1945.730 18.260 ;
        RECT 1941.270 18.060 1941.590 18.120 ;
        RECT 1945.410 18.060 1945.730 18.120 ;
      LAYER via ;
        RECT 1945.440 1687.460 1945.700 1687.720 ;
        RECT 2147.840 1686.780 2148.100 1687.040 ;
        RECT 1941.300 18.060 1941.560 18.320 ;
        RECT 1945.440 18.060 1945.700 18.320 ;
      LAYER met2 ;
        RECT 2147.760 1700.000 2148.040 1704.000 ;
        RECT 1945.440 1687.430 1945.700 1687.750 ;
        RECT 1945.500 18.350 1945.640 1687.430 ;
        RECT 2147.900 1687.070 2148.040 1700.000 ;
        RECT 2147.840 1686.750 2148.100 1687.070 ;
        RECT 1941.300 18.030 1941.560 18.350 ;
        RECT 1945.440 18.030 1945.700 18.350 ;
        RECT 1941.360 2.400 1941.500 18.030 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2118.445 18.105 2118.615 20.655 ;
      LAYER mcon ;
        RECT 2118.445 20.485 2118.615 20.655 ;
      LAYER met1 ;
        RECT 2152.870 1678.140 2153.190 1678.200 ;
        RECT 2155.630 1678.140 2155.950 1678.200 ;
        RECT 2152.870 1678.000 2155.950 1678.140 ;
        RECT 2152.870 1677.940 2153.190 1678.000 ;
        RECT 2155.630 1677.940 2155.950 1678.000 ;
        RECT 2149.280 20.840 2153.100 20.980 ;
        RECT 2118.385 20.640 2118.675 20.685 ;
        RECT 2149.280 20.640 2149.420 20.840 ;
        RECT 2152.960 20.700 2153.100 20.840 ;
        RECT 2118.385 20.500 2149.420 20.640 ;
        RECT 2118.385 20.455 2118.675 20.500 ;
        RECT 2152.870 20.440 2153.190 20.700 ;
        RECT 1959.210 18.260 1959.530 18.320 ;
        RECT 2041.550 18.260 2041.870 18.320 ;
        RECT 1959.210 18.120 2041.870 18.260 ;
        RECT 1959.210 18.060 1959.530 18.120 ;
        RECT 2041.550 18.060 2041.870 18.120 ;
        RECT 2042.930 18.260 2043.250 18.320 ;
        RECT 2118.385 18.260 2118.675 18.305 ;
        RECT 2042.930 18.120 2118.675 18.260 ;
        RECT 2042.930 18.060 2043.250 18.120 ;
        RECT 2118.385 18.075 2118.675 18.120 ;
      LAYER via ;
        RECT 2152.900 1677.940 2153.160 1678.200 ;
        RECT 2155.660 1677.940 2155.920 1678.200 ;
        RECT 2152.900 20.440 2153.160 20.700 ;
        RECT 1959.240 18.060 1959.500 18.320 ;
        RECT 2041.580 18.060 2041.840 18.320 ;
        RECT 2042.960 18.060 2043.220 18.320 ;
      LAYER met2 ;
        RECT 2156.960 1700.410 2157.240 1704.000 ;
        RECT 2155.720 1700.270 2157.240 1700.410 ;
        RECT 2155.720 1678.230 2155.860 1700.270 ;
        RECT 2156.960 1700.000 2157.240 1700.270 ;
        RECT 2152.900 1677.910 2153.160 1678.230 ;
        RECT 2155.660 1677.910 2155.920 1678.230 ;
        RECT 2152.960 20.730 2153.100 1677.910 ;
        RECT 2152.900 20.410 2153.160 20.730 ;
        RECT 1959.240 18.030 1959.500 18.350 ;
        RECT 2041.580 18.205 2041.840 18.350 ;
        RECT 2042.960 18.205 2043.220 18.350 ;
        RECT 1959.300 2.400 1959.440 18.030 ;
        RECT 2041.570 17.835 2041.850 18.205 ;
        RECT 2042.950 17.835 2043.230 18.205 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
      LAYER via2 ;
        RECT 2041.570 17.880 2041.850 18.160 ;
        RECT 2042.950 17.880 2043.230 18.160 ;
      LAYER met3 ;
        RECT 2041.545 18.170 2041.875 18.185 ;
        RECT 2042.925 18.170 2043.255 18.185 ;
        RECT 2041.545 17.870 2043.255 18.170 ;
        RECT 2041.545 17.855 2041.875 17.870 ;
        RECT 2042.925 17.855 2043.255 17.870 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2152.485 1685.125 2152.655 1685.975 ;
      LAYER mcon ;
        RECT 2152.485 1685.805 2152.655 1685.975 ;
      LAYER met1 ;
        RECT 2152.425 1685.960 2152.715 1686.005 ;
        RECT 2166.210 1685.960 2166.530 1686.020 ;
        RECT 2152.425 1685.820 2166.530 1685.960 ;
        RECT 2152.425 1685.775 2152.715 1685.820 ;
        RECT 2166.210 1685.760 2166.530 1685.820 ;
        RECT 2100.890 1685.280 2101.210 1685.340 ;
        RECT 2152.425 1685.280 2152.715 1685.325 ;
        RECT 2100.890 1685.140 2152.715 1685.280 ;
        RECT 2100.890 1685.080 2101.210 1685.140 ;
        RECT 2152.425 1685.095 2152.715 1685.140 ;
        RECT 1977.150 14.180 1977.470 14.240 ;
        RECT 2100.890 14.180 2101.210 14.240 ;
        RECT 1977.150 14.040 2101.210 14.180 ;
        RECT 1977.150 13.980 1977.470 14.040 ;
        RECT 2100.890 13.980 2101.210 14.040 ;
      LAYER via ;
        RECT 2166.240 1685.760 2166.500 1686.020 ;
        RECT 2100.920 1685.080 2101.180 1685.340 ;
        RECT 1977.180 13.980 1977.440 14.240 ;
        RECT 2100.920 13.980 2101.180 14.240 ;
      LAYER met2 ;
        RECT 2166.160 1700.000 2166.440 1704.000 ;
        RECT 2166.300 1686.050 2166.440 1700.000 ;
        RECT 2166.240 1685.730 2166.500 1686.050 ;
        RECT 2100.920 1685.050 2101.180 1685.370 ;
        RECT 2100.980 14.270 2101.120 1685.050 ;
        RECT 1977.180 13.950 1977.440 14.270 ;
        RECT 2100.920 13.950 2101.180 14.270 ;
        RECT 1977.240 2.400 1977.380 13.950 ;
        RECT 1977.030 -4.800 1977.590 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1995.090 18.940 1995.410 19.000 ;
        RECT 2174.030 18.940 2174.350 19.000 ;
        RECT 1995.090 18.800 2174.350 18.940 ;
        RECT 1995.090 18.740 1995.410 18.800 ;
        RECT 2174.030 18.740 2174.350 18.800 ;
      LAYER via ;
        RECT 1995.120 18.740 1995.380 19.000 ;
        RECT 2174.060 18.740 2174.320 19.000 ;
      LAYER met2 ;
        RECT 2175.360 1700.410 2175.640 1704.000 ;
        RECT 2174.120 1700.270 2175.640 1700.410 ;
        RECT 2174.120 19.030 2174.260 1700.270 ;
        RECT 2175.360 1700.000 2175.640 1700.270 ;
        RECT 1995.120 18.710 1995.380 19.030 ;
        RECT 2174.060 18.710 2174.320 19.030 ;
        RECT 1995.180 2.400 1995.320 18.710 ;
        RECT 1994.970 -4.800 1995.530 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2163.525 1687.335 2163.695 1689.035 ;
        RECT 2162.605 1687.165 2163.695 1687.335 ;
        RECT 2155.705 1684.785 2155.875 1686.995 ;
        RECT 2162.605 1686.825 2162.775 1687.165 ;
        RECT 2017.705 19.125 2017.875 20.655 ;
        RECT 2046.225 19.805 2046.395 20.655 ;
      LAYER mcon ;
        RECT 2163.525 1688.865 2163.695 1689.035 ;
        RECT 2155.705 1686.825 2155.875 1686.995 ;
        RECT 2017.705 20.485 2017.875 20.655 ;
        RECT 2046.225 20.485 2046.395 20.655 ;
      LAYER met1 ;
        RECT 2163.465 1689.020 2163.755 1689.065 ;
        RECT 2184.610 1689.020 2184.930 1689.080 ;
        RECT 2163.465 1688.880 2184.930 1689.020 ;
        RECT 2163.465 1688.835 2163.755 1688.880 ;
        RECT 2184.610 1688.820 2184.930 1688.880 ;
        RECT 2155.645 1686.980 2155.935 1687.025 ;
        RECT 2162.545 1686.980 2162.835 1687.025 ;
        RECT 2155.645 1686.840 2162.835 1686.980 ;
        RECT 2155.645 1686.795 2155.935 1686.840 ;
        RECT 2162.545 1686.795 2162.835 1686.840 ;
        RECT 2122.050 1684.940 2122.370 1685.000 ;
        RECT 2155.645 1684.940 2155.935 1684.985 ;
        RECT 2122.050 1684.800 2155.935 1684.940 ;
        RECT 2122.050 1684.740 2122.370 1684.800 ;
        RECT 2155.645 1684.755 2155.935 1684.800 ;
        RECT 2017.645 20.640 2017.935 20.685 ;
        RECT 2046.165 20.640 2046.455 20.685 ;
        RECT 2017.645 20.500 2046.455 20.640 ;
        RECT 2017.645 20.455 2017.935 20.500 ;
        RECT 2046.165 20.455 2046.455 20.500 ;
        RECT 2046.165 19.960 2046.455 20.005 ;
        RECT 2122.050 19.960 2122.370 20.020 ;
        RECT 2046.165 19.820 2122.370 19.960 ;
        RECT 2046.165 19.775 2046.455 19.820 ;
        RECT 2122.050 19.760 2122.370 19.820 ;
        RECT 2012.570 19.280 2012.890 19.340 ;
        RECT 2017.645 19.280 2017.935 19.325 ;
        RECT 2012.570 19.140 2017.935 19.280 ;
        RECT 2012.570 19.080 2012.890 19.140 ;
        RECT 2017.645 19.095 2017.935 19.140 ;
      LAYER via ;
        RECT 2184.640 1688.820 2184.900 1689.080 ;
        RECT 2122.080 1684.740 2122.340 1685.000 ;
        RECT 2122.080 19.760 2122.340 20.020 ;
        RECT 2012.600 19.080 2012.860 19.340 ;
      LAYER met2 ;
        RECT 2184.560 1700.000 2184.840 1704.000 ;
        RECT 2184.700 1689.110 2184.840 1700.000 ;
        RECT 2184.640 1688.790 2184.900 1689.110 ;
        RECT 2122.080 1684.710 2122.340 1685.030 ;
        RECT 2122.140 20.050 2122.280 1684.710 ;
        RECT 2122.080 19.730 2122.340 20.050 ;
        RECT 2012.600 19.050 2012.860 19.370 ;
        RECT 2012.660 2.400 2012.800 19.050 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2163.065 1683.765 2163.235 1684.615 ;
        RECT 2105.565 14.705 2105.735 16.235 ;
      LAYER mcon ;
        RECT 2163.065 1684.445 2163.235 1684.615 ;
        RECT 2105.565 16.065 2105.735 16.235 ;
      LAYER met1 ;
        RECT 2187.370 1689.020 2187.690 1689.080 ;
        RECT 2193.810 1689.020 2194.130 1689.080 ;
        RECT 2187.370 1688.880 2194.130 1689.020 ;
        RECT 2187.370 1688.820 2187.690 1688.880 ;
        RECT 2193.810 1688.820 2194.130 1688.880 ;
        RECT 2135.390 1684.600 2135.710 1684.660 ;
        RECT 2163.005 1684.600 2163.295 1684.645 ;
        RECT 2135.390 1684.460 2163.295 1684.600 ;
        RECT 2135.390 1684.400 2135.710 1684.460 ;
        RECT 2163.005 1684.415 2163.295 1684.460 ;
        RECT 2163.005 1683.920 2163.295 1683.965 ;
        RECT 2187.370 1683.920 2187.690 1683.980 ;
        RECT 2163.005 1683.780 2187.690 1683.920 ;
        RECT 2163.005 1683.735 2163.295 1683.780 ;
        RECT 2187.370 1683.720 2187.690 1683.780 ;
        RECT 2030.510 16.560 2030.830 16.620 ;
        RECT 2030.510 16.420 2066.620 16.560 ;
        RECT 2030.510 16.360 2030.830 16.420 ;
        RECT 2066.480 16.220 2066.620 16.420 ;
        RECT 2105.505 16.220 2105.795 16.265 ;
        RECT 2066.480 16.080 2105.795 16.220 ;
        RECT 2105.505 16.035 2105.795 16.080 ;
        RECT 2105.505 14.860 2105.795 14.905 ;
        RECT 2135.390 14.860 2135.710 14.920 ;
        RECT 2105.505 14.720 2135.710 14.860 ;
        RECT 2105.505 14.675 2105.795 14.720 ;
        RECT 2135.390 14.660 2135.710 14.720 ;
      LAYER via ;
        RECT 2187.400 1688.820 2187.660 1689.080 ;
        RECT 2193.840 1688.820 2194.100 1689.080 ;
        RECT 2135.420 1684.400 2135.680 1684.660 ;
        RECT 2187.400 1683.720 2187.660 1683.980 ;
        RECT 2030.540 16.360 2030.800 16.620 ;
        RECT 2135.420 14.660 2135.680 14.920 ;
      LAYER met2 ;
        RECT 2193.760 1700.000 2194.040 1704.000 ;
        RECT 2193.900 1689.110 2194.040 1700.000 ;
        RECT 2187.400 1688.790 2187.660 1689.110 ;
        RECT 2193.840 1688.790 2194.100 1689.110 ;
        RECT 2135.420 1684.370 2135.680 1684.690 ;
        RECT 2030.540 16.330 2030.800 16.650 ;
        RECT 2030.600 2.400 2030.740 16.330 ;
        RECT 2135.480 14.950 2135.620 1684.370 ;
        RECT 2187.460 1684.010 2187.600 1688.790 ;
        RECT 2187.400 1683.690 2187.660 1684.010 ;
        RECT 2135.420 14.630 2135.680 14.950 ;
        RECT 2030.390 -4.800 2030.950 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2109.705 15.725 2109.875 16.915 ;
      LAYER mcon ;
        RECT 2109.705 16.745 2109.875 16.915 ;
      LAYER met1 ;
        RECT 2156.090 1684.940 2156.410 1685.000 ;
        RECT 2156.090 1684.800 2163.680 1684.940 ;
        RECT 2156.090 1684.740 2156.410 1684.800 ;
        RECT 2163.540 1684.600 2163.680 1684.800 ;
        RECT 2203.010 1684.600 2203.330 1684.660 ;
        RECT 2163.540 1684.460 2203.330 1684.600 ;
        RECT 2203.010 1684.400 2203.330 1684.460 ;
        RECT 2048.450 16.900 2048.770 16.960 ;
        RECT 2109.645 16.900 2109.935 16.945 ;
        RECT 2048.450 16.760 2109.935 16.900 ;
        RECT 2048.450 16.700 2048.770 16.760 ;
        RECT 2109.645 16.715 2109.935 16.760 ;
        RECT 2109.645 15.880 2109.935 15.925 ;
        RECT 2156.090 15.880 2156.410 15.940 ;
        RECT 2109.645 15.740 2156.410 15.880 ;
        RECT 2109.645 15.695 2109.935 15.740 ;
        RECT 2156.090 15.680 2156.410 15.740 ;
      LAYER via ;
        RECT 2156.120 1684.740 2156.380 1685.000 ;
        RECT 2203.040 1684.400 2203.300 1684.660 ;
        RECT 2048.480 16.700 2048.740 16.960 ;
        RECT 2156.120 15.680 2156.380 15.940 ;
      LAYER met2 ;
        RECT 2202.960 1700.000 2203.240 1704.000 ;
        RECT 2156.120 1684.710 2156.380 1685.030 ;
        RECT 2048.480 16.670 2048.740 16.990 ;
        RECT 2048.540 2.400 2048.680 16.670 ;
        RECT 2156.180 15.970 2156.320 1684.710 ;
        RECT 2203.100 1684.690 2203.240 1700.000 ;
        RECT 2203.040 1684.370 2203.300 1684.690 ;
        RECT 2156.120 15.650 2156.380 15.970 ;
        RECT 2048.330 -4.800 2048.890 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1539.230 1678.140 1539.550 1678.200 ;
        RECT 1540.150 1678.140 1540.470 1678.200 ;
        RECT 1539.230 1678.000 1540.470 1678.140 ;
        RECT 1539.230 1677.940 1539.550 1678.000 ;
        RECT 1540.150 1677.940 1540.470 1678.000 ;
        RECT 765.510 67.900 765.830 67.960 ;
        RECT 1539.230 67.900 1539.550 67.960 ;
        RECT 765.510 67.760 1539.550 67.900 ;
        RECT 765.510 67.700 765.830 67.760 ;
        RECT 1539.230 67.700 1539.550 67.760 ;
      LAYER via ;
        RECT 1539.260 1677.940 1539.520 1678.200 ;
        RECT 1540.180 1677.940 1540.440 1678.200 ;
        RECT 765.540 67.700 765.800 67.960 ;
        RECT 1539.260 67.700 1539.520 67.960 ;
      LAYER met2 ;
        RECT 1541.480 1700.410 1541.760 1704.000 ;
        RECT 1540.240 1700.270 1541.760 1700.410 ;
        RECT 1540.240 1678.230 1540.380 1700.270 ;
        RECT 1541.480 1700.000 1541.760 1700.270 ;
        RECT 1539.260 1677.910 1539.520 1678.230 ;
        RECT 1540.180 1677.910 1540.440 1678.230 ;
        RECT 1539.320 67.990 1539.460 1677.910 ;
        RECT 765.540 67.670 765.800 67.990 ;
        RECT 1539.260 67.670 1539.520 67.990 ;
        RECT 765.600 16.730 765.740 67.670 ;
        RECT 763.760 16.590 765.740 16.730 ;
        RECT 763.760 2.400 763.900 16.590 ;
        RECT 763.550 -4.800 764.110 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2114.765 15.045 2114.935 16.575 ;
      LAYER mcon ;
        RECT 2114.765 16.405 2114.935 16.575 ;
      LAYER met1 ;
        RECT 2176.790 1684.260 2177.110 1684.320 ;
        RECT 2212.210 1684.260 2212.530 1684.320 ;
        RECT 2176.790 1684.120 2212.530 1684.260 ;
        RECT 2176.790 1684.060 2177.110 1684.120 ;
        RECT 2212.210 1684.060 2212.530 1684.120 ;
        RECT 2114.705 16.560 2114.995 16.605 ;
        RECT 2114.705 16.420 2158.160 16.560 ;
        RECT 2114.705 16.375 2114.995 16.420 ;
        RECT 2158.020 15.880 2158.160 16.420 ;
        RECT 2176.790 15.880 2177.110 15.940 ;
        RECT 2158.020 15.740 2177.110 15.880 ;
        RECT 2176.790 15.680 2177.110 15.740 ;
        RECT 2066.850 15.200 2067.170 15.260 ;
        RECT 2114.705 15.200 2114.995 15.245 ;
        RECT 2066.850 15.060 2114.995 15.200 ;
        RECT 2066.850 15.000 2067.170 15.060 ;
        RECT 2114.705 15.015 2114.995 15.060 ;
      LAYER via ;
        RECT 2176.820 1684.060 2177.080 1684.320 ;
        RECT 2212.240 1684.060 2212.500 1684.320 ;
        RECT 2176.820 15.680 2177.080 15.940 ;
        RECT 2066.880 15.000 2067.140 15.260 ;
      LAYER met2 ;
        RECT 2212.160 1700.000 2212.440 1704.000 ;
        RECT 2212.300 1684.350 2212.440 1700.000 ;
        RECT 2176.820 1684.030 2177.080 1684.350 ;
        RECT 2212.240 1684.030 2212.500 1684.350 ;
        RECT 2176.880 15.970 2177.020 1684.030 ;
        RECT 2176.820 15.650 2177.080 15.970 ;
        RECT 2066.880 14.970 2067.140 15.290 ;
        RECT 2066.940 8.570 2067.080 14.970 ;
        RECT 2066.480 8.430 2067.080 8.570 ;
        RECT 2066.480 2.400 2066.620 8.430 ;
        RECT 2066.270 -4.800 2066.830 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2190.590 1683.920 2190.910 1683.980 ;
        RECT 2221.410 1683.920 2221.730 1683.980 ;
        RECT 2190.590 1683.780 2221.730 1683.920 ;
        RECT 2190.590 1683.720 2190.910 1683.780 ;
        RECT 2221.410 1683.720 2221.730 1683.780 ;
        RECT 2084.330 15.540 2084.650 15.600 ;
        RECT 2190.590 15.540 2190.910 15.600 ;
        RECT 2084.330 15.400 2190.910 15.540 ;
        RECT 2084.330 15.340 2084.650 15.400 ;
        RECT 2190.590 15.340 2190.910 15.400 ;
      LAYER via ;
        RECT 2190.620 1683.720 2190.880 1683.980 ;
        RECT 2221.440 1683.720 2221.700 1683.980 ;
        RECT 2084.360 15.340 2084.620 15.600 ;
        RECT 2190.620 15.340 2190.880 15.600 ;
      LAYER met2 ;
        RECT 2221.360 1700.000 2221.640 1704.000 ;
        RECT 2221.500 1684.010 2221.640 1700.000 ;
        RECT 2190.620 1683.690 2190.880 1684.010 ;
        RECT 2221.440 1683.690 2221.700 1684.010 ;
        RECT 2190.680 15.630 2190.820 1683.690 ;
        RECT 2084.360 15.310 2084.620 15.630 ;
        RECT 2190.620 15.310 2190.880 15.630 ;
        RECT 2084.420 2.400 2084.560 15.310 ;
        RECT 2084.210 -4.800 2084.770 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2104.110 1688.340 2104.430 1688.400 ;
        RECT 2230.610 1688.340 2230.930 1688.400 ;
        RECT 2104.110 1688.200 2230.930 1688.340 ;
        RECT 2104.110 1688.140 2104.430 1688.200 ;
        RECT 2230.610 1688.140 2230.930 1688.200 ;
        RECT 2101.810 20.640 2102.130 20.700 ;
        RECT 2104.110 20.640 2104.430 20.700 ;
        RECT 2101.810 20.500 2104.430 20.640 ;
        RECT 2101.810 20.440 2102.130 20.500 ;
        RECT 2104.110 20.440 2104.430 20.500 ;
      LAYER via ;
        RECT 2104.140 1688.140 2104.400 1688.400 ;
        RECT 2230.640 1688.140 2230.900 1688.400 ;
        RECT 2101.840 20.440 2102.100 20.700 ;
        RECT 2104.140 20.440 2104.400 20.700 ;
      LAYER met2 ;
        RECT 2230.560 1700.000 2230.840 1704.000 ;
        RECT 2230.700 1688.430 2230.840 1700.000 ;
        RECT 2104.140 1688.110 2104.400 1688.430 ;
        RECT 2230.640 1688.110 2230.900 1688.430 ;
        RECT 2104.200 20.730 2104.340 1688.110 ;
        RECT 2101.840 20.410 2102.100 20.730 ;
        RECT 2104.140 20.410 2104.400 20.730 ;
        RECT 2101.900 2.400 2102.040 20.410 ;
        RECT 2101.690 -4.800 2102.250 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2124.810 1686.300 2125.130 1686.360 ;
        RECT 2239.810 1686.300 2240.130 1686.360 ;
        RECT 2124.810 1686.160 2240.130 1686.300 ;
        RECT 2124.810 1686.100 2125.130 1686.160 ;
        RECT 2239.810 1686.100 2240.130 1686.160 ;
        RECT 2119.750 16.220 2120.070 16.280 ;
        RECT 2124.810 16.220 2125.130 16.280 ;
        RECT 2119.750 16.080 2125.130 16.220 ;
        RECT 2119.750 16.020 2120.070 16.080 ;
        RECT 2124.810 16.020 2125.130 16.080 ;
      LAYER via ;
        RECT 2124.840 1686.100 2125.100 1686.360 ;
        RECT 2239.840 1686.100 2240.100 1686.360 ;
        RECT 2119.780 16.020 2120.040 16.280 ;
        RECT 2124.840 16.020 2125.100 16.280 ;
      LAYER met2 ;
        RECT 2239.760 1700.000 2240.040 1704.000 ;
        RECT 2239.900 1686.390 2240.040 1700.000 ;
        RECT 2124.840 1686.070 2125.100 1686.390 ;
        RECT 2239.840 1686.070 2240.100 1686.390 ;
        RECT 2124.900 16.310 2125.040 1686.070 ;
        RECT 2119.780 15.990 2120.040 16.310 ;
        RECT 2124.840 15.990 2125.100 16.310 ;
        RECT 2119.840 2.400 2119.980 15.990 ;
        RECT 2119.630 -4.800 2120.190 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2211.290 1689.700 2211.610 1689.760 ;
        RECT 2249.010 1689.700 2249.330 1689.760 ;
        RECT 2211.290 1689.560 2249.330 1689.700 ;
        RECT 2211.290 1689.500 2211.610 1689.560 ;
        RECT 2249.010 1689.500 2249.330 1689.560 ;
        RECT 2137.690 19.960 2138.010 20.020 ;
        RECT 2137.690 19.820 2163.220 19.960 ;
        RECT 2137.690 19.760 2138.010 19.820 ;
        RECT 2163.080 19.620 2163.220 19.820 ;
        RECT 2211.290 19.620 2211.610 19.680 ;
        RECT 2163.080 19.480 2211.610 19.620 ;
        RECT 2211.290 19.420 2211.610 19.480 ;
      LAYER via ;
        RECT 2211.320 1689.500 2211.580 1689.760 ;
        RECT 2249.040 1689.500 2249.300 1689.760 ;
        RECT 2137.720 19.760 2137.980 20.020 ;
        RECT 2211.320 19.420 2211.580 19.680 ;
      LAYER met2 ;
        RECT 2248.960 1700.000 2249.240 1704.000 ;
        RECT 2249.100 1689.790 2249.240 1700.000 ;
        RECT 2211.320 1689.470 2211.580 1689.790 ;
        RECT 2249.040 1689.470 2249.300 1689.790 ;
        RECT 2137.720 19.730 2137.980 20.050 ;
        RECT 2137.780 2.400 2137.920 19.730 ;
        RECT 2211.380 19.710 2211.520 1689.470 ;
        RECT 2211.320 19.390 2211.580 19.710 ;
        RECT 2137.570 -4.800 2138.130 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2258.210 1685.620 2258.530 1685.680 ;
        RECT 2164.000 1685.480 2258.530 1685.620 ;
        RECT 2159.310 1685.280 2159.630 1685.340 ;
        RECT 2164.000 1685.280 2164.140 1685.480 ;
        RECT 2258.210 1685.420 2258.530 1685.480 ;
        RECT 2159.310 1685.140 2164.140 1685.280 ;
        RECT 2159.310 1685.080 2159.630 1685.140 ;
        RECT 2155.630 20.640 2155.950 20.700 ;
        RECT 2159.310 20.640 2159.630 20.700 ;
        RECT 2155.630 20.500 2159.630 20.640 ;
        RECT 2155.630 20.440 2155.950 20.500 ;
        RECT 2159.310 20.440 2159.630 20.500 ;
      LAYER via ;
        RECT 2159.340 1685.080 2159.600 1685.340 ;
        RECT 2258.240 1685.420 2258.500 1685.680 ;
        RECT 2155.660 20.440 2155.920 20.700 ;
        RECT 2159.340 20.440 2159.600 20.700 ;
      LAYER met2 ;
        RECT 2258.160 1700.000 2258.440 1704.000 ;
        RECT 2258.300 1685.710 2258.440 1700.000 ;
        RECT 2258.240 1685.390 2258.500 1685.710 ;
        RECT 2159.340 1685.050 2159.600 1685.370 ;
        RECT 2159.400 20.730 2159.540 1685.050 ;
        RECT 2155.660 20.410 2155.920 20.730 ;
        RECT 2159.340 20.410 2159.600 20.730 ;
        RECT 2155.720 2.400 2155.860 20.410 ;
        RECT 2155.510 -4.800 2156.070 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2267.410 1684.600 2267.730 1684.660 ;
        RECT 2235.760 1684.460 2267.730 1684.600 ;
        RECT 2231.990 1683.920 2232.310 1683.980 ;
        RECT 2235.760 1683.920 2235.900 1684.460 ;
        RECT 2267.410 1684.400 2267.730 1684.460 ;
        RECT 2231.990 1683.780 2235.900 1683.920 ;
        RECT 2231.990 1683.720 2232.310 1683.780 ;
        RECT 2172.650 18.600 2172.970 18.660 ;
        RECT 2231.990 18.600 2232.310 18.660 ;
        RECT 2172.650 18.460 2232.310 18.600 ;
        RECT 2172.650 18.400 2172.970 18.460 ;
        RECT 2231.990 18.400 2232.310 18.460 ;
      LAYER via ;
        RECT 2232.020 1683.720 2232.280 1683.980 ;
        RECT 2267.440 1684.400 2267.700 1684.660 ;
        RECT 2172.680 18.400 2172.940 18.660 ;
        RECT 2232.020 18.400 2232.280 18.660 ;
      LAYER met2 ;
        RECT 2267.360 1700.000 2267.640 1704.000 ;
        RECT 2267.500 1684.690 2267.640 1700.000 ;
        RECT 2267.440 1684.370 2267.700 1684.690 ;
        RECT 2232.020 1683.690 2232.280 1684.010 ;
        RECT 2232.080 18.690 2232.220 1683.690 ;
        RECT 2172.680 18.370 2172.940 18.690 ;
        RECT 2232.020 18.370 2232.280 18.690 ;
        RECT 2172.740 9.250 2172.880 18.370 ;
        RECT 2172.740 9.110 2173.340 9.250 ;
        RECT 2173.200 2.400 2173.340 9.110 ;
        RECT 2172.990 -4.800 2173.550 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2238.890 1683.920 2239.210 1683.980 ;
        RECT 2276.610 1683.920 2276.930 1683.980 ;
        RECT 2238.890 1683.780 2276.930 1683.920 ;
        RECT 2238.890 1683.720 2239.210 1683.780 ;
        RECT 2276.610 1683.720 2276.930 1683.780 ;
        RECT 2191.050 18.940 2191.370 19.000 ;
        RECT 2238.890 18.940 2239.210 19.000 ;
        RECT 2191.050 18.800 2239.210 18.940 ;
        RECT 2191.050 18.740 2191.370 18.800 ;
        RECT 2238.890 18.740 2239.210 18.800 ;
      LAYER via ;
        RECT 2238.920 1683.720 2239.180 1683.980 ;
        RECT 2276.640 1683.720 2276.900 1683.980 ;
        RECT 2191.080 18.740 2191.340 19.000 ;
        RECT 2238.920 18.740 2239.180 19.000 ;
      LAYER met2 ;
        RECT 2276.560 1700.000 2276.840 1704.000 ;
        RECT 2276.700 1684.010 2276.840 1700.000 ;
        RECT 2238.920 1683.690 2239.180 1684.010 ;
        RECT 2276.640 1683.690 2276.900 1684.010 ;
        RECT 2238.980 19.030 2239.120 1683.690 ;
        RECT 2191.080 18.710 2191.340 19.030 ;
        RECT 2238.920 18.710 2239.180 19.030 ;
        RECT 2191.140 2.400 2191.280 18.710 ;
        RECT 2190.930 -4.800 2191.490 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2246.250 1689.360 2246.570 1689.420 ;
        RECT 2285.810 1689.360 2286.130 1689.420 ;
        RECT 2246.250 1689.220 2286.130 1689.360 ;
        RECT 2246.250 1689.160 2246.570 1689.220 ;
        RECT 2285.810 1689.160 2286.130 1689.220 ;
        RECT 2245.790 16.900 2246.110 16.960 ;
        RECT 2238.520 16.760 2246.110 16.900 ;
        RECT 2208.990 16.560 2209.310 16.620 ;
        RECT 2238.520 16.560 2238.660 16.760 ;
        RECT 2245.790 16.700 2246.110 16.760 ;
        RECT 2208.990 16.420 2238.660 16.560 ;
        RECT 2208.990 16.360 2209.310 16.420 ;
      LAYER via ;
        RECT 2246.280 1689.160 2246.540 1689.420 ;
        RECT 2285.840 1689.160 2286.100 1689.420 ;
        RECT 2209.020 16.360 2209.280 16.620 ;
        RECT 2245.820 16.700 2246.080 16.960 ;
      LAYER met2 ;
        RECT 2285.760 1700.000 2286.040 1704.000 ;
        RECT 2285.900 1689.450 2286.040 1700.000 ;
        RECT 2246.280 1689.130 2246.540 1689.450 ;
        RECT 2285.840 1689.130 2286.100 1689.450 ;
        RECT 2246.340 1672.530 2246.480 1689.130 ;
        RECT 2245.880 1672.390 2246.480 1672.530 ;
        RECT 2245.880 16.990 2246.020 1672.390 ;
        RECT 2245.820 16.670 2246.080 16.990 ;
        RECT 2209.020 16.330 2209.280 16.650 ;
        RECT 2209.080 2.400 2209.220 16.330 ;
        RECT 2208.870 -4.800 2209.430 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2259.590 1690.040 2259.910 1690.100 ;
        RECT 2295.010 1690.040 2295.330 1690.100 ;
        RECT 2259.590 1689.900 2295.330 1690.040 ;
        RECT 2259.590 1689.840 2259.910 1689.900 ;
        RECT 2295.010 1689.840 2295.330 1689.900 ;
        RECT 2226.930 20.300 2227.250 20.360 ;
        RECT 2259.590 20.300 2259.910 20.360 ;
        RECT 2226.930 20.160 2259.910 20.300 ;
        RECT 2226.930 20.100 2227.250 20.160 ;
        RECT 2259.590 20.100 2259.910 20.160 ;
      LAYER via ;
        RECT 2259.620 1689.840 2259.880 1690.100 ;
        RECT 2295.040 1689.840 2295.300 1690.100 ;
        RECT 2226.960 20.100 2227.220 20.360 ;
        RECT 2259.620 20.100 2259.880 20.360 ;
      LAYER met2 ;
        RECT 2294.960 1700.000 2295.240 1704.000 ;
        RECT 2295.100 1690.130 2295.240 1700.000 ;
        RECT 2259.620 1689.810 2259.880 1690.130 ;
        RECT 2295.040 1689.810 2295.300 1690.130 ;
        RECT 2259.680 20.390 2259.820 1689.810 ;
        RECT 2226.960 20.070 2227.220 20.390 ;
        RECT 2259.620 20.070 2259.880 20.390 ;
        RECT 2227.020 2.400 2227.160 20.070 ;
        RECT 2226.810 -4.800 2227.370 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1546.665 1497.445 1546.835 1545.555 ;
        RECT 1546.665 1400.885 1546.835 1448.655 ;
        RECT 1546.665 1304.325 1546.835 1352.095 ;
        RECT 1546.665 1256.045 1546.835 1303.815 ;
        RECT 1546.665 1110.865 1546.835 1158.975 ;
        RECT 1546.665 917.745 1546.835 1007.335 ;
        RECT 1546.205 448.205 1546.375 524.195 ;
        RECT 1546.665 386.325 1546.835 400.435 ;
        RECT 1546.665 186.405 1546.835 234.515 ;
      LAYER mcon ;
        RECT 1546.665 1545.385 1546.835 1545.555 ;
        RECT 1546.665 1448.485 1546.835 1448.655 ;
        RECT 1546.665 1351.925 1546.835 1352.095 ;
        RECT 1546.665 1303.645 1546.835 1303.815 ;
        RECT 1546.665 1158.805 1546.835 1158.975 ;
        RECT 1546.665 1007.165 1546.835 1007.335 ;
        RECT 1546.205 524.025 1546.375 524.195 ;
        RECT 1546.665 400.265 1546.835 400.435 ;
        RECT 1546.665 234.345 1546.835 234.515 ;
      LAYER met1 ;
        RECT 1547.050 1642.440 1547.370 1642.500 ;
        RECT 1548.430 1642.440 1548.750 1642.500 ;
        RECT 1547.050 1642.300 1548.750 1642.440 ;
        RECT 1547.050 1642.240 1547.370 1642.300 ;
        RECT 1548.430 1642.240 1548.750 1642.300 ;
        RECT 1546.590 1545.540 1546.910 1545.600 ;
        RECT 1546.395 1545.400 1546.910 1545.540 ;
        RECT 1546.590 1545.340 1546.910 1545.400 ;
        RECT 1546.605 1497.600 1546.895 1497.645 ;
        RECT 1547.050 1497.600 1547.370 1497.660 ;
        RECT 1546.605 1497.460 1547.370 1497.600 ;
        RECT 1546.605 1497.415 1546.895 1497.460 ;
        RECT 1547.050 1497.400 1547.370 1497.460 ;
        RECT 1546.590 1449.320 1546.910 1449.380 ;
        RECT 1547.970 1449.320 1548.290 1449.380 ;
        RECT 1546.590 1449.180 1548.290 1449.320 ;
        RECT 1546.590 1449.120 1546.910 1449.180 ;
        RECT 1547.970 1449.120 1548.290 1449.180 ;
        RECT 1546.590 1448.640 1546.910 1448.700 ;
        RECT 1546.395 1448.500 1546.910 1448.640 ;
        RECT 1546.590 1448.440 1546.910 1448.500 ;
        RECT 1546.605 1401.040 1546.895 1401.085 ;
        RECT 1547.050 1401.040 1547.370 1401.100 ;
        RECT 1546.605 1400.900 1547.370 1401.040 ;
        RECT 1546.605 1400.855 1546.895 1400.900 ;
        RECT 1547.050 1400.840 1547.370 1400.900 ;
        RECT 1546.590 1352.760 1546.910 1352.820 ;
        RECT 1547.970 1352.760 1548.290 1352.820 ;
        RECT 1546.590 1352.620 1548.290 1352.760 ;
        RECT 1546.590 1352.560 1546.910 1352.620 ;
        RECT 1547.970 1352.560 1548.290 1352.620 ;
        RECT 1546.590 1352.080 1546.910 1352.140 ;
        RECT 1546.395 1351.940 1546.910 1352.080 ;
        RECT 1546.590 1351.880 1546.910 1351.940 ;
        RECT 1546.605 1304.480 1546.895 1304.525 ;
        RECT 1547.050 1304.480 1547.370 1304.540 ;
        RECT 1546.605 1304.340 1547.370 1304.480 ;
        RECT 1546.605 1304.295 1546.895 1304.340 ;
        RECT 1547.050 1304.280 1547.370 1304.340 ;
        RECT 1546.605 1303.800 1546.895 1303.845 ;
        RECT 1547.050 1303.800 1547.370 1303.860 ;
        RECT 1546.605 1303.660 1547.370 1303.800 ;
        RECT 1546.605 1303.615 1546.895 1303.660 ;
        RECT 1547.050 1303.600 1547.370 1303.660 ;
        RECT 1546.590 1256.200 1546.910 1256.260 ;
        RECT 1546.395 1256.060 1546.910 1256.200 ;
        RECT 1546.590 1256.000 1546.910 1256.060 ;
        RECT 1547.510 1207.580 1547.830 1207.640 ;
        RECT 1547.970 1207.580 1548.290 1207.640 ;
        RECT 1547.510 1207.440 1548.290 1207.580 ;
        RECT 1547.510 1207.380 1547.830 1207.440 ;
        RECT 1547.970 1207.380 1548.290 1207.440 ;
        RECT 1546.590 1172.900 1546.910 1172.960 ;
        RECT 1547.970 1172.900 1548.290 1172.960 ;
        RECT 1546.590 1172.760 1548.290 1172.900 ;
        RECT 1546.590 1172.700 1546.910 1172.760 ;
        RECT 1547.970 1172.700 1548.290 1172.760 ;
        RECT 1546.590 1158.960 1546.910 1159.020 ;
        RECT 1546.395 1158.820 1546.910 1158.960 ;
        RECT 1546.590 1158.760 1546.910 1158.820 ;
        RECT 1546.605 1111.020 1546.895 1111.065 ;
        RECT 1547.510 1111.020 1547.830 1111.080 ;
        RECT 1546.605 1110.880 1547.830 1111.020 ;
        RECT 1546.605 1110.835 1546.895 1110.880 ;
        RECT 1547.510 1110.820 1547.830 1110.880 ;
        RECT 1546.590 1014.800 1546.910 1014.860 ;
        RECT 1547.050 1014.800 1547.370 1014.860 ;
        RECT 1546.590 1014.660 1547.370 1014.800 ;
        RECT 1546.590 1014.600 1546.910 1014.660 ;
        RECT 1547.050 1014.600 1547.370 1014.660 ;
        RECT 1546.605 1007.320 1546.895 1007.365 ;
        RECT 1547.050 1007.320 1547.370 1007.380 ;
        RECT 1546.605 1007.180 1547.370 1007.320 ;
        RECT 1546.605 1007.135 1546.895 1007.180 ;
        RECT 1547.050 1007.120 1547.370 1007.180 ;
        RECT 1546.605 917.900 1546.895 917.945 ;
        RECT 1547.510 917.900 1547.830 917.960 ;
        RECT 1546.605 917.760 1547.830 917.900 ;
        RECT 1546.605 917.715 1546.895 917.760 ;
        RECT 1547.510 917.700 1547.830 917.760 ;
        RECT 1547.510 870.100 1547.830 870.360 ;
        RECT 1547.600 869.340 1547.740 870.100 ;
        RECT 1547.510 869.080 1547.830 869.340 ;
        RECT 1546.590 738.180 1546.910 738.440 ;
        RECT 1546.680 738.040 1546.820 738.180 ;
        RECT 1547.050 738.040 1547.370 738.100 ;
        RECT 1546.680 737.900 1547.370 738.040 ;
        RECT 1547.050 737.840 1547.370 737.900 ;
        RECT 1547.050 717.640 1547.370 717.700 ;
        RECT 1548.430 717.640 1548.750 717.700 ;
        RECT 1547.050 717.500 1548.750 717.640 ;
        RECT 1547.050 717.440 1547.370 717.500 ;
        RECT 1548.430 717.440 1548.750 717.500 ;
        RECT 1547.510 620.740 1547.830 620.800 ;
        RECT 1547.510 620.600 1548.200 620.740 ;
        RECT 1547.510 620.540 1547.830 620.600 ;
        RECT 1546.590 620.060 1546.910 620.120 ;
        RECT 1548.060 620.060 1548.200 620.600 ;
        RECT 1546.590 619.920 1548.200 620.060 ;
        RECT 1546.590 619.860 1546.910 619.920 ;
        RECT 1546.130 531.320 1546.450 531.380 ;
        RECT 1546.590 531.320 1546.910 531.380 ;
        RECT 1546.130 531.180 1546.910 531.320 ;
        RECT 1546.130 531.120 1546.450 531.180 ;
        RECT 1546.590 531.120 1546.910 531.180 ;
        RECT 1546.130 524.180 1546.450 524.240 ;
        RECT 1545.935 524.040 1546.450 524.180 ;
        RECT 1546.130 523.980 1546.450 524.040 ;
        RECT 1546.145 448.360 1546.435 448.405 ;
        RECT 1546.590 448.360 1546.910 448.420 ;
        RECT 1546.145 448.220 1546.910 448.360 ;
        RECT 1546.145 448.175 1546.435 448.220 ;
        RECT 1546.590 448.160 1546.910 448.220 ;
        RECT 1546.590 400.420 1546.910 400.480 ;
        RECT 1546.395 400.280 1546.910 400.420 ;
        RECT 1546.590 400.220 1546.910 400.280 ;
        RECT 1546.130 386.480 1546.450 386.540 ;
        RECT 1546.605 386.480 1546.895 386.525 ;
        RECT 1546.130 386.340 1546.895 386.480 ;
        RECT 1546.130 386.280 1546.450 386.340 ;
        RECT 1546.605 386.295 1546.895 386.340 ;
        RECT 1546.130 338.340 1546.450 338.600 ;
        RECT 1546.220 338.200 1546.360 338.340 ;
        RECT 1546.590 338.200 1546.910 338.260 ;
        RECT 1546.220 338.060 1546.910 338.200 ;
        RECT 1546.590 338.000 1546.910 338.060 ;
        RECT 1546.590 255.380 1546.910 255.640 ;
        RECT 1546.680 254.900 1546.820 255.380 ;
        RECT 1547.050 254.900 1547.370 254.960 ;
        RECT 1546.680 254.760 1547.370 254.900 ;
        RECT 1547.050 254.700 1547.370 254.760 ;
        RECT 1546.605 234.500 1546.895 234.545 ;
        RECT 1547.050 234.500 1547.370 234.560 ;
        RECT 1546.605 234.360 1547.370 234.500 ;
        RECT 1546.605 234.315 1546.895 234.360 ;
        RECT 1547.050 234.300 1547.370 234.360 ;
        RECT 1546.590 186.560 1546.910 186.620 ;
        RECT 1546.395 186.420 1546.910 186.560 ;
        RECT 1546.590 186.360 1546.910 186.420 ;
        RECT 786.210 71.640 786.530 71.700 ;
        RECT 1546.590 71.640 1546.910 71.700 ;
        RECT 786.210 71.500 1546.910 71.640 ;
        RECT 786.210 71.440 786.530 71.500 ;
        RECT 1546.590 71.440 1546.910 71.500 ;
      LAYER via ;
        RECT 1547.080 1642.240 1547.340 1642.500 ;
        RECT 1548.460 1642.240 1548.720 1642.500 ;
        RECT 1546.620 1545.340 1546.880 1545.600 ;
        RECT 1547.080 1497.400 1547.340 1497.660 ;
        RECT 1546.620 1449.120 1546.880 1449.380 ;
        RECT 1548.000 1449.120 1548.260 1449.380 ;
        RECT 1546.620 1448.440 1546.880 1448.700 ;
        RECT 1547.080 1400.840 1547.340 1401.100 ;
        RECT 1546.620 1352.560 1546.880 1352.820 ;
        RECT 1548.000 1352.560 1548.260 1352.820 ;
        RECT 1546.620 1351.880 1546.880 1352.140 ;
        RECT 1547.080 1304.280 1547.340 1304.540 ;
        RECT 1547.080 1303.600 1547.340 1303.860 ;
        RECT 1546.620 1256.000 1546.880 1256.260 ;
        RECT 1547.540 1207.380 1547.800 1207.640 ;
        RECT 1548.000 1207.380 1548.260 1207.640 ;
        RECT 1546.620 1172.700 1546.880 1172.960 ;
        RECT 1548.000 1172.700 1548.260 1172.960 ;
        RECT 1546.620 1158.760 1546.880 1159.020 ;
        RECT 1547.540 1110.820 1547.800 1111.080 ;
        RECT 1546.620 1014.600 1546.880 1014.860 ;
        RECT 1547.080 1014.600 1547.340 1014.860 ;
        RECT 1547.080 1007.120 1547.340 1007.380 ;
        RECT 1547.540 917.700 1547.800 917.960 ;
        RECT 1547.540 870.100 1547.800 870.360 ;
        RECT 1547.540 869.080 1547.800 869.340 ;
        RECT 1546.620 738.180 1546.880 738.440 ;
        RECT 1547.080 737.840 1547.340 738.100 ;
        RECT 1547.080 717.440 1547.340 717.700 ;
        RECT 1548.460 717.440 1548.720 717.700 ;
        RECT 1547.540 620.540 1547.800 620.800 ;
        RECT 1546.620 619.860 1546.880 620.120 ;
        RECT 1546.160 531.120 1546.420 531.380 ;
        RECT 1546.620 531.120 1546.880 531.380 ;
        RECT 1546.160 523.980 1546.420 524.240 ;
        RECT 1546.620 448.160 1546.880 448.420 ;
        RECT 1546.620 400.220 1546.880 400.480 ;
        RECT 1546.160 386.280 1546.420 386.540 ;
        RECT 1546.160 338.340 1546.420 338.600 ;
        RECT 1546.620 338.000 1546.880 338.260 ;
        RECT 1546.620 255.380 1546.880 255.640 ;
        RECT 1547.080 254.700 1547.340 254.960 ;
        RECT 1547.080 234.300 1547.340 234.560 ;
        RECT 1546.620 186.360 1546.880 186.620 ;
        RECT 786.240 71.440 786.500 71.700 ;
        RECT 1546.620 71.440 1546.880 71.700 ;
      LAYER met2 ;
        RECT 1550.680 1700.410 1550.960 1704.000 ;
        RECT 1548.520 1700.270 1550.960 1700.410 ;
        RECT 1548.520 1642.530 1548.660 1700.270 ;
        RECT 1550.680 1700.000 1550.960 1700.270 ;
        RECT 1547.080 1642.210 1547.340 1642.530 ;
        RECT 1548.460 1642.210 1548.720 1642.530 ;
        RECT 1547.140 1559.650 1547.280 1642.210 ;
        RECT 1546.680 1559.510 1547.280 1559.650 ;
        RECT 1546.680 1545.630 1546.820 1559.510 ;
        RECT 1546.620 1545.310 1546.880 1545.630 ;
        RECT 1547.080 1497.370 1547.340 1497.690 ;
        RECT 1547.140 1497.205 1547.280 1497.370 ;
        RECT 1547.070 1496.835 1547.350 1497.205 ;
        RECT 1547.990 1496.835 1548.270 1497.205 ;
        RECT 1548.060 1449.410 1548.200 1496.835 ;
        RECT 1546.620 1449.090 1546.880 1449.410 ;
        RECT 1548.000 1449.090 1548.260 1449.410 ;
        RECT 1546.680 1448.730 1546.820 1449.090 ;
        RECT 1546.620 1448.410 1546.880 1448.730 ;
        RECT 1547.080 1400.810 1547.340 1401.130 ;
        RECT 1547.140 1400.645 1547.280 1400.810 ;
        RECT 1547.070 1400.275 1547.350 1400.645 ;
        RECT 1547.990 1400.275 1548.270 1400.645 ;
        RECT 1548.060 1352.850 1548.200 1400.275 ;
        RECT 1546.620 1352.530 1546.880 1352.850 ;
        RECT 1548.000 1352.530 1548.260 1352.850 ;
        RECT 1546.680 1352.170 1546.820 1352.530 ;
        RECT 1546.620 1351.850 1546.880 1352.170 ;
        RECT 1547.080 1304.250 1547.340 1304.570 ;
        RECT 1547.140 1303.890 1547.280 1304.250 ;
        RECT 1547.080 1303.570 1547.340 1303.890 ;
        RECT 1546.620 1255.970 1546.880 1256.290 ;
        RECT 1546.680 1255.805 1546.820 1255.970 ;
        RECT 1546.610 1255.435 1546.890 1255.805 ;
        RECT 1547.530 1255.435 1547.810 1255.805 ;
        RECT 1547.600 1207.670 1547.740 1255.435 ;
        RECT 1547.540 1207.350 1547.800 1207.670 ;
        RECT 1548.000 1207.350 1548.260 1207.670 ;
        RECT 1548.060 1172.990 1548.200 1207.350 ;
        RECT 1546.620 1172.670 1546.880 1172.990 ;
        RECT 1548.000 1172.670 1548.260 1172.990 ;
        RECT 1546.680 1159.050 1546.820 1172.670 ;
        RECT 1546.620 1158.730 1546.880 1159.050 ;
        RECT 1547.540 1110.790 1547.800 1111.110 ;
        RECT 1547.600 1055.885 1547.740 1110.790 ;
        RECT 1546.610 1055.515 1546.890 1055.885 ;
        RECT 1547.530 1055.515 1547.810 1055.885 ;
        RECT 1546.680 1014.890 1546.820 1055.515 ;
        RECT 1546.620 1014.570 1546.880 1014.890 ;
        RECT 1547.080 1014.570 1547.340 1014.890 ;
        RECT 1547.140 1007.410 1547.280 1014.570 ;
        RECT 1547.080 1007.090 1547.340 1007.410 ;
        RECT 1547.540 917.670 1547.800 917.990 ;
        RECT 1547.600 870.390 1547.740 917.670 ;
        RECT 1547.540 870.070 1547.800 870.390 ;
        RECT 1547.540 869.050 1547.800 869.370 ;
        RECT 1547.600 773.685 1547.740 869.050 ;
        RECT 1547.530 773.315 1547.810 773.685 ;
        RECT 1546.610 772.635 1546.890 773.005 ;
        RECT 1546.680 738.470 1546.820 772.635 ;
        RECT 1546.620 738.150 1546.880 738.470 ;
        RECT 1547.080 737.810 1547.340 738.130 ;
        RECT 1547.140 717.730 1547.280 737.810 ;
        RECT 1547.080 717.410 1547.340 717.730 ;
        RECT 1548.460 717.410 1548.720 717.730 ;
        RECT 1548.520 669.645 1548.660 717.410 ;
        RECT 1547.530 669.275 1547.810 669.645 ;
        RECT 1548.450 669.275 1548.730 669.645 ;
        RECT 1547.600 620.830 1547.740 669.275 ;
        RECT 1547.540 620.510 1547.800 620.830 ;
        RECT 1546.620 619.830 1546.880 620.150 ;
        RECT 1546.680 531.410 1546.820 619.830 ;
        RECT 1546.160 531.090 1546.420 531.410 ;
        RECT 1546.620 531.090 1546.880 531.410 ;
        RECT 1546.220 524.270 1546.360 531.090 ;
        RECT 1546.160 523.950 1546.420 524.270 ;
        RECT 1546.620 448.130 1546.880 448.450 ;
        RECT 1546.680 400.510 1546.820 448.130 ;
        RECT 1546.620 400.190 1546.880 400.510 ;
        RECT 1546.160 386.250 1546.420 386.570 ;
        RECT 1546.220 338.630 1546.360 386.250 ;
        RECT 1546.160 338.310 1546.420 338.630 ;
        RECT 1546.620 337.970 1546.880 338.290 ;
        RECT 1546.680 255.670 1546.820 337.970 ;
        RECT 1546.620 255.350 1546.880 255.670 ;
        RECT 1547.080 254.670 1547.340 254.990 ;
        RECT 1547.140 234.590 1547.280 254.670 ;
        RECT 1547.080 234.270 1547.340 234.590 ;
        RECT 1546.620 186.330 1546.880 186.650 ;
        RECT 1546.680 137.770 1546.820 186.330 ;
        RECT 1546.680 137.630 1547.280 137.770 ;
        RECT 1547.140 90.965 1547.280 137.630 ;
        RECT 1547.070 90.595 1547.350 90.965 ;
        RECT 1546.610 89.915 1546.890 90.285 ;
        RECT 1546.680 71.730 1546.820 89.915 ;
        RECT 786.240 71.410 786.500 71.730 ;
        RECT 1546.620 71.410 1546.880 71.730 ;
        RECT 786.300 16.730 786.440 71.410 ;
        RECT 781.700 16.590 786.440 16.730 ;
        RECT 781.700 2.400 781.840 16.590 ;
        RECT 781.490 -4.800 782.050 2.400 ;
      LAYER via2 ;
        RECT 1547.070 1496.880 1547.350 1497.160 ;
        RECT 1547.990 1496.880 1548.270 1497.160 ;
        RECT 1547.070 1400.320 1547.350 1400.600 ;
        RECT 1547.990 1400.320 1548.270 1400.600 ;
        RECT 1546.610 1255.480 1546.890 1255.760 ;
        RECT 1547.530 1255.480 1547.810 1255.760 ;
        RECT 1546.610 1055.560 1546.890 1055.840 ;
        RECT 1547.530 1055.560 1547.810 1055.840 ;
        RECT 1547.530 773.360 1547.810 773.640 ;
        RECT 1546.610 772.680 1546.890 772.960 ;
        RECT 1547.530 669.320 1547.810 669.600 ;
        RECT 1548.450 669.320 1548.730 669.600 ;
        RECT 1547.070 90.640 1547.350 90.920 ;
        RECT 1546.610 89.960 1546.890 90.240 ;
      LAYER met3 ;
        RECT 1547.045 1497.170 1547.375 1497.185 ;
        RECT 1547.965 1497.170 1548.295 1497.185 ;
        RECT 1547.045 1496.870 1548.295 1497.170 ;
        RECT 1547.045 1496.855 1547.375 1496.870 ;
        RECT 1547.965 1496.855 1548.295 1496.870 ;
        RECT 1547.045 1400.610 1547.375 1400.625 ;
        RECT 1547.965 1400.610 1548.295 1400.625 ;
        RECT 1547.045 1400.310 1548.295 1400.610 ;
        RECT 1547.045 1400.295 1547.375 1400.310 ;
        RECT 1547.965 1400.295 1548.295 1400.310 ;
        RECT 1546.585 1255.770 1546.915 1255.785 ;
        RECT 1547.505 1255.770 1547.835 1255.785 ;
        RECT 1546.585 1255.470 1547.835 1255.770 ;
        RECT 1546.585 1255.455 1546.915 1255.470 ;
        RECT 1547.505 1255.455 1547.835 1255.470 ;
        RECT 1546.585 1055.850 1546.915 1055.865 ;
        RECT 1547.505 1055.850 1547.835 1055.865 ;
        RECT 1546.585 1055.550 1547.835 1055.850 ;
        RECT 1546.585 1055.535 1546.915 1055.550 ;
        RECT 1547.505 1055.535 1547.835 1055.550 ;
        RECT 1547.505 773.650 1547.835 773.665 ;
        RECT 1545.910 773.350 1547.835 773.650 ;
        RECT 1545.910 772.970 1546.210 773.350 ;
        RECT 1547.505 773.335 1547.835 773.350 ;
        RECT 1546.585 772.970 1546.915 772.985 ;
        RECT 1545.910 772.670 1546.915 772.970 ;
        RECT 1546.585 772.655 1546.915 772.670 ;
        RECT 1547.505 669.610 1547.835 669.625 ;
        RECT 1548.425 669.610 1548.755 669.625 ;
        RECT 1547.505 669.310 1548.755 669.610 ;
        RECT 1547.505 669.295 1547.835 669.310 ;
        RECT 1548.425 669.295 1548.755 669.310 ;
        RECT 1547.045 90.930 1547.375 90.945 ;
        RECT 1545.910 90.630 1547.375 90.930 ;
        RECT 1545.910 90.250 1546.210 90.630 ;
        RECT 1547.045 90.615 1547.375 90.630 ;
        RECT 1546.585 90.250 1546.915 90.265 ;
        RECT 1545.910 89.950 1546.915 90.250 ;
        RECT 1546.585 89.935 1546.915 89.950 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2266.490 1686.980 2266.810 1687.040 ;
        RECT 2303.750 1686.980 2304.070 1687.040 ;
        RECT 2266.490 1686.840 2304.070 1686.980 ;
        RECT 2266.490 1686.780 2266.810 1686.840 ;
        RECT 2303.750 1686.780 2304.070 1686.840 ;
        RECT 2244.870 19.280 2245.190 19.340 ;
        RECT 2266.490 19.280 2266.810 19.340 ;
        RECT 2244.870 19.140 2266.810 19.280 ;
        RECT 2244.870 19.080 2245.190 19.140 ;
        RECT 2266.490 19.080 2266.810 19.140 ;
      LAYER via ;
        RECT 2266.520 1686.780 2266.780 1687.040 ;
        RECT 2303.780 1686.780 2304.040 1687.040 ;
        RECT 2244.900 19.080 2245.160 19.340 ;
        RECT 2266.520 19.080 2266.780 19.340 ;
      LAYER met2 ;
        RECT 2303.700 1700.000 2303.980 1704.000 ;
        RECT 2303.840 1687.070 2303.980 1700.000 ;
        RECT 2266.520 1686.750 2266.780 1687.070 ;
        RECT 2303.780 1686.750 2304.040 1687.070 ;
        RECT 2266.580 19.370 2266.720 1686.750 ;
        RECT 2244.900 19.050 2245.160 19.370 ;
        RECT 2266.520 19.050 2266.780 19.370 ;
        RECT 2244.960 2.400 2245.100 19.050 ;
        RECT 2244.750 -4.800 2245.310 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2300.990 1683.920 2301.310 1683.980 ;
        RECT 2312.950 1683.920 2313.270 1683.980 ;
        RECT 2300.990 1683.780 2313.270 1683.920 ;
        RECT 2300.990 1683.720 2301.310 1683.780 ;
        RECT 2312.950 1683.720 2313.270 1683.780 ;
        RECT 2262.350 17.580 2262.670 17.640 ;
        RECT 2300.990 17.580 2301.310 17.640 ;
        RECT 2262.350 17.440 2301.310 17.580 ;
        RECT 2262.350 17.380 2262.670 17.440 ;
        RECT 2300.990 17.380 2301.310 17.440 ;
      LAYER via ;
        RECT 2301.020 1683.720 2301.280 1683.980 ;
        RECT 2312.980 1683.720 2313.240 1683.980 ;
        RECT 2262.380 17.380 2262.640 17.640 ;
        RECT 2301.020 17.380 2301.280 17.640 ;
      LAYER met2 ;
        RECT 2312.900 1700.000 2313.180 1704.000 ;
        RECT 2313.040 1684.010 2313.180 1700.000 ;
        RECT 2301.020 1683.690 2301.280 1684.010 ;
        RECT 2312.980 1683.690 2313.240 1684.010 ;
        RECT 2301.080 17.670 2301.220 1683.690 ;
        RECT 2262.380 17.350 2262.640 17.670 ;
        RECT 2301.020 17.350 2301.280 17.670 ;
        RECT 2262.440 2.400 2262.580 17.350 ;
        RECT 2262.230 -4.800 2262.790 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2314.790 1684.600 2315.110 1684.660 ;
        RECT 2322.150 1684.600 2322.470 1684.660 ;
        RECT 2314.790 1684.460 2322.470 1684.600 ;
        RECT 2314.790 1684.400 2315.110 1684.460 ;
        RECT 2322.150 1684.400 2322.470 1684.460 ;
        RECT 2280.750 19.960 2281.070 20.020 ;
        RECT 2314.790 19.960 2315.110 20.020 ;
        RECT 2280.750 19.820 2315.110 19.960 ;
        RECT 2280.750 19.760 2281.070 19.820 ;
        RECT 2314.790 19.760 2315.110 19.820 ;
      LAYER via ;
        RECT 2314.820 1684.400 2315.080 1684.660 ;
        RECT 2322.180 1684.400 2322.440 1684.660 ;
        RECT 2280.780 19.760 2281.040 20.020 ;
        RECT 2314.820 19.760 2315.080 20.020 ;
      LAYER met2 ;
        RECT 2322.100 1700.000 2322.380 1704.000 ;
        RECT 2322.240 1684.690 2322.380 1700.000 ;
        RECT 2314.820 1684.370 2315.080 1684.690 ;
        RECT 2322.180 1684.370 2322.440 1684.690 ;
        RECT 2314.880 20.050 2315.020 1684.370 ;
        RECT 2280.780 19.730 2281.040 20.050 ;
        RECT 2314.820 19.730 2315.080 20.050 ;
        RECT 2280.840 9.930 2280.980 19.730 ;
        RECT 2280.380 9.790 2280.980 9.930 ;
        RECT 2280.380 2.400 2280.520 9.790 ;
        RECT 2280.170 -4.800 2280.730 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2321.690 1684.940 2322.010 1685.000 ;
        RECT 2331.350 1684.940 2331.670 1685.000 ;
        RECT 2321.690 1684.800 2331.670 1684.940 ;
        RECT 2321.690 1684.740 2322.010 1684.800 ;
        RECT 2331.350 1684.740 2331.670 1684.800 ;
        RECT 2298.230 18.940 2298.550 19.000 ;
        RECT 2321.690 18.940 2322.010 19.000 ;
        RECT 2298.230 18.800 2322.010 18.940 ;
        RECT 2298.230 18.740 2298.550 18.800 ;
        RECT 2321.690 18.740 2322.010 18.800 ;
      LAYER via ;
        RECT 2321.720 1684.740 2321.980 1685.000 ;
        RECT 2331.380 1684.740 2331.640 1685.000 ;
        RECT 2298.260 18.740 2298.520 19.000 ;
        RECT 2321.720 18.740 2321.980 19.000 ;
      LAYER met2 ;
        RECT 2331.300 1700.000 2331.580 1704.000 ;
        RECT 2331.440 1685.030 2331.580 1700.000 ;
        RECT 2321.720 1684.710 2321.980 1685.030 ;
        RECT 2331.380 1684.710 2331.640 1685.030 ;
        RECT 2321.780 19.030 2321.920 1684.710 ;
        RECT 2298.260 18.710 2298.520 19.030 ;
        RECT 2321.720 18.710 2321.980 19.030 ;
        RECT 2298.320 2.400 2298.460 18.710 ;
        RECT 2298.110 -4.800 2298.670 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2318.010 1689.020 2318.330 1689.080 ;
        RECT 2340.550 1689.020 2340.870 1689.080 ;
        RECT 2318.010 1688.880 2340.870 1689.020 ;
        RECT 2318.010 1688.820 2318.330 1688.880 ;
        RECT 2340.550 1688.820 2340.870 1688.880 ;
      LAYER via ;
        RECT 2318.040 1688.820 2318.300 1689.080 ;
        RECT 2340.580 1688.820 2340.840 1689.080 ;
      LAYER met2 ;
        RECT 2340.500 1700.000 2340.780 1704.000 ;
        RECT 2340.640 1689.110 2340.780 1700.000 ;
        RECT 2318.040 1688.790 2318.300 1689.110 ;
        RECT 2340.580 1688.790 2340.840 1689.110 ;
        RECT 2318.100 16.730 2318.240 1688.790 ;
        RECT 2316.260 16.590 2318.240 16.730 ;
        RECT 2316.260 2.400 2316.400 16.590 ;
        RECT 2316.050 -4.800 2316.610 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2338.710 1684.260 2339.030 1684.320 ;
        RECT 2349.750 1684.260 2350.070 1684.320 ;
        RECT 2338.710 1684.120 2350.070 1684.260 ;
        RECT 2338.710 1684.060 2339.030 1684.120 ;
        RECT 2349.750 1684.060 2350.070 1684.120 ;
        RECT 2334.110 18.600 2334.430 18.660 ;
        RECT 2338.710 18.600 2339.030 18.660 ;
        RECT 2334.110 18.460 2339.030 18.600 ;
        RECT 2334.110 18.400 2334.430 18.460 ;
        RECT 2338.710 18.400 2339.030 18.460 ;
      LAYER via ;
        RECT 2338.740 1684.060 2339.000 1684.320 ;
        RECT 2349.780 1684.060 2350.040 1684.320 ;
        RECT 2334.140 18.400 2334.400 18.660 ;
        RECT 2338.740 18.400 2339.000 18.660 ;
      LAYER met2 ;
        RECT 2349.700 1700.000 2349.980 1704.000 ;
        RECT 2349.840 1684.350 2349.980 1700.000 ;
        RECT 2338.740 1684.030 2339.000 1684.350 ;
        RECT 2349.780 1684.030 2350.040 1684.350 ;
        RECT 2338.800 18.690 2338.940 1684.030 ;
        RECT 2334.140 18.370 2334.400 18.690 ;
        RECT 2338.740 18.370 2339.000 18.690 ;
        RECT 2334.200 2.400 2334.340 18.370 ;
        RECT 2333.990 -4.800 2334.550 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2351.590 20.640 2351.910 20.700 ;
        RECT 2353.890 20.640 2354.210 20.700 ;
        RECT 2351.590 20.500 2354.210 20.640 ;
        RECT 2351.590 20.440 2351.910 20.500 ;
        RECT 2353.890 20.440 2354.210 20.500 ;
      LAYER via ;
        RECT 2351.620 20.440 2351.880 20.700 ;
        RECT 2353.920 20.440 2354.180 20.700 ;
      LAYER met2 ;
        RECT 2358.900 1700.410 2359.180 1704.000 ;
        RECT 2356.740 1700.270 2359.180 1700.410 ;
        RECT 2356.740 1678.650 2356.880 1700.270 ;
        RECT 2358.900 1700.000 2359.180 1700.270 ;
        RECT 2353.980 1678.510 2356.880 1678.650 ;
        RECT 2353.980 20.730 2354.120 1678.510 ;
        RECT 2351.620 20.410 2351.880 20.730 ;
        RECT 2353.920 20.410 2354.180 20.730 ;
        RECT 2351.680 2.400 2351.820 20.410 ;
        RECT 2351.470 -4.800 2352.030 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2366.770 20.640 2367.090 20.700 ;
        RECT 2369.530 20.640 2369.850 20.700 ;
        RECT 2366.770 20.500 2369.850 20.640 ;
        RECT 2366.770 20.440 2367.090 20.500 ;
        RECT 2369.530 20.440 2369.850 20.500 ;
      LAYER via ;
        RECT 2366.800 20.440 2367.060 20.700 ;
        RECT 2369.560 20.440 2369.820 20.700 ;
      LAYER met2 ;
        RECT 2368.100 1700.410 2368.380 1704.000 ;
        RECT 2366.860 1700.270 2368.380 1700.410 ;
        RECT 2366.860 20.730 2367.000 1700.270 ;
        RECT 2368.100 1700.000 2368.380 1700.270 ;
        RECT 2366.800 20.410 2367.060 20.730 ;
        RECT 2369.560 20.410 2369.820 20.730 ;
        RECT 2369.620 2.400 2369.760 20.410 ;
        RECT 2369.410 -4.800 2369.970 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2377.350 1688.340 2377.670 1688.400 ;
        RECT 2388.390 1688.340 2388.710 1688.400 ;
        RECT 2377.350 1688.200 2388.710 1688.340 ;
        RECT 2377.350 1688.140 2377.670 1688.200 ;
        RECT 2388.390 1688.140 2388.710 1688.200 ;
      LAYER via ;
        RECT 2377.380 1688.140 2377.640 1688.400 ;
        RECT 2388.420 1688.140 2388.680 1688.400 ;
      LAYER met2 ;
        RECT 2377.300 1700.000 2377.580 1704.000 ;
        RECT 2377.440 1688.430 2377.580 1700.000 ;
        RECT 2377.380 1688.110 2377.640 1688.430 ;
        RECT 2388.420 1688.110 2388.680 1688.430 ;
        RECT 2388.480 37.130 2388.620 1688.110 ;
        RECT 2387.560 36.990 2388.620 37.130 ;
        RECT 2387.560 2.400 2387.700 36.990 ;
        RECT 2387.350 -4.800 2387.910 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2401.805 1538.925 2401.975 1587.035 ;
        RECT 2401.805 1442.025 2401.975 1490.475 ;
        RECT 2401.345 1007.505 2401.515 1014.815 ;
        RECT 2401.345 766.105 2401.515 821.015 ;
        RECT 2402.265 476.085 2402.435 524.195 ;
        RECT 2402.265 385.645 2402.435 427.635 ;
        RECT 2401.805 89.845 2401.975 137.955 ;
      LAYER mcon ;
        RECT 2401.805 1586.865 2401.975 1587.035 ;
        RECT 2401.805 1490.305 2401.975 1490.475 ;
        RECT 2401.345 1014.645 2401.515 1014.815 ;
        RECT 2401.345 820.845 2401.515 821.015 ;
        RECT 2402.265 524.025 2402.435 524.195 ;
        RECT 2402.265 427.465 2402.435 427.635 ;
        RECT 2401.805 137.785 2401.975 137.955 ;
      LAYER met1 ;
        RECT 2386.550 1635.640 2386.870 1635.700 ;
        RECT 2401.730 1635.640 2402.050 1635.700 ;
        RECT 2386.550 1635.500 2402.050 1635.640 ;
        RECT 2386.550 1635.440 2386.870 1635.500 ;
        RECT 2401.730 1635.440 2402.050 1635.500 ;
        RECT 2401.730 1587.020 2402.050 1587.080 ;
        RECT 2401.535 1586.880 2402.050 1587.020 ;
        RECT 2401.730 1586.820 2402.050 1586.880 ;
        RECT 2401.730 1539.080 2402.050 1539.140 ;
        RECT 2401.535 1538.940 2402.050 1539.080 ;
        RECT 2401.730 1538.880 2402.050 1538.940 ;
        RECT 2401.730 1490.460 2402.050 1490.520 ;
        RECT 2401.535 1490.320 2402.050 1490.460 ;
        RECT 2401.730 1490.260 2402.050 1490.320 ;
        RECT 2401.730 1442.180 2402.050 1442.240 ;
        RECT 2401.535 1442.040 2402.050 1442.180 ;
        RECT 2401.730 1441.980 2402.050 1442.040 ;
        RECT 2400.810 1345.620 2401.130 1345.680 ;
        RECT 2401.730 1345.620 2402.050 1345.680 ;
        RECT 2400.810 1345.480 2402.050 1345.620 ;
        RECT 2400.810 1345.420 2401.130 1345.480 ;
        RECT 2401.730 1345.420 2402.050 1345.480 ;
        RECT 2400.810 1249.060 2401.130 1249.120 ;
        RECT 2401.730 1249.060 2402.050 1249.120 ;
        RECT 2400.810 1248.920 2402.050 1249.060 ;
        RECT 2400.810 1248.860 2401.130 1248.920 ;
        RECT 2401.730 1248.860 2402.050 1248.920 ;
        RECT 2400.810 1152.500 2401.130 1152.560 ;
        RECT 2401.730 1152.500 2402.050 1152.560 ;
        RECT 2400.810 1152.360 2402.050 1152.500 ;
        RECT 2400.810 1152.300 2401.130 1152.360 ;
        RECT 2401.730 1152.300 2402.050 1152.360 ;
        RECT 2401.285 1014.800 2401.575 1014.845 ;
        RECT 2401.730 1014.800 2402.050 1014.860 ;
        RECT 2401.285 1014.660 2402.050 1014.800 ;
        RECT 2401.285 1014.615 2401.575 1014.660 ;
        RECT 2401.730 1014.600 2402.050 1014.660 ;
        RECT 2401.270 1007.660 2401.590 1007.720 ;
        RECT 2401.075 1007.520 2401.590 1007.660 ;
        RECT 2401.270 1007.460 2401.590 1007.520 ;
        RECT 2401.270 979.920 2401.590 980.180 ;
        RECT 2401.360 979.440 2401.500 979.920 ;
        RECT 2401.730 979.440 2402.050 979.500 ;
        RECT 2401.360 979.300 2402.050 979.440 ;
        RECT 2401.730 979.240 2402.050 979.300 ;
        RECT 2401.730 893.900 2402.050 894.160 ;
        RECT 2401.820 893.480 2401.960 893.900 ;
        RECT 2401.730 893.220 2402.050 893.480 ;
        RECT 2401.730 845.480 2402.050 845.540 ;
        RECT 2402.650 845.480 2402.970 845.540 ;
        RECT 2401.730 845.340 2402.970 845.480 ;
        RECT 2401.730 845.280 2402.050 845.340 ;
        RECT 2402.650 845.280 2402.970 845.340 ;
        RECT 2401.285 821.000 2401.575 821.045 ;
        RECT 2401.730 821.000 2402.050 821.060 ;
        RECT 2401.285 820.860 2402.050 821.000 ;
        RECT 2401.285 820.815 2401.575 820.860 ;
        RECT 2401.730 820.800 2402.050 820.860 ;
        RECT 2401.270 766.260 2401.590 766.320 ;
        RECT 2401.075 766.120 2401.590 766.260 ;
        RECT 2401.270 766.060 2401.590 766.120 ;
        RECT 2401.270 717.640 2401.590 717.700 ;
        RECT 2402.190 717.640 2402.510 717.700 ;
        RECT 2401.270 717.500 2402.510 717.640 ;
        RECT 2401.270 717.440 2401.590 717.500 ;
        RECT 2402.190 717.440 2402.510 717.500 ;
        RECT 2402.190 524.180 2402.510 524.240 ;
        RECT 2401.995 524.040 2402.510 524.180 ;
        RECT 2402.190 523.980 2402.510 524.040 ;
        RECT 2402.205 476.240 2402.495 476.285 ;
        RECT 2402.650 476.240 2402.970 476.300 ;
        RECT 2402.205 476.100 2402.970 476.240 ;
        RECT 2402.205 476.055 2402.495 476.100 ;
        RECT 2402.650 476.040 2402.970 476.100 ;
        RECT 2402.190 427.620 2402.510 427.680 ;
        RECT 2401.995 427.480 2402.510 427.620 ;
        RECT 2402.190 427.420 2402.510 427.480 ;
        RECT 2402.205 385.800 2402.495 385.845 ;
        RECT 2402.650 385.800 2402.970 385.860 ;
        RECT 2402.205 385.660 2402.970 385.800 ;
        RECT 2402.205 385.615 2402.495 385.660 ;
        RECT 2402.650 385.600 2402.970 385.660 ;
        RECT 2401.270 337.860 2401.590 337.920 ;
        RECT 2402.190 337.860 2402.510 337.920 ;
        RECT 2401.270 337.720 2402.510 337.860 ;
        RECT 2401.270 337.660 2401.590 337.720 ;
        RECT 2402.190 337.660 2402.510 337.720 ;
        RECT 2401.730 289.580 2402.050 289.640 ;
        RECT 2402.650 289.580 2402.970 289.640 ;
        RECT 2401.730 289.440 2402.970 289.580 ;
        RECT 2401.730 289.380 2402.050 289.440 ;
        RECT 2402.650 289.380 2402.970 289.440 ;
        RECT 2401.270 193.700 2401.590 193.760 ;
        RECT 2402.650 193.700 2402.970 193.760 ;
        RECT 2401.270 193.560 2402.970 193.700 ;
        RECT 2401.270 193.500 2401.590 193.560 ;
        RECT 2402.650 193.500 2402.970 193.560 ;
        RECT 2401.270 158.820 2401.590 159.080 ;
        RECT 2401.360 158.340 2401.500 158.820 ;
        RECT 2401.730 158.340 2402.050 158.400 ;
        RECT 2401.360 158.200 2402.050 158.340 ;
        RECT 2401.730 158.140 2402.050 158.200 ;
        RECT 2401.730 137.940 2402.050 138.000 ;
        RECT 2401.535 137.800 2402.050 137.940 ;
        RECT 2401.730 137.740 2402.050 137.800 ;
        RECT 2401.730 90.000 2402.050 90.060 ;
        RECT 2401.535 89.860 2402.050 90.000 ;
        RECT 2401.730 89.800 2402.050 89.860 ;
        RECT 2401.730 5.000 2402.050 5.060 ;
        RECT 2405.410 5.000 2405.730 5.060 ;
        RECT 2401.730 4.860 2405.730 5.000 ;
        RECT 2401.730 4.800 2402.050 4.860 ;
        RECT 2405.410 4.800 2405.730 4.860 ;
      LAYER via ;
        RECT 2386.580 1635.440 2386.840 1635.700 ;
        RECT 2401.760 1635.440 2402.020 1635.700 ;
        RECT 2401.760 1586.820 2402.020 1587.080 ;
        RECT 2401.760 1538.880 2402.020 1539.140 ;
        RECT 2401.760 1490.260 2402.020 1490.520 ;
        RECT 2401.760 1441.980 2402.020 1442.240 ;
        RECT 2400.840 1345.420 2401.100 1345.680 ;
        RECT 2401.760 1345.420 2402.020 1345.680 ;
        RECT 2400.840 1248.860 2401.100 1249.120 ;
        RECT 2401.760 1248.860 2402.020 1249.120 ;
        RECT 2400.840 1152.300 2401.100 1152.560 ;
        RECT 2401.760 1152.300 2402.020 1152.560 ;
        RECT 2401.760 1014.600 2402.020 1014.860 ;
        RECT 2401.300 1007.460 2401.560 1007.720 ;
        RECT 2401.300 979.920 2401.560 980.180 ;
        RECT 2401.760 979.240 2402.020 979.500 ;
        RECT 2401.760 893.900 2402.020 894.160 ;
        RECT 2401.760 893.220 2402.020 893.480 ;
        RECT 2401.760 845.280 2402.020 845.540 ;
        RECT 2402.680 845.280 2402.940 845.540 ;
        RECT 2401.760 820.800 2402.020 821.060 ;
        RECT 2401.300 766.060 2401.560 766.320 ;
        RECT 2401.300 717.440 2401.560 717.700 ;
        RECT 2402.220 717.440 2402.480 717.700 ;
        RECT 2402.220 523.980 2402.480 524.240 ;
        RECT 2402.680 476.040 2402.940 476.300 ;
        RECT 2402.220 427.420 2402.480 427.680 ;
        RECT 2402.680 385.600 2402.940 385.860 ;
        RECT 2401.300 337.660 2401.560 337.920 ;
        RECT 2402.220 337.660 2402.480 337.920 ;
        RECT 2401.760 289.380 2402.020 289.640 ;
        RECT 2402.680 289.380 2402.940 289.640 ;
        RECT 2401.300 193.500 2401.560 193.760 ;
        RECT 2402.680 193.500 2402.940 193.760 ;
        RECT 2401.300 158.820 2401.560 159.080 ;
        RECT 2401.760 158.140 2402.020 158.400 ;
        RECT 2401.760 137.740 2402.020 138.000 ;
        RECT 2401.760 89.800 2402.020 90.060 ;
        RECT 2401.760 4.800 2402.020 5.060 ;
        RECT 2405.440 4.800 2405.700 5.060 ;
      LAYER met2 ;
        RECT 2386.500 1700.000 2386.780 1704.000 ;
        RECT 2386.640 1635.730 2386.780 1700.000 ;
        RECT 2386.580 1635.410 2386.840 1635.730 ;
        RECT 2401.760 1635.410 2402.020 1635.730 ;
        RECT 2401.820 1587.110 2401.960 1635.410 ;
        RECT 2401.760 1586.790 2402.020 1587.110 ;
        RECT 2401.760 1538.850 2402.020 1539.170 ;
        RECT 2401.820 1490.550 2401.960 1538.850 ;
        RECT 2401.760 1490.230 2402.020 1490.550 ;
        RECT 2401.760 1441.950 2402.020 1442.270 ;
        RECT 2401.820 1393.845 2401.960 1441.950 ;
        RECT 2400.830 1393.475 2401.110 1393.845 ;
        RECT 2401.750 1393.475 2402.030 1393.845 ;
        RECT 2400.900 1345.710 2401.040 1393.475 ;
        RECT 2400.840 1345.390 2401.100 1345.710 ;
        RECT 2401.760 1345.390 2402.020 1345.710 ;
        RECT 2401.820 1297.285 2401.960 1345.390 ;
        RECT 2400.830 1296.915 2401.110 1297.285 ;
        RECT 2401.750 1296.915 2402.030 1297.285 ;
        RECT 2400.900 1249.150 2401.040 1296.915 ;
        RECT 2400.840 1248.830 2401.100 1249.150 ;
        RECT 2401.760 1248.830 2402.020 1249.150 ;
        RECT 2401.820 1208.885 2401.960 1248.830 ;
        RECT 2401.750 1208.515 2402.030 1208.885 ;
        RECT 2401.750 1207.835 2402.030 1208.205 ;
        RECT 2401.820 1200.725 2401.960 1207.835 ;
        RECT 2400.830 1200.355 2401.110 1200.725 ;
        RECT 2401.750 1200.355 2402.030 1200.725 ;
        RECT 2400.900 1152.590 2401.040 1200.355 ;
        RECT 2400.840 1152.270 2401.100 1152.590 ;
        RECT 2401.760 1152.270 2402.020 1152.590 ;
        RECT 2401.820 1104.165 2401.960 1152.270 ;
        RECT 2400.830 1103.795 2401.110 1104.165 ;
        RECT 2401.750 1103.795 2402.030 1104.165 ;
        RECT 2400.900 1055.885 2401.040 1103.795 ;
        RECT 2400.830 1055.515 2401.110 1055.885 ;
        RECT 2401.750 1055.515 2402.030 1055.885 ;
        RECT 2401.820 1014.890 2401.960 1055.515 ;
        RECT 2401.760 1014.570 2402.020 1014.890 ;
        RECT 2401.300 1007.430 2401.560 1007.750 ;
        RECT 2401.360 980.210 2401.500 1007.430 ;
        RECT 2401.300 979.890 2401.560 980.210 ;
        RECT 2401.760 979.210 2402.020 979.530 ;
        RECT 2401.820 931.330 2401.960 979.210 ;
        RECT 2401.820 931.190 2402.420 931.330 ;
        RECT 2402.280 917.730 2402.420 931.190 ;
        RECT 2401.820 917.590 2402.420 917.730 ;
        RECT 2401.820 894.190 2401.960 917.590 ;
        RECT 2401.760 893.870 2402.020 894.190 ;
        RECT 2401.760 893.190 2402.020 893.510 ;
        RECT 2401.820 845.570 2401.960 893.190 ;
        RECT 2401.760 845.250 2402.020 845.570 ;
        RECT 2402.680 845.250 2402.940 845.570 ;
        RECT 2402.740 821.285 2402.880 845.250 ;
        RECT 2401.750 820.915 2402.030 821.285 ;
        RECT 2402.670 820.915 2402.950 821.285 ;
        RECT 2401.760 820.770 2402.020 820.915 ;
        RECT 2401.300 766.030 2401.560 766.350 ;
        RECT 2401.360 717.730 2401.500 766.030 ;
        RECT 2401.300 717.410 2401.560 717.730 ;
        RECT 2402.220 717.410 2402.480 717.730 ;
        RECT 2402.280 579.885 2402.420 717.410 ;
        RECT 2401.290 579.515 2401.570 579.885 ;
        RECT 2402.210 579.515 2402.490 579.885 ;
        RECT 2401.360 555.290 2401.500 579.515 ;
        RECT 2401.360 555.150 2402.420 555.290 ;
        RECT 2402.280 524.270 2402.420 555.150 ;
        RECT 2402.220 523.950 2402.480 524.270 ;
        RECT 2402.680 476.010 2402.940 476.330 ;
        RECT 2402.740 448.530 2402.880 476.010 ;
        RECT 2402.280 448.390 2402.880 448.530 ;
        RECT 2402.280 427.710 2402.420 448.390 ;
        RECT 2402.220 427.390 2402.480 427.710 ;
        RECT 2402.680 385.570 2402.940 385.890 ;
        RECT 2402.740 338.370 2402.880 385.570 ;
        RECT 2402.280 338.230 2402.880 338.370 ;
        RECT 2402.280 337.950 2402.420 338.230 ;
        RECT 2401.300 337.630 2401.560 337.950 ;
        RECT 2402.220 337.630 2402.480 337.950 ;
        RECT 2401.360 290.090 2401.500 337.630 ;
        RECT 2401.360 289.950 2401.960 290.090 ;
        RECT 2401.820 289.670 2401.960 289.950 ;
        RECT 2401.760 289.350 2402.020 289.670 ;
        RECT 2402.680 289.350 2402.940 289.670 ;
        RECT 2402.740 193.790 2402.880 289.350 ;
        RECT 2401.300 193.470 2401.560 193.790 ;
        RECT 2402.680 193.470 2402.940 193.790 ;
        RECT 2401.360 159.110 2401.500 193.470 ;
        RECT 2401.300 158.790 2401.560 159.110 ;
        RECT 2401.760 158.110 2402.020 158.430 ;
        RECT 2401.820 138.030 2401.960 158.110 ;
        RECT 2401.760 137.710 2402.020 138.030 ;
        RECT 2401.760 89.770 2402.020 90.090 ;
        RECT 2401.820 5.090 2401.960 89.770 ;
        RECT 2401.760 4.770 2402.020 5.090 ;
        RECT 2405.440 4.770 2405.700 5.090 ;
        RECT 2405.500 2.400 2405.640 4.770 ;
        RECT 2405.290 -4.800 2405.850 2.400 ;
      LAYER via2 ;
        RECT 2400.830 1393.520 2401.110 1393.800 ;
        RECT 2401.750 1393.520 2402.030 1393.800 ;
        RECT 2400.830 1296.960 2401.110 1297.240 ;
        RECT 2401.750 1296.960 2402.030 1297.240 ;
        RECT 2401.750 1208.560 2402.030 1208.840 ;
        RECT 2401.750 1207.880 2402.030 1208.160 ;
        RECT 2400.830 1200.400 2401.110 1200.680 ;
        RECT 2401.750 1200.400 2402.030 1200.680 ;
        RECT 2400.830 1103.840 2401.110 1104.120 ;
        RECT 2401.750 1103.840 2402.030 1104.120 ;
        RECT 2400.830 1055.560 2401.110 1055.840 ;
        RECT 2401.750 1055.560 2402.030 1055.840 ;
        RECT 2401.750 820.960 2402.030 821.240 ;
        RECT 2402.670 820.960 2402.950 821.240 ;
        RECT 2401.290 579.560 2401.570 579.840 ;
        RECT 2402.210 579.560 2402.490 579.840 ;
      LAYER met3 ;
        RECT 2400.805 1393.810 2401.135 1393.825 ;
        RECT 2401.725 1393.810 2402.055 1393.825 ;
        RECT 2400.805 1393.510 2402.055 1393.810 ;
        RECT 2400.805 1393.495 2401.135 1393.510 ;
        RECT 2401.725 1393.495 2402.055 1393.510 ;
        RECT 2400.805 1297.250 2401.135 1297.265 ;
        RECT 2401.725 1297.250 2402.055 1297.265 ;
        RECT 2400.805 1296.950 2402.055 1297.250 ;
        RECT 2400.805 1296.935 2401.135 1296.950 ;
        RECT 2401.725 1296.935 2402.055 1296.950 ;
        RECT 2401.725 1208.850 2402.055 1208.865 ;
        RECT 2401.725 1208.550 2402.730 1208.850 ;
        RECT 2401.725 1208.535 2402.055 1208.550 ;
        RECT 2401.725 1208.170 2402.055 1208.185 ;
        RECT 2402.430 1208.170 2402.730 1208.550 ;
        RECT 2401.725 1207.870 2402.730 1208.170 ;
        RECT 2401.725 1207.855 2402.055 1207.870 ;
        RECT 2400.805 1200.690 2401.135 1200.705 ;
        RECT 2401.725 1200.690 2402.055 1200.705 ;
        RECT 2400.805 1200.390 2402.055 1200.690 ;
        RECT 2400.805 1200.375 2401.135 1200.390 ;
        RECT 2401.725 1200.375 2402.055 1200.390 ;
        RECT 2400.805 1104.130 2401.135 1104.145 ;
        RECT 2401.725 1104.130 2402.055 1104.145 ;
        RECT 2400.805 1103.830 2402.055 1104.130 ;
        RECT 2400.805 1103.815 2401.135 1103.830 ;
        RECT 2401.725 1103.815 2402.055 1103.830 ;
        RECT 2400.805 1055.850 2401.135 1055.865 ;
        RECT 2401.725 1055.850 2402.055 1055.865 ;
        RECT 2400.805 1055.550 2402.055 1055.850 ;
        RECT 2400.805 1055.535 2401.135 1055.550 ;
        RECT 2401.725 1055.535 2402.055 1055.550 ;
        RECT 2401.725 821.250 2402.055 821.265 ;
        RECT 2402.645 821.250 2402.975 821.265 ;
        RECT 2401.725 820.950 2402.975 821.250 ;
        RECT 2401.725 820.935 2402.055 820.950 ;
        RECT 2402.645 820.935 2402.975 820.950 ;
        RECT 2401.265 579.850 2401.595 579.865 ;
        RECT 2402.185 579.850 2402.515 579.865 ;
        RECT 2401.265 579.550 2402.515 579.850 ;
        RECT 2401.265 579.535 2401.595 579.550 ;
        RECT 2402.185 579.535 2402.515 579.550 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 800.010 71.980 800.330 72.040 ;
        RECT 1559.930 71.980 1560.250 72.040 ;
        RECT 800.010 71.840 1560.250 71.980 ;
        RECT 800.010 71.780 800.330 71.840 ;
        RECT 1559.930 71.780 1560.250 71.840 ;
      LAYER via ;
        RECT 800.040 71.780 800.300 72.040 ;
        RECT 1559.960 71.780 1560.220 72.040 ;
      LAYER met2 ;
        RECT 1559.880 1700.000 1560.160 1704.000 ;
        RECT 1560.020 72.070 1560.160 1700.000 ;
        RECT 800.040 71.750 800.300 72.070 ;
        RECT 1559.960 71.750 1560.220 72.070 ;
        RECT 800.100 17.410 800.240 71.750 ;
        RECT 799.640 17.270 800.240 17.410 ;
        RECT 799.640 2.400 799.780 17.270 ;
        RECT 799.430 -4.800 799.990 2.400 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1477.665 1490.985 1477.835 1538.755 ;
        RECT 1478.125 1466.165 1478.295 1490.475 ;
        RECT 1477.205 1317.245 1477.375 1369.775 ;
        RECT 1477.665 1256.045 1477.835 1304.155 ;
        RECT 1477.665 1013.965 1477.835 1048.815 ;
        RECT 1478.585 917.405 1478.755 1000.535 ;
        RECT 1477.665 517.565 1477.835 565.675 ;
      LAYER mcon ;
        RECT 1477.665 1538.585 1477.835 1538.755 ;
        RECT 1478.125 1490.305 1478.295 1490.475 ;
        RECT 1477.205 1369.605 1477.375 1369.775 ;
        RECT 1477.665 1303.985 1477.835 1304.155 ;
        RECT 1477.665 1048.645 1477.835 1048.815 ;
        RECT 1478.585 1000.365 1478.755 1000.535 ;
        RECT 1477.665 565.505 1477.835 565.675 ;
      LAYER met1 ;
        RECT 1478.970 1656.380 1479.290 1656.440 ;
        RECT 1478.140 1656.240 1479.290 1656.380 ;
        RECT 1478.140 1656.100 1478.280 1656.240 ;
        RECT 1478.970 1656.180 1479.290 1656.240 ;
        RECT 1478.050 1655.840 1478.370 1656.100 ;
        RECT 1477.590 1538.740 1477.910 1538.800 ;
        RECT 1477.395 1538.600 1477.910 1538.740 ;
        RECT 1477.590 1538.540 1477.910 1538.600 ;
        RECT 1477.605 1491.140 1477.895 1491.185 ;
        RECT 1477.605 1491.000 1478.280 1491.140 ;
        RECT 1477.605 1490.955 1477.895 1491.000 ;
        RECT 1478.140 1490.505 1478.280 1491.000 ;
        RECT 1478.065 1490.275 1478.355 1490.505 ;
        RECT 1478.065 1466.320 1478.355 1466.365 ;
        RECT 1478.510 1466.320 1478.830 1466.380 ;
        RECT 1478.065 1466.180 1478.830 1466.320 ;
        RECT 1478.065 1466.135 1478.355 1466.180 ;
        RECT 1478.510 1466.120 1478.830 1466.180 ;
        RECT 1477.130 1400.700 1477.450 1400.760 ;
        RECT 1478.510 1400.700 1478.830 1400.760 ;
        RECT 1477.130 1400.560 1478.830 1400.700 ;
        RECT 1477.130 1400.500 1477.450 1400.560 ;
        RECT 1478.510 1400.500 1478.830 1400.560 ;
        RECT 1477.130 1369.760 1477.450 1369.820 ;
        RECT 1476.935 1369.620 1477.450 1369.760 ;
        RECT 1477.130 1369.560 1477.450 1369.620 ;
        RECT 1477.145 1317.400 1477.435 1317.445 ;
        RECT 1478.050 1317.400 1478.370 1317.460 ;
        RECT 1477.145 1317.260 1478.370 1317.400 ;
        RECT 1477.145 1317.215 1477.435 1317.260 ;
        RECT 1478.050 1317.200 1478.370 1317.260 ;
        RECT 1477.605 1304.140 1477.895 1304.185 ;
        RECT 1478.050 1304.140 1478.370 1304.200 ;
        RECT 1477.605 1304.000 1478.370 1304.140 ;
        RECT 1477.605 1303.955 1477.895 1304.000 ;
        RECT 1478.050 1303.940 1478.370 1304.000 ;
        RECT 1477.590 1256.200 1477.910 1256.260 ;
        RECT 1477.395 1256.060 1477.910 1256.200 ;
        RECT 1477.590 1256.000 1477.910 1256.060 ;
        RECT 1478.510 1207.580 1478.830 1207.640 ;
        RECT 1478.970 1207.580 1479.290 1207.640 ;
        RECT 1478.510 1207.440 1479.290 1207.580 ;
        RECT 1478.510 1207.380 1478.830 1207.440 ;
        RECT 1478.970 1207.380 1479.290 1207.440 ;
        RECT 1477.590 1159.300 1477.910 1159.360 ;
        RECT 1478.970 1159.300 1479.290 1159.360 ;
        RECT 1477.590 1159.160 1479.290 1159.300 ;
        RECT 1477.590 1159.100 1477.910 1159.160 ;
        RECT 1478.970 1159.100 1479.290 1159.160 ;
        RECT 1477.590 1111.020 1477.910 1111.080 ;
        RECT 1478.970 1111.020 1479.290 1111.080 ;
        RECT 1477.590 1110.880 1479.290 1111.020 ;
        RECT 1477.590 1110.820 1477.910 1110.880 ;
        RECT 1478.970 1110.820 1479.290 1110.880 ;
        RECT 1477.590 1048.800 1477.910 1048.860 ;
        RECT 1477.395 1048.660 1477.910 1048.800 ;
        RECT 1477.590 1048.600 1477.910 1048.660 ;
        RECT 1477.590 1014.120 1477.910 1014.180 ;
        RECT 1477.395 1013.980 1477.910 1014.120 ;
        RECT 1477.590 1013.920 1477.910 1013.980 ;
        RECT 1477.590 1000.520 1477.910 1000.580 ;
        RECT 1478.525 1000.520 1478.815 1000.565 ;
        RECT 1477.590 1000.380 1478.815 1000.520 ;
        RECT 1477.590 1000.320 1477.910 1000.380 ;
        RECT 1478.525 1000.335 1478.815 1000.380 ;
        RECT 1478.510 917.560 1478.830 917.620 ;
        RECT 1478.315 917.420 1478.830 917.560 ;
        RECT 1478.510 917.360 1478.830 917.420 ;
        RECT 1478.050 862.820 1478.370 862.880 ;
        RECT 1478.510 862.820 1478.830 862.880 ;
        RECT 1478.050 862.680 1478.830 862.820 ;
        RECT 1478.050 862.620 1478.370 862.680 ;
        RECT 1478.510 862.620 1478.830 862.680 ;
        RECT 1478.050 724.440 1478.370 724.500 ;
        RECT 1478.510 724.440 1478.830 724.500 ;
        RECT 1478.050 724.300 1478.830 724.440 ;
        RECT 1478.050 724.240 1478.370 724.300 ;
        RECT 1478.510 724.240 1478.830 724.300 ;
        RECT 1477.590 620.740 1477.910 620.800 ;
        RECT 1478.050 620.740 1478.370 620.800 ;
        RECT 1477.590 620.600 1478.370 620.740 ;
        RECT 1477.590 620.540 1477.910 620.600 ;
        RECT 1478.050 620.540 1478.370 620.600 ;
        RECT 1477.590 565.660 1477.910 565.720 ;
        RECT 1477.395 565.520 1477.910 565.660 ;
        RECT 1477.590 565.460 1477.910 565.520 ;
        RECT 1477.590 517.720 1477.910 517.780 ;
        RECT 1477.395 517.580 1477.910 517.720 ;
        RECT 1477.590 517.520 1477.910 517.580 ;
        RECT 1477.590 476.040 1477.910 476.300 ;
        RECT 1477.680 475.560 1477.820 476.040 ;
        RECT 1478.050 475.560 1478.370 475.620 ;
        RECT 1477.680 475.420 1478.370 475.560 ;
        RECT 1478.050 475.360 1478.370 475.420 ;
        RECT 1477.590 427.960 1477.910 428.020 ;
        RECT 1478.050 427.960 1478.370 428.020 ;
        RECT 1477.590 427.820 1478.370 427.960 ;
        RECT 1477.590 427.760 1477.910 427.820 ;
        RECT 1478.050 427.760 1478.370 427.820 ;
        RECT 1477.590 186.560 1477.910 186.620 ;
        RECT 1478.510 186.560 1478.830 186.620 ;
        RECT 1477.590 186.420 1478.830 186.560 ;
        RECT 1477.590 186.360 1477.910 186.420 ;
        RECT 1478.510 186.360 1478.830 186.420 ;
        RECT 648.210 75.720 648.530 75.780 ;
        RECT 1477.590 75.720 1477.910 75.780 ;
        RECT 648.210 75.580 1477.910 75.720 ;
        RECT 648.210 75.520 648.530 75.580 ;
        RECT 1477.590 75.520 1477.910 75.580 ;
      LAYER via ;
        RECT 1479.000 1656.180 1479.260 1656.440 ;
        RECT 1478.080 1655.840 1478.340 1656.100 ;
        RECT 1477.620 1538.540 1477.880 1538.800 ;
        RECT 1478.540 1466.120 1478.800 1466.380 ;
        RECT 1477.160 1400.500 1477.420 1400.760 ;
        RECT 1478.540 1400.500 1478.800 1400.760 ;
        RECT 1477.160 1369.560 1477.420 1369.820 ;
        RECT 1478.080 1317.200 1478.340 1317.460 ;
        RECT 1478.080 1303.940 1478.340 1304.200 ;
        RECT 1477.620 1256.000 1477.880 1256.260 ;
        RECT 1478.540 1207.380 1478.800 1207.640 ;
        RECT 1479.000 1207.380 1479.260 1207.640 ;
        RECT 1477.620 1159.100 1477.880 1159.360 ;
        RECT 1479.000 1159.100 1479.260 1159.360 ;
        RECT 1477.620 1110.820 1477.880 1111.080 ;
        RECT 1479.000 1110.820 1479.260 1111.080 ;
        RECT 1477.620 1048.600 1477.880 1048.860 ;
        RECT 1477.620 1013.920 1477.880 1014.180 ;
        RECT 1477.620 1000.320 1477.880 1000.580 ;
        RECT 1478.540 917.360 1478.800 917.620 ;
        RECT 1478.080 862.620 1478.340 862.880 ;
        RECT 1478.540 862.620 1478.800 862.880 ;
        RECT 1478.080 724.240 1478.340 724.500 ;
        RECT 1478.540 724.240 1478.800 724.500 ;
        RECT 1477.620 620.540 1477.880 620.800 ;
        RECT 1478.080 620.540 1478.340 620.800 ;
        RECT 1477.620 565.460 1477.880 565.720 ;
        RECT 1477.620 517.520 1477.880 517.780 ;
        RECT 1477.620 476.040 1477.880 476.300 ;
        RECT 1478.080 475.360 1478.340 475.620 ;
        RECT 1477.620 427.760 1477.880 428.020 ;
        RECT 1478.080 427.760 1478.340 428.020 ;
        RECT 1477.620 186.360 1477.880 186.620 ;
        RECT 1478.540 186.360 1478.800 186.620 ;
        RECT 648.240 75.520 648.500 75.780 ;
        RECT 1477.620 75.520 1477.880 75.780 ;
      LAYER met2 ;
        RECT 1480.300 1700.410 1480.580 1704.000 ;
        RECT 1479.060 1700.270 1480.580 1700.410 ;
        RECT 1479.060 1656.470 1479.200 1700.270 ;
        RECT 1480.300 1700.000 1480.580 1700.270 ;
        RECT 1479.000 1656.150 1479.260 1656.470 ;
        RECT 1478.080 1655.810 1478.340 1656.130 ;
        RECT 1478.140 1559.650 1478.280 1655.810 ;
        RECT 1477.680 1559.510 1478.280 1559.650 ;
        RECT 1477.680 1538.830 1477.820 1559.510 ;
        RECT 1477.620 1538.510 1477.880 1538.830 ;
        RECT 1478.540 1466.090 1478.800 1466.410 ;
        RECT 1478.600 1400.790 1478.740 1466.090 ;
        RECT 1477.160 1400.470 1477.420 1400.790 ;
        RECT 1478.540 1400.470 1478.800 1400.790 ;
        RECT 1477.220 1369.850 1477.360 1400.470 ;
        RECT 1477.160 1369.530 1477.420 1369.850 ;
        RECT 1478.080 1317.170 1478.340 1317.490 ;
        RECT 1478.140 1304.230 1478.280 1317.170 ;
        RECT 1478.080 1303.910 1478.340 1304.230 ;
        RECT 1477.620 1255.970 1477.880 1256.290 ;
        RECT 1477.680 1231.890 1477.820 1255.970 ;
        RECT 1477.680 1231.750 1478.740 1231.890 ;
        RECT 1478.600 1207.670 1478.740 1231.750 ;
        RECT 1478.540 1207.350 1478.800 1207.670 ;
        RECT 1479.000 1207.350 1479.260 1207.670 ;
        RECT 1479.060 1159.390 1479.200 1207.350 ;
        RECT 1477.620 1159.070 1477.880 1159.390 ;
        RECT 1479.000 1159.070 1479.260 1159.390 ;
        RECT 1477.680 1111.110 1477.820 1159.070 ;
        RECT 1477.620 1110.790 1477.880 1111.110 ;
        RECT 1479.000 1110.790 1479.260 1111.110 ;
        RECT 1479.060 1080.250 1479.200 1110.790 ;
        RECT 1477.680 1080.110 1479.200 1080.250 ;
        RECT 1477.680 1048.890 1477.820 1080.110 ;
        RECT 1477.620 1048.570 1477.880 1048.890 ;
        RECT 1477.620 1013.890 1477.880 1014.210 ;
        RECT 1477.680 1000.610 1477.820 1013.890 ;
        RECT 1477.620 1000.290 1477.880 1000.610 ;
        RECT 1478.540 917.330 1478.800 917.650 ;
        RECT 1478.600 862.910 1478.740 917.330 ;
        RECT 1478.080 862.590 1478.340 862.910 ;
        RECT 1478.540 862.590 1478.800 862.910 ;
        RECT 1478.140 787.170 1478.280 862.590 ;
        RECT 1478.140 787.030 1478.740 787.170 ;
        RECT 1478.600 766.090 1478.740 787.030 ;
        RECT 1478.140 765.950 1478.740 766.090 ;
        RECT 1478.140 724.530 1478.280 765.950 ;
        RECT 1478.080 724.210 1478.340 724.530 ;
        RECT 1478.540 724.210 1478.800 724.530 ;
        RECT 1478.600 676.445 1478.740 724.210 ;
        RECT 1477.610 676.075 1477.890 676.445 ;
        RECT 1478.530 676.075 1478.810 676.445 ;
        RECT 1477.680 645.050 1477.820 676.075 ;
        RECT 1477.220 644.910 1477.820 645.050 ;
        RECT 1477.220 626.690 1477.360 644.910 ;
        RECT 1477.220 626.550 1478.280 626.690 ;
        RECT 1478.140 620.830 1478.280 626.550 ;
        RECT 1477.620 620.510 1477.880 620.830 ;
        RECT 1478.080 620.510 1478.340 620.830 ;
        RECT 1477.680 567.530 1477.820 620.510 ;
        RECT 1477.680 567.390 1478.280 567.530 ;
        RECT 1478.140 566.170 1478.280 567.390 ;
        RECT 1477.680 566.030 1478.280 566.170 ;
        RECT 1477.680 565.750 1477.820 566.030 ;
        RECT 1477.620 565.430 1477.880 565.750 ;
        RECT 1477.620 517.490 1477.880 517.810 ;
        RECT 1477.680 476.330 1477.820 517.490 ;
        RECT 1477.620 476.010 1477.880 476.330 ;
        RECT 1478.080 475.330 1478.340 475.650 ;
        RECT 1478.140 428.050 1478.280 475.330 ;
        RECT 1477.620 427.730 1477.880 428.050 ;
        RECT 1478.080 427.730 1478.340 428.050 ;
        RECT 1477.680 282.610 1477.820 427.730 ;
        RECT 1477.680 282.470 1478.740 282.610 ;
        RECT 1478.600 186.650 1478.740 282.470 ;
        RECT 1477.620 186.330 1477.880 186.650 ;
        RECT 1478.540 186.330 1478.800 186.650 ;
        RECT 1477.680 75.810 1477.820 186.330 ;
        RECT 648.240 75.490 648.500 75.810 ;
        RECT 1477.620 75.490 1477.880 75.810 ;
        RECT 648.300 17.410 648.440 75.490 ;
        RECT 645.080 17.270 648.440 17.410 ;
        RECT 645.080 2.400 645.220 17.270 ;
        RECT 644.870 -4.800 645.430 2.400 ;
      LAYER via2 ;
        RECT 1477.610 676.120 1477.890 676.400 ;
        RECT 1478.530 676.120 1478.810 676.400 ;
      LAYER met3 ;
        RECT 1477.585 676.410 1477.915 676.425 ;
        RECT 1478.505 676.410 1478.835 676.425 ;
        RECT 1477.585 676.110 1478.835 676.410 ;
        RECT 1477.585 676.095 1477.915 676.110 ;
        RECT 1478.505 676.095 1478.835 676.110 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2398.970 1687.660 2399.290 1687.720 ;
        RECT 2429.790 1687.660 2430.110 1687.720 ;
        RECT 2398.970 1687.520 2430.110 1687.660 ;
        RECT 2398.970 1687.460 2399.290 1687.520 ;
        RECT 2429.790 1687.460 2430.110 1687.520 ;
      LAYER via ;
        RECT 2399.000 1687.460 2399.260 1687.720 ;
        RECT 2429.820 1687.460 2430.080 1687.720 ;
      LAYER met2 ;
        RECT 2398.920 1700.000 2399.200 1704.000 ;
        RECT 2399.060 1687.750 2399.200 1700.000 ;
        RECT 2399.000 1687.430 2399.260 1687.750 ;
        RECT 2429.820 1687.430 2430.080 1687.750 ;
        RECT 2429.880 3.130 2430.020 1687.430 ;
        RECT 2428.960 2.990 2430.020 3.130 ;
        RECT 2428.960 2.400 2429.100 2.990 ;
        RECT 2428.750 -4.800 2429.310 2.400 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2408.170 1683.920 2408.490 1683.980 ;
        RECT 2414.610 1683.920 2414.930 1683.980 ;
        RECT 2408.170 1683.780 2414.930 1683.920 ;
        RECT 2408.170 1683.720 2408.490 1683.780 ;
        RECT 2414.610 1683.720 2414.930 1683.780 ;
        RECT 2414.610 16.900 2414.930 16.960 ;
        RECT 2446.810 16.900 2447.130 16.960 ;
        RECT 2414.610 16.760 2447.130 16.900 ;
        RECT 2414.610 16.700 2414.930 16.760 ;
        RECT 2446.810 16.700 2447.130 16.760 ;
      LAYER via ;
        RECT 2408.200 1683.720 2408.460 1683.980 ;
        RECT 2414.640 1683.720 2414.900 1683.980 ;
        RECT 2414.640 16.700 2414.900 16.960 ;
        RECT 2446.840 16.700 2447.100 16.960 ;
      LAYER met2 ;
        RECT 2408.120 1700.000 2408.400 1704.000 ;
        RECT 2408.260 1684.010 2408.400 1700.000 ;
        RECT 2408.200 1683.690 2408.460 1684.010 ;
        RECT 2414.640 1683.690 2414.900 1684.010 ;
        RECT 2414.700 16.990 2414.840 1683.690 ;
        RECT 2414.640 16.670 2414.900 16.990 ;
        RECT 2446.840 16.670 2447.100 16.990 ;
        RECT 2446.900 2.400 2447.040 16.670 ;
        RECT 2446.690 -4.800 2447.250 2.400 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2417.370 1683.920 2417.690 1683.980 ;
        RECT 2421.510 1683.920 2421.830 1683.980 ;
        RECT 2417.370 1683.780 2421.830 1683.920 ;
        RECT 2417.370 1683.720 2417.690 1683.780 ;
        RECT 2421.510 1683.720 2421.830 1683.780 ;
        RECT 2421.510 18.260 2421.830 18.320 ;
        RECT 2464.750 18.260 2465.070 18.320 ;
        RECT 2421.510 18.120 2465.070 18.260 ;
        RECT 2421.510 18.060 2421.830 18.120 ;
        RECT 2464.750 18.060 2465.070 18.120 ;
      LAYER via ;
        RECT 2417.400 1683.720 2417.660 1683.980 ;
        RECT 2421.540 1683.720 2421.800 1683.980 ;
        RECT 2421.540 18.060 2421.800 18.320 ;
        RECT 2464.780 18.060 2465.040 18.320 ;
      LAYER met2 ;
        RECT 2417.320 1700.000 2417.600 1704.000 ;
        RECT 2417.460 1684.010 2417.600 1700.000 ;
        RECT 2417.400 1683.690 2417.660 1684.010 ;
        RECT 2421.540 1683.690 2421.800 1684.010 ;
        RECT 2421.600 18.350 2421.740 1683.690 ;
        RECT 2421.540 18.030 2421.800 18.350 ;
        RECT 2464.780 18.030 2465.040 18.350 ;
        RECT 2464.840 2.400 2464.980 18.030 ;
        RECT 2464.630 -4.800 2465.190 2.400 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2426.570 1687.320 2426.890 1687.380 ;
        RECT 2466.590 1687.320 2466.910 1687.380 ;
        RECT 2426.570 1687.180 2466.910 1687.320 ;
        RECT 2426.570 1687.120 2426.890 1687.180 ;
        RECT 2466.590 1687.120 2466.910 1687.180 ;
        RECT 2466.590 15.880 2466.910 15.940 ;
        RECT 2482.690 15.880 2483.010 15.940 ;
        RECT 2466.590 15.740 2483.010 15.880 ;
        RECT 2466.590 15.680 2466.910 15.740 ;
        RECT 2482.690 15.680 2483.010 15.740 ;
      LAYER via ;
        RECT 2426.600 1687.120 2426.860 1687.380 ;
        RECT 2466.620 1687.120 2466.880 1687.380 ;
        RECT 2466.620 15.680 2466.880 15.940 ;
        RECT 2482.720 15.680 2482.980 15.940 ;
      LAYER met2 ;
        RECT 2426.520 1700.000 2426.800 1704.000 ;
        RECT 2426.660 1687.410 2426.800 1700.000 ;
        RECT 2426.600 1687.090 2426.860 1687.410 ;
        RECT 2466.620 1687.090 2466.880 1687.410 ;
        RECT 2466.680 15.970 2466.820 1687.090 ;
        RECT 2466.620 15.650 2466.880 15.970 ;
        RECT 2482.720 15.650 2482.980 15.970 ;
        RECT 2482.780 2.400 2482.920 15.650 ;
        RECT 2482.570 -4.800 2483.130 2.400 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2435.770 1688.680 2436.090 1688.740 ;
        RECT 2498.790 1688.680 2499.110 1688.740 ;
        RECT 2435.770 1688.540 2499.110 1688.680 ;
        RECT 2435.770 1688.480 2436.090 1688.540 ;
        RECT 2498.790 1688.480 2499.110 1688.540 ;
        RECT 2498.790 2.960 2499.110 3.020 ;
        RECT 2500.630 2.960 2500.950 3.020 ;
        RECT 2498.790 2.820 2500.950 2.960 ;
        RECT 2498.790 2.760 2499.110 2.820 ;
        RECT 2500.630 2.760 2500.950 2.820 ;
      LAYER via ;
        RECT 2435.800 1688.480 2436.060 1688.740 ;
        RECT 2498.820 1688.480 2499.080 1688.740 ;
        RECT 2498.820 2.760 2499.080 3.020 ;
        RECT 2500.660 2.760 2500.920 3.020 ;
      LAYER met2 ;
        RECT 2435.720 1700.000 2436.000 1704.000 ;
        RECT 2435.860 1688.770 2436.000 1700.000 ;
        RECT 2435.800 1688.450 2436.060 1688.770 ;
        RECT 2498.820 1688.450 2499.080 1688.770 ;
        RECT 2498.880 3.050 2499.020 1688.450 ;
        RECT 2498.820 2.730 2499.080 3.050 ;
        RECT 2500.660 2.730 2500.920 3.050 ;
        RECT 2500.720 2.400 2500.860 2.730 ;
        RECT 2500.510 -4.800 2501.070 2.400 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2444.970 1689.020 2445.290 1689.080 ;
        RECT 2513.050 1689.020 2513.370 1689.080 ;
        RECT 2444.970 1688.880 2513.370 1689.020 ;
        RECT 2444.970 1688.820 2445.290 1688.880 ;
        RECT 2513.050 1688.820 2513.370 1688.880 ;
      LAYER via ;
        RECT 2445.000 1688.820 2445.260 1689.080 ;
        RECT 2513.080 1688.820 2513.340 1689.080 ;
      LAYER met2 ;
        RECT 2444.920 1700.000 2445.200 1704.000 ;
        RECT 2445.060 1689.110 2445.200 1700.000 ;
        RECT 2445.000 1688.790 2445.260 1689.110 ;
        RECT 2513.080 1688.790 2513.340 1689.110 ;
        RECT 2513.140 16.730 2513.280 1688.790 ;
        RECT 2513.140 16.590 2518.340 16.730 ;
        RECT 2518.200 2.400 2518.340 16.590 ;
        RECT 2517.990 -4.800 2518.550 2.400 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2495.185 1687.845 2495.355 1690.055 ;
        RECT 2511.745 1686.485 2511.915 1688.015 ;
      LAYER mcon ;
        RECT 2495.185 1689.885 2495.355 1690.055 ;
        RECT 2511.745 1687.845 2511.915 1688.015 ;
      LAYER met1 ;
        RECT 2454.170 1690.040 2454.490 1690.100 ;
        RECT 2495.125 1690.040 2495.415 1690.085 ;
        RECT 2454.170 1689.900 2495.415 1690.040 ;
        RECT 2454.170 1689.840 2454.490 1689.900 ;
        RECT 2495.125 1689.855 2495.415 1689.900 ;
        RECT 2495.125 1688.000 2495.415 1688.045 ;
        RECT 2511.685 1688.000 2511.975 1688.045 ;
        RECT 2495.125 1687.860 2511.975 1688.000 ;
        RECT 2495.125 1687.815 2495.415 1687.860 ;
        RECT 2511.685 1687.815 2511.975 1687.860 ;
        RECT 2511.685 1686.640 2511.975 1686.685 ;
        RECT 2533.290 1686.640 2533.610 1686.700 ;
        RECT 2511.685 1686.500 2533.610 1686.640 ;
        RECT 2511.685 1686.455 2511.975 1686.500 ;
        RECT 2533.290 1686.440 2533.610 1686.500 ;
        RECT 2533.290 2.960 2533.610 3.020 ;
        RECT 2536.050 2.960 2536.370 3.020 ;
        RECT 2533.290 2.820 2536.370 2.960 ;
        RECT 2533.290 2.760 2533.610 2.820 ;
        RECT 2536.050 2.760 2536.370 2.820 ;
      LAYER via ;
        RECT 2454.200 1689.840 2454.460 1690.100 ;
        RECT 2533.320 1686.440 2533.580 1686.700 ;
        RECT 2533.320 2.760 2533.580 3.020 ;
        RECT 2536.080 2.760 2536.340 3.020 ;
      LAYER met2 ;
        RECT 2454.120 1700.000 2454.400 1704.000 ;
        RECT 2454.260 1690.130 2454.400 1700.000 ;
        RECT 2454.200 1689.810 2454.460 1690.130 ;
        RECT 2533.320 1686.410 2533.580 1686.730 ;
        RECT 2533.380 3.050 2533.520 1686.410 ;
        RECT 2533.320 2.730 2533.580 3.050 ;
        RECT 2536.080 2.730 2536.340 3.050 ;
        RECT 2536.140 2.400 2536.280 2.730 ;
        RECT 2535.930 -4.800 2536.490 2.400 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2553.990 1688.340 2554.310 1688.400 ;
        RECT 2494.740 1688.200 2554.310 1688.340 ;
        RECT 2463.370 1688.000 2463.690 1688.060 ;
        RECT 2494.740 1688.000 2494.880 1688.200 ;
        RECT 2553.990 1688.140 2554.310 1688.200 ;
        RECT 2463.370 1687.860 2494.880 1688.000 ;
        RECT 2463.370 1687.800 2463.690 1687.860 ;
      LAYER via ;
        RECT 2463.400 1687.800 2463.660 1688.060 ;
        RECT 2554.020 1688.140 2554.280 1688.400 ;
      LAYER met2 ;
        RECT 2463.320 1700.000 2463.600 1704.000 ;
        RECT 2463.460 1688.090 2463.600 1700.000 ;
        RECT 2554.020 1688.110 2554.280 1688.430 ;
        RECT 2463.400 1687.770 2463.660 1688.090 ;
        RECT 2554.080 2.400 2554.220 1688.110 ;
        RECT 2553.870 -4.800 2554.430 2.400 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2472.570 1687.660 2472.890 1687.720 ;
        RECT 2567.790 1687.660 2568.110 1687.720 ;
        RECT 2472.570 1687.520 2568.110 1687.660 ;
        RECT 2472.570 1687.460 2472.890 1687.520 ;
        RECT 2567.790 1687.460 2568.110 1687.520 ;
        RECT 2567.790 2.960 2568.110 3.020 ;
        RECT 2571.930 2.960 2572.250 3.020 ;
        RECT 2567.790 2.820 2572.250 2.960 ;
        RECT 2567.790 2.760 2568.110 2.820 ;
        RECT 2571.930 2.760 2572.250 2.820 ;
      LAYER via ;
        RECT 2472.600 1687.460 2472.860 1687.720 ;
        RECT 2567.820 1687.460 2568.080 1687.720 ;
        RECT 2567.820 2.760 2568.080 3.020 ;
        RECT 2571.960 2.760 2572.220 3.020 ;
      LAYER met2 ;
        RECT 2472.520 1700.000 2472.800 1704.000 ;
        RECT 2472.660 1687.750 2472.800 1700.000 ;
        RECT 2472.600 1687.430 2472.860 1687.750 ;
        RECT 2567.820 1687.430 2568.080 1687.750 ;
        RECT 2567.880 3.050 2568.020 1687.430 ;
        RECT 2567.820 2.730 2568.080 3.050 ;
        RECT 2571.960 2.730 2572.220 3.050 ;
        RECT 2572.020 2.400 2572.160 2.730 ;
        RECT 2571.810 -4.800 2572.370 2.400 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2481.310 1687.320 2481.630 1687.380 ;
        RECT 2481.310 1687.180 2554.680 1687.320 ;
        RECT 2481.310 1687.120 2481.630 1687.180 ;
        RECT 2554.540 1686.980 2554.680 1687.180 ;
        RECT 2588.030 1686.980 2588.350 1687.040 ;
        RECT 2554.540 1686.840 2588.350 1686.980 ;
        RECT 2588.030 1686.780 2588.350 1686.840 ;
      LAYER via ;
        RECT 2481.340 1687.120 2481.600 1687.380 ;
        RECT 2588.060 1686.780 2588.320 1687.040 ;
      LAYER met2 ;
        RECT 2481.260 1700.000 2481.540 1704.000 ;
        RECT 2481.400 1687.410 2481.540 1700.000 ;
        RECT 2481.340 1687.090 2481.600 1687.410 ;
        RECT 2588.060 1686.750 2588.320 1687.070 ;
        RECT 2588.120 3.130 2588.260 1686.750 ;
        RECT 2588.120 2.990 2589.640 3.130 ;
        RECT 2589.500 2.400 2589.640 2.990 ;
        RECT 2589.290 -4.800 2589.850 2.400 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1567.290 1689.360 1567.610 1689.420 ;
        RECT 1570.510 1689.360 1570.830 1689.420 ;
        RECT 1567.290 1689.220 1570.830 1689.360 ;
        RECT 1567.290 1689.160 1567.610 1689.220 ;
        RECT 1570.510 1689.160 1570.830 1689.220 ;
        RECT 827.610 71.300 827.930 71.360 ;
        RECT 1567.290 71.300 1567.610 71.360 ;
        RECT 827.610 71.160 1567.610 71.300 ;
        RECT 827.610 71.100 827.930 71.160 ;
        RECT 1567.290 71.100 1567.610 71.160 ;
      LAYER via ;
        RECT 1567.320 1689.160 1567.580 1689.420 ;
        RECT 1570.540 1689.160 1570.800 1689.420 ;
        RECT 827.640 71.100 827.900 71.360 ;
        RECT 1567.320 71.100 1567.580 71.360 ;
      LAYER met2 ;
        RECT 1572.300 1700.410 1572.580 1704.000 ;
        RECT 1570.600 1700.270 1572.580 1700.410 ;
        RECT 1570.600 1689.450 1570.740 1700.270 ;
        RECT 1572.300 1700.000 1572.580 1700.270 ;
        RECT 1567.320 1689.130 1567.580 1689.450 ;
        RECT 1570.540 1689.130 1570.800 1689.450 ;
        RECT 1567.380 71.390 1567.520 1689.130 ;
        RECT 827.640 71.070 827.900 71.390 ;
        RECT 1567.320 71.070 1567.580 71.390 ;
        RECT 827.700 16.730 827.840 71.070 ;
        RECT 823.560 16.590 827.840 16.730 ;
        RECT 823.560 2.400 823.700 16.590 ;
        RECT 823.350 -4.800 823.910 2.400 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2601.830 1686.640 2602.150 1686.700 ;
        RECT 2539.360 1686.500 2602.150 1686.640 ;
        RECT 2490.510 1685.960 2490.830 1686.020 ;
        RECT 2539.360 1685.960 2539.500 1686.500 ;
        RECT 2601.830 1686.440 2602.150 1686.500 ;
        RECT 2490.510 1685.820 2539.500 1685.960 ;
        RECT 2490.510 1685.760 2490.830 1685.820 ;
        RECT 2601.830 2.960 2602.150 3.020 ;
        RECT 2607.350 2.960 2607.670 3.020 ;
        RECT 2601.830 2.820 2607.670 2.960 ;
        RECT 2601.830 2.760 2602.150 2.820 ;
        RECT 2607.350 2.760 2607.670 2.820 ;
      LAYER via ;
        RECT 2490.540 1685.760 2490.800 1686.020 ;
        RECT 2601.860 1686.440 2602.120 1686.700 ;
        RECT 2601.860 2.760 2602.120 3.020 ;
        RECT 2607.380 2.760 2607.640 3.020 ;
      LAYER met2 ;
        RECT 2490.460 1700.000 2490.740 1704.000 ;
        RECT 2490.600 1686.050 2490.740 1700.000 ;
        RECT 2601.860 1686.410 2602.120 1686.730 ;
        RECT 2490.540 1685.730 2490.800 1686.050 ;
        RECT 2601.920 3.050 2602.060 1686.410 ;
        RECT 2601.860 2.730 2602.120 3.050 ;
        RECT 2607.380 2.730 2607.640 3.050 ;
        RECT 2607.440 2.400 2607.580 2.730 ;
        RECT 2607.230 -4.800 2607.790 2.400 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2499.710 1688.680 2500.030 1688.740 ;
        RECT 2504.310 1688.680 2504.630 1688.740 ;
        RECT 2499.710 1688.540 2504.630 1688.680 ;
        RECT 2499.710 1688.480 2500.030 1688.540 ;
        RECT 2504.310 1688.480 2504.630 1688.540 ;
        RECT 2504.310 18.940 2504.630 19.000 ;
        RECT 2625.290 18.940 2625.610 19.000 ;
        RECT 2504.310 18.800 2625.610 18.940 ;
        RECT 2504.310 18.740 2504.630 18.800 ;
        RECT 2625.290 18.740 2625.610 18.800 ;
      LAYER via ;
        RECT 2499.740 1688.480 2500.000 1688.740 ;
        RECT 2504.340 1688.480 2504.600 1688.740 ;
        RECT 2504.340 18.740 2504.600 19.000 ;
        RECT 2625.320 18.740 2625.580 19.000 ;
      LAYER met2 ;
        RECT 2499.660 1700.000 2499.940 1704.000 ;
        RECT 2499.800 1688.770 2499.940 1700.000 ;
        RECT 2499.740 1688.450 2500.000 1688.770 ;
        RECT 2504.340 1688.450 2504.600 1688.770 ;
        RECT 2504.400 19.030 2504.540 1688.450 ;
        RECT 2504.340 18.710 2504.600 19.030 ;
        RECT 2625.320 18.710 2625.580 19.030 ;
        RECT 2625.380 2.400 2625.520 18.710 ;
        RECT 2625.170 -4.800 2625.730 2.400 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2511.210 17.240 2511.530 17.300 ;
        RECT 2643.230 17.240 2643.550 17.300 ;
        RECT 2511.210 17.100 2643.550 17.240 ;
        RECT 2511.210 17.040 2511.530 17.100 ;
        RECT 2643.230 17.040 2643.550 17.100 ;
      LAYER via ;
        RECT 2511.240 17.040 2511.500 17.300 ;
        RECT 2643.260 17.040 2643.520 17.300 ;
      LAYER met2 ;
        RECT 2508.860 1700.410 2509.140 1704.000 ;
        RECT 2508.860 1700.270 2511.440 1700.410 ;
        RECT 2508.860 1700.000 2509.140 1700.270 ;
        RECT 2511.300 17.330 2511.440 1700.270 ;
        RECT 2511.240 17.010 2511.500 17.330 ;
        RECT 2643.260 17.010 2643.520 17.330 ;
        RECT 2643.320 2.400 2643.460 17.010 ;
        RECT 2643.110 -4.800 2643.670 2.400 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2622.145 1683.765 2622.315 1686.995 ;
      LAYER mcon ;
        RECT 2622.145 1686.825 2622.315 1686.995 ;
      LAYER met1 ;
        RECT 2517.190 1689.700 2517.510 1689.760 ;
        RECT 2518.110 1689.700 2518.430 1689.760 ;
        RECT 2517.190 1689.560 2518.430 1689.700 ;
        RECT 2517.190 1689.500 2517.510 1689.560 ;
        RECT 2518.110 1689.500 2518.430 1689.560 ;
        RECT 2622.085 1686.980 2622.375 1687.025 ;
        RECT 2656.570 1686.980 2656.890 1687.040 ;
        RECT 2622.085 1686.840 2656.890 1686.980 ;
        RECT 2622.085 1686.795 2622.375 1686.840 ;
        RECT 2656.570 1686.780 2656.890 1686.840 ;
        RECT 2517.190 1683.920 2517.510 1683.980 ;
        RECT 2622.085 1683.920 2622.375 1683.965 ;
        RECT 2517.190 1683.780 2622.375 1683.920 ;
        RECT 2517.190 1683.720 2517.510 1683.780 ;
        RECT 2622.085 1683.735 2622.375 1683.780 ;
      LAYER via ;
        RECT 2517.220 1689.500 2517.480 1689.760 ;
        RECT 2518.140 1689.500 2518.400 1689.760 ;
        RECT 2656.600 1686.780 2656.860 1687.040 ;
        RECT 2517.220 1683.720 2517.480 1683.980 ;
      LAYER met2 ;
        RECT 2518.060 1700.000 2518.340 1704.000 ;
        RECT 2518.200 1689.790 2518.340 1700.000 ;
        RECT 2517.220 1689.470 2517.480 1689.790 ;
        RECT 2518.140 1689.470 2518.400 1689.790 ;
        RECT 2517.280 1684.010 2517.420 1689.470 ;
        RECT 2656.600 1686.750 2656.860 1687.070 ;
        RECT 2517.220 1683.690 2517.480 1684.010 ;
        RECT 2656.660 16.730 2656.800 1686.750 ;
        RECT 2656.660 16.590 2661.400 16.730 ;
        RECT 2661.260 2.400 2661.400 16.590 ;
        RECT 2661.050 -4.800 2661.610 2.400 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2527.310 1688.680 2527.630 1688.740 ;
        RECT 2531.910 1688.680 2532.230 1688.740 ;
        RECT 2527.310 1688.540 2532.230 1688.680 ;
        RECT 2527.310 1688.480 2527.630 1688.540 ;
        RECT 2531.910 1688.480 2532.230 1688.540 ;
        RECT 2531.910 15.200 2532.230 15.260 ;
        RECT 2678.650 15.200 2678.970 15.260 ;
        RECT 2531.910 15.060 2678.970 15.200 ;
        RECT 2531.910 15.000 2532.230 15.060 ;
        RECT 2678.650 15.000 2678.970 15.060 ;
      LAYER via ;
        RECT 2527.340 1688.480 2527.600 1688.740 ;
        RECT 2531.940 1688.480 2532.200 1688.740 ;
        RECT 2531.940 15.000 2532.200 15.260 ;
        RECT 2678.680 15.000 2678.940 15.260 ;
      LAYER met2 ;
        RECT 2527.260 1700.000 2527.540 1704.000 ;
        RECT 2527.400 1688.770 2527.540 1700.000 ;
        RECT 2527.340 1688.450 2527.600 1688.770 ;
        RECT 2531.940 1688.450 2532.200 1688.770 ;
        RECT 2532.000 15.290 2532.140 1688.450 ;
        RECT 2531.940 14.970 2532.200 15.290 ;
        RECT 2678.680 14.970 2678.940 15.290 ;
        RECT 2678.740 2.400 2678.880 14.970 ;
        RECT 2678.530 -4.800 2679.090 2.400 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2536.510 1685.620 2536.830 1685.680 ;
        RECT 2691.070 1685.620 2691.390 1685.680 ;
        RECT 2536.510 1685.480 2691.390 1685.620 ;
        RECT 2536.510 1685.420 2536.830 1685.480 ;
        RECT 2691.070 1685.420 2691.390 1685.480 ;
      LAYER via ;
        RECT 2536.540 1685.420 2536.800 1685.680 ;
        RECT 2691.100 1685.420 2691.360 1685.680 ;
      LAYER met2 ;
        RECT 2536.460 1700.000 2536.740 1704.000 ;
        RECT 2536.600 1685.710 2536.740 1700.000 ;
        RECT 2536.540 1685.390 2536.800 1685.710 ;
        RECT 2691.100 1685.390 2691.360 1685.710 ;
        RECT 2691.160 16.730 2691.300 1685.390 ;
        RECT 2691.160 16.590 2696.820 16.730 ;
        RECT 2696.680 2.400 2696.820 16.590 ;
        RECT 2696.470 -4.800 2697.030 2.400 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2545.250 1685.960 2545.570 1686.020 ;
        RECT 2701.190 1685.960 2701.510 1686.020 ;
        RECT 2545.250 1685.820 2701.510 1685.960 ;
        RECT 2545.250 1685.760 2545.570 1685.820 ;
        RECT 2701.190 1685.760 2701.510 1685.820 ;
        RECT 2701.190 16.560 2701.510 16.620 ;
        RECT 2714.530 16.560 2714.850 16.620 ;
        RECT 2701.190 16.420 2714.850 16.560 ;
        RECT 2701.190 16.360 2701.510 16.420 ;
        RECT 2714.530 16.360 2714.850 16.420 ;
      LAYER via ;
        RECT 2545.280 1685.760 2545.540 1686.020 ;
        RECT 2701.220 1685.760 2701.480 1686.020 ;
        RECT 2701.220 16.360 2701.480 16.620 ;
        RECT 2714.560 16.360 2714.820 16.620 ;
      LAYER met2 ;
        RECT 2545.660 1700.410 2545.940 1704.000 ;
        RECT 2545.340 1700.270 2545.940 1700.410 ;
        RECT 2545.340 1686.050 2545.480 1700.270 ;
        RECT 2545.660 1700.000 2545.940 1700.270 ;
        RECT 2545.280 1685.730 2545.540 1686.050 ;
        RECT 2701.220 1685.730 2701.480 1686.050 ;
        RECT 2701.280 16.650 2701.420 1685.730 ;
        RECT 2701.220 16.330 2701.480 16.650 ;
        RECT 2714.560 16.330 2714.820 16.650 ;
        RECT 2714.620 2.400 2714.760 16.330 ;
        RECT 2714.410 -4.800 2714.970 2.400 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2700.805 15.045 2700.975 16.575 ;
      LAYER mcon ;
        RECT 2700.805 16.405 2700.975 16.575 ;
      LAYER met1 ;
        RECT 2554.910 1687.320 2555.230 1687.380 ;
        RECT 2559.050 1687.320 2559.370 1687.380 ;
        RECT 2554.910 1687.180 2559.370 1687.320 ;
        RECT 2554.910 1687.120 2555.230 1687.180 ;
        RECT 2559.050 1687.120 2559.370 1687.180 ;
        RECT 2700.745 16.560 2701.035 16.605 ;
        RECT 2584.440 16.420 2701.035 16.560 ;
        RECT 2559.050 16.220 2559.370 16.280 ;
        RECT 2584.440 16.220 2584.580 16.420 ;
        RECT 2700.745 16.375 2701.035 16.420 ;
        RECT 2559.050 16.080 2584.580 16.220 ;
        RECT 2559.050 16.020 2559.370 16.080 ;
        RECT 2700.745 15.200 2701.035 15.245 ;
        RECT 2732.470 15.200 2732.790 15.260 ;
        RECT 2700.745 15.060 2732.790 15.200 ;
        RECT 2700.745 15.015 2701.035 15.060 ;
        RECT 2732.470 15.000 2732.790 15.060 ;
      LAYER via ;
        RECT 2554.940 1687.120 2555.200 1687.380 ;
        RECT 2559.080 1687.120 2559.340 1687.380 ;
        RECT 2559.080 16.020 2559.340 16.280 ;
        RECT 2732.500 15.000 2732.760 15.260 ;
      LAYER met2 ;
        RECT 2554.860 1700.000 2555.140 1704.000 ;
        RECT 2555.000 1687.410 2555.140 1700.000 ;
        RECT 2554.940 1687.090 2555.200 1687.410 ;
        RECT 2559.080 1687.090 2559.340 1687.410 ;
        RECT 2559.140 16.310 2559.280 1687.090 ;
        RECT 2559.080 15.990 2559.340 16.310 ;
        RECT 2732.500 14.970 2732.760 15.290 ;
        RECT 2732.560 2.400 2732.700 14.970 ;
        RECT 2732.350 -4.800 2732.910 2.400 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2564.110 1690.040 2564.430 1690.100 ;
        RECT 2736.150 1690.040 2736.470 1690.100 ;
        RECT 2564.110 1689.900 2736.470 1690.040 ;
        RECT 2564.110 1689.840 2564.430 1689.900 ;
        RECT 2736.150 1689.840 2736.470 1689.900 ;
        RECT 2736.150 16.560 2736.470 16.620 ;
        RECT 2750.410 16.560 2750.730 16.620 ;
        RECT 2736.150 16.420 2750.730 16.560 ;
        RECT 2736.150 16.360 2736.470 16.420 ;
        RECT 2750.410 16.360 2750.730 16.420 ;
      LAYER via ;
        RECT 2564.140 1689.840 2564.400 1690.100 ;
        RECT 2736.180 1689.840 2736.440 1690.100 ;
        RECT 2736.180 16.360 2736.440 16.620 ;
        RECT 2750.440 16.360 2750.700 16.620 ;
      LAYER met2 ;
        RECT 2564.060 1700.000 2564.340 1704.000 ;
        RECT 2564.200 1690.130 2564.340 1700.000 ;
        RECT 2564.140 1689.810 2564.400 1690.130 ;
        RECT 2736.180 1689.810 2736.440 1690.130 ;
        RECT 2736.240 16.650 2736.380 1689.810 ;
        RECT 2736.180 16.330 2736.440 16.650 ;
        RECT 2750.440 16.330 2750.700 16.650 ;
        RECT 2750.500 2.400 2750.640 16.330 ;
        RECT 2750.290 -4.800 2750.850 2.400 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2573.310 1689.360 2573.630 1689.420 ;
        RECT 2766.970 1689.360 2767.290 1689.420 ;
        RECT 2573.310 1689.220 2767.290 1689.360 ;
        RECT 2573.310 1689.160 2573.630 1689.220 ;
        RECT 2766.970 1689.160 2767.290 1689.220 ;
      LAYER via ;
        RECT 2573.340 1689.160 2573.600 1689.420 ;
        RECT 2767.000 1689.160 2767.260 1689.420 ;
      LAYER met2 ;
        RECT 2573.260 1700.000 2573.540 1704.000 ;
        RECT 2573.400 1689.450 2573.540 1700.000 ;
        RECT 2573.340 1689.130 2573.600 1689.450 ;
        RECT 2767.000 1689.130 2767.260 1689.450 ;
        RECT 2767.060 16.730 2767.200 1689.130 ;
        RECT 2767.060 16.590 2768.120 16.730 ;
        RECT 2767.980 2.400 2768.120 16.590 ;
        RECT 2767.770 -4.800 2768.330 2.400 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 841.410 70.960 841.730 71.020 ;
        RECT 1580.630 70.960 1580.950 71.020 ;
        RECT 841.410 70.820 1580.950 70.960 ;
        RECT 841.410 70.760 841.730 70.820 ;
        RECT 1580.630 70.760 1580.950 70.820 ;
      LAYER via ;
        RECT 841.440 70.760 841.700 71.020 ;
        RECT 1580.660 70.760 1580.920 71.020 ;
      LAYER met2 ;
        RECT 1581.500 1700.410 1581.780 1704.000 ;
        RECT 1580.720 1700.270 1581.780 1700.410 ;
        RECT 1580.720 71.050 1580.860 1700.270 ;
        RECT 1581.500 1700.000 1581.780 1700.270 ;
        RECT 841.440 70.730 841.700 71.050 ;
        RECT 1580.660 70.730 1580.920 71.050 ;
        RECT 841.500 17.410 841.640 70.730 ;
        RECT 841.040 17.270 841.640 17.410 ;
        RECT 841.040 2.400 841.180 17.270 ;
        RECT 840.830 -4.800 841.390 2.400 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2582.510 1684.940 2582.830 1685.000 ;
        RECT 2587.110 1684.940 2587.430 1685.000 ;
        RECT 2582.510 1684.800 2587.430 1684.940 ;
        RECT 2582.510 1684.740 2582.830 1684.800 ;
        RECT 2587.110 1684.740 2587.430 1684.800 ;
        RECT 2587.110 20.640 2587.430 20.700 ;
        RECT 2785.830 20.640 2786.150 20.700 ;
        RECT 2587.110 20.500 2786.150 20.640 ;
        RECT 2587.110 20.440 2587.430 20.500 ;
        RECT 2785.830 20.440 2786.150 20.500 ;
      LAYER via ;
        RECT 2582.540 1684.740 2582.800 1685.000 ;
        RECT 2587.140 1684.740 2587.400 1685.000 ;
        RECT 2587.140 20.440 2587.400 20.700 ;
        RECT 2785.860 20.440 2786.120 20.700 ;
      LAYER met2 ;
        RECT 2582.460 1700.000 2582.740 1704.000 ;
        RECT 2582.600 1685.030 2582.740 1700.000 ;
        RECT 2582.540 1684.710 2582.800 1685.030 ;
        RECT 2587.140 1684.710 2587.400 1685.030 ;
        RECT 2587.200 20.730 2587.340 1684.710 ;
        RECT 2587.140 20.410 2587.400 20.730 ;
        RECT 2785.860 20.410 2786.120 20.730 ;
        RECT 2785.920 2.400 2786.060 20.410 ;
        RECT 2785.710 -4.800 2786.270 2.400 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2591.710 1688.680 2592.030 1688.740 ;
        RECT 2801.470 1688.680 2801.790 1688.740 ;
        RECT 2591.710 1688.540 2801.790 1688.680 ;
        RECT 2591.710 1688.480 2592.030 1688.540 ;
        RECT 2801.470 1688.480 2801.790 1688.540 ;
      LAYER via ;
        RECT 2591.740 1688.480 2592.000 1688.740 ;
        RECT 2801.500 1688.480 2801.760 1688.740 ;
      LAYER met2 ;
        RECT 2591.660 1700.000 2591.940 1704.000 ;
        RECT 2591.800 1688.770 2591.940 1700.000 ;
        RECT 2591.740 1688.450 2592.000 1688.770 ;
        RECT 2801.500 1688.450 2801.760 1688.770 ;
        RECT 2801.560 17.410 2801.700 1688.450 ;
        RECT 2801.560 17.270 2804.000 17.410 ;
        RECT 2803.860 2.400 2804.000 17.270 ;
        RECT 2803.650 -4.800 2804.210 2.400 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2600.910 19.620 2601.230 19.680 ;
        RECT 2821.710 19.620 2822.030 19.680 ;
        RECT 2600.910 19.480 2822.030 19.620 ;
        RECT 2600.910 19.420 2601.230 19.480 ;
        RECT 2821.710 19.420 2822.030 19.480 ;
      LAYER via ;
        RECT 2600.940 19.420 2601.200 19.680 ;
        RECT 2821.740 19.420 2822.000 19.680 ;
      LAYER met2 ;
        RECT 2600.860 1700.000 2601.140 1704.000 ;
        RECT 2601.000 19.710 2601.140 1700.000 ;
        RECT 2600.940 19.390 2601.200 19.710 ;
        RECT 2821.740 19.390 2822.000 19.710 ;
        RECT 2821.800 2.400 2821.940 19.390 ;
        RECT 2821.590 -4.800 2822.150 2.400 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2646.525 1686.145 2646.695 1687.675 ;
      LAYER mcon ;
        RECT 2646.525 1687.505 2646.695 1687.675 ;
      LAYER met1 ;
        RECT 2646.465 1687.660 2646.755 1687.705 ;
        RECT 2835.970 1687.660 2836.290 1687.720 ;
        RECT 2646.465 1687.520 2836.290 1687.660 ;
        RECT 2646.465 1687.475 2646.755 1687.520 ;
        RECT 2835.970 1687.460 2836.290 1687.520 ;
        RECT 2610.110 1686.300 2610.430 1686.360 ;
        RECT 2646.465 1686.300 2646.755 1686.345 ;
        RECT 2610.110 1686.160 2646.755 1686.300 ;
        RECT 2610.110 1686.100 2610.430 1686.160 ;
        RECT 2646.465 1686.115 2646.755 1686.160 ;
      LAYER via ;
        RECT 2836.000 1687.460 2836.260 1687.720 ;
        RECT 2610.140 1686.100 2610.400 1686.360 ;
      LAYER met2 ;
        RECT 2610.060 1700.000 2610.340 1704.000 ;
        RECT 2610.200 1686.390 2610.340 1700.000 ;
        RECT 2836.000 1687.430 2836.260 1687.750 ;
        RECT 2610.140 1686.070 2610.400 1686.390 ;
        RECT 2836.060 16.730 2836.200 1687.430 ;
        RECT 2836.060 16.590 2839.420 16.730 ;
        RECT 2839.280 2.400 2839.420 16.590 ;
        RECT 2839.070 -4.800 2839.630 2.400 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2621.610 18.260 2621.930 18.320 ;
        RECT 2857.130 18.260 2857.450 18.320 ;
        RECT 2621.610 18.120 2857.450 18.260 ;
        RECT 2621.610 18.060 2621.930 18.120 ;
        RECT 2857.130 18.060 2857.450 18.120 ;
      LAYER via ;
        RECT 2621.640 18.060 2621.900 18.320 ;
        RECT 2857.160 18.060 2857.420 18.320 ;
      LAYER met2 ;
        RECT 2619.260 1700.410 2619.540 1704.000 ;
        RECT 2619.260 1700.270 2621.840 1700.410 ;
        RECT 2619.260 1700.000 2619.540 1700.270 ;
        RECT 2621.700 18.350 2621.840 1700.270 ;
        RECT 2621.640 18.030 2621.900 18.350 ;
        RECT 2857.160 18.030 2857.420 18.350 ;
        RECT 2857.220 2.400 2857.360 18.030 ;
        RECT 2857.010 -4.800 2857.570 2.400 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2628.460 1700.000 2628.740 1704.000 ;
        RECT 2628.600 16.845 2628.740 1700.000 ;
        RECT 2628.530 16.475 2628.810 16.845 ;
        RECT 2875.090 16.475 2875.370 16.845 ;
        RECT 2875.160 2.400 2875.300 16.475 ;
        RECT 2874.950 -4.800 2875.510 2.400 ;
      LAYER via2 ;
        RECT 2628.530 16.520 2628.810 16.800 ;
        RECT 2875.090 16.520 2875.370 16.800 ;
      LAYER met3 ;
        RECT 2628.505 16.810 2628.835 16.825 ;
        RECT 2875.065 16.810 2875.395 16.825 ;
        RECT 2628.505 16.510 2875.395 16.810 ;
        RECT 2628.505 16.495 2628.835 16.510 ;
        RECT 2875.065 16.495 2875.395 16.510 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2845.705 16.745 2845.875 17.595 ;
      LAYER mcon ;
        RECT 2845.705 17.425 2845.875 17.595 ;
      LAYER met1 ;
        RECT 2637.710 1683.920 2638.030 1683.980 ;
        RECT 2642.310 1683.920 2642.630 1683.980 ;
        RECT 2637.710 1683.780 2642.630 1683.920 ;
        RECT 2637.710 1683.720 2638.030 1683.780 ;
        RECT 2642.310 1683.720 2642.630 1683.780 ;
        RECT 2642.310 17.580 2642.630 17.640 ;
        RECT 2845.645 17.580 2845.935 17.625 ;
        RECT 2642.310 17.440 2845.935 17.580 ;
        RECT 2642.310 17.380 2642.630 17.440 ;
        RECT 2845.645 17.395 2845.935 17.440 ;
        RECT 2845.645 16.900 2845.935 16.945 ;
        RECT 2893.010 16.900 2893.330 16.960 ;
        RECT 2845.645 16.760 2893.330 16.900 ;
        RECT 2845.645 16.715 2845.935 16.760 ;
        RECT 2893.010 16.700 2893.330 16.760 ;
      LAYER via ;
        RECT 2637.740 1683.720 2638.000 1683.980 ;
        RECT 2642.340 1683.720 2642.600 1683.980 ;
        RECT 2642.340 17.380 2642.600 17.640 ;
        RECT 2893.040 16.700 2893.300 16.960 ;
      LAYER met2 ;
        RECT 2637.660 1700.000 2637.940 1704.000 ;
        RECT 2637.800 1684.010 2637.940 1700.000 ;
        RECT 2637.740 1683.690 2638.000 1684.010 ;
        RECT 2642.340 1683.690 2642.600 1684.010 ;
        RECT 2642.400 17.670 2642.540 1683.690 ;
        RECT 2642.340 17.350 2642.600 17.670 ;
        RECT 2893.040 16.670 2893.300 16.990 ;
        RECT 2893.100 2.400 2893.240 16.670 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2646.910 1688.000 2647.230 1688.060 ;
        RECT 2866.790 1688.000 2867.110 1688.060 ;
        RECT 2646.910 1687.860 2867.110 1688.000 ;
        RECT 2646.910 1687.800 2647.230 1687.860 ;
        RECT 2866.790 1687.800 2867.110 1687.860 ;
        RECT 2866.790 17.920 2867.110 17.980 ;
        RECT 2910.950 17.920 2911.270 17.980 ;
        RECT 2866.790 17.780 2911.270 17.920 ;
        RECT 2866.790 17.720 2867.110 17.780 ;
        RECT 2910.950 17.720 2911.270 17.780 ;
      LAYER via ;
        RECT 2646.940 1687.800 2647.200 1688.060 ;
        RECT 2866.820 1687.800 2867.080 1688.060 ;
        RECT 2866.820 17.720 2867.080 17.980 ;
        RECT 2910.980 17.720 2911.240 17.980 ;
      LAYER met2 ;
        RECT 2646.860 1700.000 2647.140 1704.000 ;
        RECT 2647.000 1688.090 2647.140 1700.000 ;
        RECT 2646.940 1687.770 2647.200 1688.090 ;
        RECT 2866.820 1687.770 2867.080 1688.090 ;
        RECT 2866.880 18.010 2867.020 1687.770 ;
        RECT 2866.820 17.690 2867.080 18.010 ;
        RECT 2910.980 17.690 2911.240 18.010 ;
        RECT 2911.040 2.400 2911.180 17.690 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 858.890 45.120 859.210 45.180 ;
        RECT 1588.450 45.120 1588.770 45.180 ;
        RECT 858.890 44.980 1588.770 45.120 ;
        RECT 858.890 44.920 859.210 44.980 ;
        RECT 1588.450 44.920 1588.770 44.980 ;
      LAYER via ;
        RECT 858.920 44.920 859.180 45.180 ;
        RECT 1588.480 44.920 1588.740 45.180 ;
      LAYER met2 ;
        RECT 1590.700 1700.410 1590.980 1704.000 ;
        RECT 1588.540 1700.270 1590.980 1700.410 ;
        RECT 1588.540 45.210 1588.680 1700.270 ;
        RECT 1590.700 1700.000 1590.980 1700.270 ;
        RECT 858.920 44.890 859.180 45.210 ;
        RECT 1588.480 44.890 1588.740 45.210 ;
        RECT 858.980 2.400 859.120 44.890 ;
        RECT 858.770 -4.800 859.330 2.400 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1594.965 1497.445 1595.135 1545.555 ;
        RECT 1595.425 476.085 1595.595 524.195 ;
        RECT 1594.965 89.845 1595.135 137.955 ;
      LAYER mcon ;
        RECT 1594.965 1545.385 1595.135 1545.555 ;
        RECT 1595.425 524.025 1595.595 524.195 ;
        RECT 1594.965 137.785 1595.135 137.955 ;
      LAYER met1 ;
        RECT 1594.890 1676.780 1595.210 1676.840 ;
        RECT 1598.110 1676.780 1598.430 1676.840 ;
        RECT 1594.890 1676.640 1598.430 1676.780 ;
        RECT 1594.890 1676.580 1595.210 1676.640 ;
        RECT 1598.110 1676.580 1598.430 1676.640 ;
        RECT 1594.430 1559.140 1594.750 1559.200 ;
        RECT 1595.350 1559.140 1595.670 1559.200 ;
        RECT 1594.430 1559.000 1595.670 1559.140 ;
        RECT 1594.430 1558.940 1594.750 1559.000 ;
        RECT 1595.350 1558.940 1595.670 1559.000 ;
        RECT 1594.905 1545.540 1595.195 1545.585 ;
        RECT 1595.350 1545.540 1595.670 1545.600 ;
        RECT 1594.905 1545.400 1595.670 1545.540 ;
        RECT 1594.905 1545.355 1595.195 1545.400 ;
        RECT 1595.350 1545.340 1595.670 1545.400 ;
        RECT 1594.890 1497.600 1595.210 1497.660 ;
        RECT 1594.695 1497.460 1595.210 1497.600 ;
        RECT 1594.890 1497.400 1595.210 1497.460 ;
        RECT 1594.890 1400.700 1595.210 1400.760 ;
        RECT 1595.350 1400.700 1595.670 1400.760 ;
        RECT 1594.890 1400.560 1595.670 1400.700 ;
        RECT 1594.890 1400.500 1595.210 1400.560 ;
        RECT 1595.350 1400.500 1595.670 1400.560 ;
        RECT 1594.890 1304.140 1595.210 1304.200 ;
        RECT 1595.350 1304.140 1595.670 1304.200 ;
        RECT 1594.890 1304.000 1595.670 1304.140 ;
        RECT 1594.890 1303.940 1595.210 1304.000 ;
        RECT 1595.350 1303.940 1595.670 1304.000 ;
        RECT 1594.890 1159.300 1595.210 1159.360 ;
        RECT 1595.350 1159.300 1595.670 1159.360 ;
        RECT 1594.890 1159.160 1595.670 1159.300 ;
        RECT 1594.890 1159.100 1595.210 1159.160 ;
        RECT 1595.350 1159.100 1595.670 1159.160 ;
        RECT 1594.890 1062.740 1595.210 1062.800 ;
        RECT 1595.350 1062.740 1595.670 1062.800 ;
        RECT 1594.890 1062.600 1595.670 1062.740 ;
        RECT 1594.890 1062.540 1595.210 1062.600 ;
        RECT 1595.350 1062.540 1595.670 1062.600 ;
        RECT 1594.890 1014.120 1595.210 1014.180 ;
        RECT 1595.350 1014.120 1595.670 1014.180 ;
        RECT 1594.890 1013.980 1595.670 1014.120 ;
        RECT 1594.890 1013.920 1595.210 1013.980 ;
        RECT 1595.350 1013.920 1595.670 1013.980 ;
        RECT 1594.430 835.280 1594.750 835.340 ;
        RECT 1595.350 835.280 1595.670 835.340 ;
        RECT 1594.430 835.140 1595.670 835.280 ;
        RECT 1594.430 835.080 1594.750 835.140 ;
        RECT 1595.350 835.080 1595.670 835.140 ;
        RECT 1594.430 738.380 1594.750 738.440 ;
        RECT 1595.350 738.380 1595.670 738.440 ;
        RECT 1594.430 738.240 1595.670 738.380 ;
        RECT 1594.430 738.180 1594.750 738.240 ;
        RECT 1595.350 738.180 1595.670 738.240 ;
        RECT 1594.430 641.820 1594.750 641.880 ;
        RECT 1595.350 641.820 1595.670 641.880 ;
        RECT 1594.430 641.680 1595.670 641.820 ;
        RECT 1594.430 641.620 1594.750 641.680 ;
        RECT 1595.350 641.620 1595.670 641.680 ;
        RECT 1595.350 531.460 1595.670 531.720 ;
        RECT 1595.440 531.040 1595.580 531.460 ;
        RECT 1595.350 530.780 1595.670 531.040 ;
        RECT 1595.350 524.180 1595.670 524.240 ;
        RECT 1595.155 524.040 1595.670 524.180 ;
        RECT 1595.350 523.980 1595.670 524.040 ;
        RECT 1595.350 476.240 1595.670 476.300 ;
        RECT 1595.155 476.100 1595.670 476.240 ;
        RECT 1595.350 476.040 1595.670 476.100 ;
        RECT 1595.350 379.680 1595.670 379.740 ;
        RECT 1595.810 379.680 1596.130 379.740 ;
        RECT 1595.350 379.540 1596.130 379.680 ;
        RECT 1595.350 379.480 1595.670 379.540 ;
        RECT 1595.810 379.480 1596.130 379.540 ;
        RECT 1594.890 338.200 1595.210 338.260 ;
        RECT 1595.350 338.200 1595.670 338.260 ;
        RECT 1594.890 338.060 1595.670 338.200 ;
        RECT 1594.890 338.000 1595.210 338.060 ;
        RECT 1595.350 338.000 1595.670 338.060 ;
        RECT 1594.890 137.940 1595.210 138.000 ;
        RECT 1594.695 137.800 1595.210 137.940 ;
        RECT 1594.890 137.740 1595.210 137.800 ;
        RECT 1594.890 90.000 1595.210 90.060 ;
        RECT 1594.695 89.860 1595.210 90.000 ;
        RECT 1594.890 89.800 1595.210 89.860 ;
        RECT 876.830 45.460 877.150 45.520 ;
        RECT 1595.350 45.460 1595.670 45.520 ;
        RECT 876.830 45.320 1595.670 45.460 ;
        RECT 876.830 45.260 877.150 45.320 ;
        RECT 1595.350 45.260 1595.670 45.320 ;
      LAYER via ;
        RECT 1594.920 1676.580 1595.180 1676.840 ;
        RECT 1598.140 1676.580 1598.400 1676.840 ;
        RECT 1594.460 1558.940 1594.720 1559.200 ;
        RECT 1595.380 1558.940 1595.640 1559.200 ;
        RECT 1595.380 1545.340 1595.640 1545.600 ;
        RECT 1594.920 1497.400 1595.180 1497.660 ;
        RECT 1594.920 1400.500 1595.180 1400.760 ;
        RECT 1595.380 1400.500 1595.640 1400.760 ;
        RECT 1594.920 1303.940 1595.180 1304.200 ;
        RECT 1595.380 1303.940 1595.640 1304.200 ;
        RECT 1594.920 1159.100 1595.180 1159.360 ;
        RECT 1595.380 1159.100 1595.640 1159.360 ;
        RECT 1594.920 1062.540 1595.180 1062.800 ;
        RECT 1595.380 1062.540 1595.640 1062.800 ;
        RECT 1594.920 1013.920 1595.180 1014.180 ;
        RECT 1595.380 1013.920 1595.640 1014.180 ;
        RECT 1594.460 835.080 1594.720 835.340 ;
        RECT 1595.380 835.080 1595.640 835.340 ;
        RECT 1594.460 738.180 1594.720 738.440 ;
        RECT 1595.380 738.180 1595.640 738.440 ;
        RECT 1594.460 641.620 1594.720 641.880 ;
        RECT 1595.380 641.620 1595.640 641.880 ;
        RECT 1595.380 531.460 1595.640 531.720 ;
        RECT 1595.380 530.780 1595.640 531.040 ;
        RECT 1595.380 523.980 1595.640 524.240 ;
        RECT 1595.380 476.040 1595.640 476.300 ;
        RECT 1595.380 379.480 1595.640 379.740 ;
        RECT 1595.840 379.480 1596.100 379.740 ;
        RECT 1594.920 338.000 1595.180 338.260 ;
        RECT 1595.380 338.000 1595.640 338.260 ;
        RECT 1594.920 137.740 1595.180 138.000 ;
        RECT 1594.920 89.800 1595.180 90.060 ;
        RECT 876.860 45.260 877.120 45.520 ;
        RECT 1595.380 45.260 1595.640 45.520 ;
      LAYER met2 ;
        RECT 1599.900 1700.410 1600.180 1704.000 ;
        RECT 1598.200 1700.270 1600.180 1700.410 ;
        RECT 1598.200 1676.870 1598.340 1700.270 ;
        RECT 1599.900 1700.000 1600.180 1700.270 ;
        RECT 1594.920 1676.550 1595.180 1676.870 ;
        RECT 1598.140 1676.550 1598.400 1676.870 ;
        RECT 1594.980 1580.730 1595.120 1676.550 ;
        RECT 1594.520 1580.590 1595.120 1580.730 ;
        RECT 1594.520 1559.230 1594.660 1580.590 ;
        RECT 1594.460 1558.910 1594.720 1559.230 ;
        RECT 1595.380 1558.910 1595.640 1559.230 ;
        RECT 1595.440 1545.630 1595.580 1558.910 ;
        RECT 1595.380 1545.310 1595.640 1545.630 ;
        RECT 1594.920 1497.370 1595.180 1497.690 ;
        RECT 1594.980 1473.290 1595.120 1497.370 ;
        RECT 1594.980 1473.150 1595.580 1473.290 ;
        RECT 1595.440 1414.130 1595.580 1473.150 ;
        RECT 1594.980 1413.990 1595.580 1414.130 ;
        RECT 1594.980 1400.790 1595.120 1413.990 ;
        RECT 1594.920 1400.470 1595.180 1400.790 ;
        RECT 1595.380 1400.470 1595.640 1400.790 ;
        RECT 1595.440 1317.570 1595.580 1400.470 ;
        RECT 1594.980 1317.430 1595.580 1317.570 ;
        RECT 1594.980 1304.230 1595.120 1317.430 ;
        RECT 1594.920 1303.910 1595.180 1304.230 ;
        RECT 1595.380 1303.910 1595.640 1304.230 ;
        RECT 1595.440 1221.010 1595.580 1303.910 ;
        RECT 1594.980 1220.870 1595.580 1221.010 ;
        RECT 1594.980 1159.390 1595.120 1220.870 ;
        RECT 1594.920 1159.070 1595.180 1159.390 ;
        RECT 1595.380 1159.070 1595.640 1159.390 ;
        RECT 1595.440 1124.450 1595.580 1159.070 ;
        RECT 1594.980 1124.310 1595.580 1124.450 ;
        RECT 1594.980 1062.830 1595.120 1124.310 ;
        RECT 1594.920 1062.510 1595.180 1062.830 ;
        RECT 1595.380 1062.510 1595.640 1062.830 ;
        RECT 1595.440 1027.890 1595.580 1062.510 ;
        RECT 1594.980 1027.750 1595.580 1027.890 ;
        RECT 1594.980 1014.210 1595.120 1027.750 ;
        RECT 1594.920 1013.890 1595.180 1014.210 ;
        RECT 1595.380 1013.890 1595.640 1014.210 ;
        RECT 1595.440 835.370 1595.580 1013.890 ;
        RECT 1594.460 835.050 1594.720 835.370 ;
        RECT 1595.380 835.050 1595.640 835.370 ;
        RECT 1594.520 834.770 1594.660 835.050 ;
        RECT 1594.520 834.630 1595.120 834.770 ;
        RECT 1594.980 796.690 1595.120 834.630 ;
        RECT 1594.980 796.550 1595.580 796.690 ;
        RECT 1595.440 738.470 1595.580 796.550 ;
        RECT 1594.460 738.210 1594.720 738.470 ;
        RECT 1594.460 738.150 1595.120 738.210 ;
        RECT 1595.380 738.150 1595.640 738.470 ;
        RECT 1594.520 738.070 1595.120 738.150 ;
        RECT 1594.980 689.250 1595.120 738.070 ;
        RECT 1594.980 689.110 1595.580 689.250 ;
        RECT 1595.440 641.910 1595.580 689.110 ;
        RECT 1594.460 641.650 1594.720 641.910 ;
        RECT 1595.380 641.650 1595.640 641.910 ;
        RECT 1594.460 641.590 1595.640 641.650 ;
        RECT 1594.520 641.510 1595.580 641.590 ;
        RECT 1595.440 573.085 1595.580 641.510 ;
        RECT 1595.370 572.715 1595.650 573.085 ;
        RECT 1595.370 572.035 1595.650 572.405 ;
        RECT 1595.440 531.750 1595.580 572.035 ;
        RECT 1595.380 531.430 1595.640 531.750 ;
        RECT 1595.380 530.750 1595.640 531.070 ;
        RECT 1595.440 524.270 1595.580 530.750 ;
        RECT 1595.380 523.950 1595.640 524.270 ;
        RECT 1595.380 476.010 1595.640 476.330 ;
        RECT 1595.440 427.450 1595.580 476.010 ;
        RECT 1595.440 427.310 1596.040 427.450 ;
        RECT 1595.900 379.770 1596.040 427.310 ;
        RECT 1595.380 379.450 1595.640 379.770 ;
        RECT 1595.840 379.450 1596.100 379.770 ;
        RECT 1595.440 338.290 1595.580 379.450 ;
        RECT 1594.920 337.970 1595.180 338.290 ;
        RECT 1595.380 337.970 1595.640 338.290 ;
        RECT 1594.980 303.690 1595.120 337.970 ;
        RECT 1594.980 303.550 1595.580 303.690 ;
        RECT 1595.440 255.410 1595.580 303.550 ;
        RECT 1594.520 255.270 1595.580 255.410 ;
        RECT 1594.520 254.730 1594.660 255.270 ;
        RECT 1594.520 254.590 1595.120 254.730 ;
        RECT 1594.980 138.030 1595.120 254.590 ;
        RECT 1594.920 137.710 1595.180 138.030 ;
        RECT 1594.920 89.770 1595.180 90.090 ;
        RECT 1594.980 72.490 1595.120 89.770 ;
        RECT 1594.980 72.350 1595.580 72.490 ;
        RECT 1595.440 45.550 1595.580 72.350 ;
        RECT 876.860 45.230 877.120 45.550 ;
        RECT 1595.380 45.230 1595.640 45.550 ;
        RECT 876.920 2.400 877.060 45.230 ;
        RECT 876.710 -4.800 877.270 2.400 ;
      LAYER via2 ;
        RECT 1595.370 572.760 1595.650 573.040 ;
        RECT 1595.370 572.080 1595.650 572.360 ;
      LAYER met3 ;
        RECT 1595.345 573.050 1595.675 573.065 ;
        RECT 1594.670 572.750 1595.675 573.050 ;
        RECT 1594.670 572.370 1594.970 572.750 ;
        RECT 1595.345 572.735 1595.675 572.750 ;
        RECT 1595.345 572.370 1595.675 572.385 ;
        RECT 1594.670 572.070 1595.675 572.370 ;
        RECT 1595.345 572.055 1595.675 572.070 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 894.770 45.800 895.090 45.860 ;
        RECT 1607.770 45.800 1608.090 45.860 ;
        RECT 894.770 45.660 1608.090 45.800 ;
        RECT 894.770 45.600 895.090 45.660 ;
        RECT 1607.770 45.600 1608.090 45.660 ;
      LAYER via ;
        RECT 894.800 45.600 895.060 45.860 ;
        RECT 1607.800 45.600 1608.060 45.860 ;
      LAYER met2 ;
        RECT 1609.100 1700.410 1609.380 1704.000 ;
        RECT 1607.860 1700.270 1609.380 1700.410 ;
        RECT 1607.860 821.965 1608.000 1700.270 ;
        RECT 1609.100 1700.000 1609.380 1700.270 ;
        RECT 1607.790 821.595 1608.070 821.965 ;
        RECT 1607.790 820.915 1608.070 821.285 ;
        RECT 1607.860 45.890 1608.000 820.915 ;
        RECT 894.800 45.570 895.060 45.890 ;
        RECT 1607.800 45.570 1608.060 45.890 ;
        RECT 894.860 2.400 895.000 45.570 ;
        RECT 894.650 -4.800 895.210 2.400 ;
      LAYER via2 ;
        RECT 1607.790 821.640 1608.070 821.920 ;
        RECT 1607.790 820.960 1608.070 821.240 ;
      LAYER met3 ;
        RECT 1607.765 821.930 1608.095 821.945 ;
        RECT 1607.550 821.615 1608.095 821.930 ;
        RECT 1607.550 821.265 1607.850 821.615 ;
        RECT 1607.550 820.950 1608.095 821.265 ;
        RECT 1607.765 820.935 1608.095 820.950 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 912.710 46.140 913.030 46.200 ;
        RECT 1616.050 46.140 1616.370 46.200 ;
        RECT 912.710 46.000 1616.370 46.140 ;
        RECT 912.710 45.940 913.030 46.000 ;
        RECT 1616.050 45.940 1616.370 46.000 ;
      LAYER via ;
        RECT 912.740 45.940 913.000 46.200 ;
        RECT 1616.080 45.940 1616.340 46.200 ;
      LAYER met2 ;
        RECT 1618.300 1700.410 1618.580 1704.000 ;
        RECT 1616.140 1700.270 1618.580 1700.410 ;
        RECT 1616.140 46.230 1616.280 1700.270 ;
        RECT 1618.300 1700.000 1618.580 1700.270 ;
        RECT 912.740 45.910 913.000 46.230 ;
        RECT 1616.080 45.910 1616.340 46.230 ;
        RECT 912.800 2.400 912.940 45.910 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1622.105 1304.325 1622.275 1318.095 ;
        RECT 1622.105 1207.765 1622.275 1221.535 ;
        RECT 1622.105 917.745 1622.275 932.195 ;
        RECT 1622.565 572.645 1622.735 594.235 ;
        RECT 1622.565 483.225 1622.735 531.335 ;
        RECT 1622.565 282.965 1622.735 331.075 ;
        RECT 1622.565 144.925 1622.735 200.855 ;
        RECT 1622.105 89.845 1622.275 137.955 ;
      LAYER mcon ;
        RECT 1622.105 1317.925 1622.275 1318.095 ;
        RECT 1622.105 1221.365 1622.275 1221.535 ;
        RECT 1622.105 932.025 1622.275 932.195 ;
        RECT 1622.565 594.065 1622.735 594.235 ;
        RECT 1622.565 531.165 1622.735 531.335 ;
        RECT 1622.565 330.905 1622.735 331.075 ;
        RECT 1622.565 200.685 1622.735 200.855 ;
        RECT 1622.105 137.785 1622.275 137.955 ;
      LAYER met1 ;
        RECT 1622.030 1659.440 1622.350 1659.500 ;
        RECT 1625.250 1659.440 1625.570 1659.500 ;
        RECT 1622.030 1659.300 1625.570 1659.440 ;
        RECT 1622.030 1659.240 1622.350 1659.300 ;
        RECT 1625.250 1659.240 1625.570 1659.300 ;
        RECT 1622.490 1449.320 1622.810 1449.380 ;
        RECT 1623.410 1449.320 1623.730 1449.380 ;
        RECT 1622.490 1449.180 1623.730 1449.320 ;
        RECT 1622.490 1449.120 1622.810 1449.180 ;
        RECT 1623.410 1449.120 1623.730 1449.180 ;
        RECT 1622.030 1401.040 1622.350 1401.100 ;
        RECT 1623.410 1401.040 1623.730 1401.100 ;
        RECT 1622.030 1400.900 1623.730 1401.040 ;
        RECT 1622.030 1400.840 1622.350 1400.900 ;
        RECT 1623.410 1400.840 1623.730 1400.900 ;
        RECT 1622.030 1318.080 1622.350 1318.140 ;
        RECT 1621.835 1317.940 1622.350 1318.080 ;
        RECT 1622.030 1317.880 1622.350 1317.940 ;
        RECT 1622.030 1304.480 1622.350 1304.540 ;
        RECT 1621.835 1304.340 1622.350 1304.480 ;
        RECT 1622.030 1304.280 1622.350 1304.340 ;
        RECT 1622.030 1221.520 1622.350 1221.580 ;
        RECT 1621.835 1221.380 1622.350 1221.520 ;
        RECT 1622.030 1221.320 1622.350 1221.380 ;
        RECT 1622.030 1207.920 1622.350 1207.980 ;
        RECT 1621.835 1207.780 1622.350 1207.920 ;
        RECT 1622.030 1207.720 1622.350 1207.780 ;
        RECT 1622.030 1207.240 1622.350 1207.300 ;
        RECT 1622.490 1207.240 1622.810 1207.300 ;
        RECT 1622.030 1207.100 1622.810 1207.240 ;
        RECT 1622.030 1207.040 1622.350 1207.100 ;
        RECT 1622.490 1207.040 1622.810 1207.100 ;
        RECT 1622.490 1080.080 1622.810 1080.140 ;
        RECT 1623.410 1080.080 1623.730 1080.140 ;
        RECT 1622.490 1079.940 1623.730 1080.080 ;
        RECT 1622.490 1079.880 1622.810 1079.940 ;
        RECT 1623.410 1079.880 1623.730 1079.940 ;
        RECT 1622.490 1007.320 1622.810 1007.380 ;
        RECT 1623.410 1007.320 1623.730 1007.380 ;
        RECT 1622.490 1007.180 1623.730 1007.320 ;
        RECT 1622.490 1007.120 1622.810 1007.180 ;
        RECT 1623.410 1007.120 1623.730 1007.180 ;
        RECT 1622.045 932.180 1622.335 932.225 ;
        RECT 1622.490 932.180 1622.810 932.240 ;
        RECT 1622.045 932.040 1622.810 932.180 ;
        RECT 1622.045 931.995 1622.335 932.040 ;
        RECT 1622.490 931.980 1622.810 932.040 ;
        RECT 1622.030 917.900 1622.350 917.960 ;
        RECT 1621.835 917.760 1622.350 917.900 ;
        RECT 1622.030 917.700 1622.350 917.760 ;
        RECT 1622.030 869.620 1622.350 869.680 ;
        RECT 1622.490 869.620 1622.810 869.680 ;
        RECT 1622.030 869.480 1622.810 869.620 ;
        RECT 1622.030 869.420 1622.350 869.480 ;
        RECT 1622.490 869.420 1622.810 869.480 ;
        RECT 1622.490 787.000 1622.810 787.060 ;
        RECT 1622.120 786.860 1622.810 787.000 ;
        RECT 1622.120 786.380 1622.260 786.860 ;
        RECT 1622.490 786.800 1622.810 786.860 ;
        RECT 1622.030 786.120 1622.350 786.380 ;
        RECT 1622.490 594.220 1622.810 594.280 ;
        RECT 1622.295 594.080 1622.810 594.220 ;
        RECT 1622.490 594.020 1622.810 594.080 ;
        RECT 1622.490 572.800 1622.810 572.860 ;
        RECT 1622.295 572.660 1622.810 572.800 ;
        RECT 1622.490 572.600 1622.810 572.660 ;
        RECT 1622.490 531.320 1622.810 531.380 ;
        RECT 1622.295 531.180 1622.810 531.320 ;
        RECT 1622.490 531.120 1622.810 531.180 ;
        RECT 1622.490 483.380 1622.810 483.440 ;
        RECT 1622.295 483.240 1622.810 483.380 ;
        RECT 1622.490 483.180 1622.810 483.240 ;
        RECT 1622.490 434.760 1622.810 434.820 ;
        RECT 1622.950 434.760 1623.270 434.820 ;
        RECT 1622.490 434.620 1623.270 434.760 ;
        RECT 1622.490 434.560 1622.810 434.620 ;
        RECT 1622.950 434.560 1623.270 434.620 ;
        RECT 1622.490 331.060 1622.810 331.120 ;
        RECT 1622.295 330.920 1622.810 331.060 ;
        RECT 1622.490 330.860 1622.810 330.920 ;
        RECT 1622.490 283.120 1622.810 283.180 ;
        RECT 1622.295 282.980 1622.810 283.120 ;
        RECT 1622.490 282.920 1622.810 282.980 ;
        RECT 1622.490 200.840 1622.810 200.900 ;
        RECT 1622.295 200.700 1622.810 200.840 ;
        RECT 1622.490 200.640 1622.810 200.700 ;
        RECT 1622.490 145.080 1622.810 145.140 ;
        RECT 1622.295 144.940 1622.810 145.080 ;
        RECT 1622.490 144.880 1622.810 144.940 ;
        RECT 1622.045 137.940 1622.335 137.985 ;
        RECT 1622.490 137.940 1622.810 138.000 ;
        RECT 1622.045 137.800 1622.810 137.940 ;
        RECT 1622.045 137.755 1622.335 137.800 ;
        RECT 1622.490 137.740 1622.810 137.800 ;
        RECT 1622.030 90.000 1622.350 90.060 ;
        RECT 1621.835 89.860 1622.350 90.000 ;
        RECT 1622.030 89.800 1622.350 89.860 ;
        RECT 930.190 46.480 930.510 46.540 ;
        RECT 1622.030 46.480 1622.350 46.540 ;
        RECT 930.190 46.340 1622.350 46.480 ;
        RECT 930.190 46.280 930.510 46.340 ;
        RECT 1622.030 46.280 1622.350 46.340 ;
      LAYER via ;
        RECT 1622.060 1659.240 1622.320 1659.500 ;
        RECT 1625.280 1659.240 1625.540 1659.500 ;
        RECT 1622.520 1449.120 1622.780 1449.380 ;
        RECT 1623.440 1449.120 1623.700 1449.380 ;
        RECT 1622.060 1400.840 1622.320 1401.100 ;
        RECT 1623.440 1400.840 1623.700 1401.100 ;
        RECT 1622.060 1317.880 1622.320 1318.140 ;
        RECT 1622.060 1304.280 1622.320 1304.540 ;
        RECT 1622.060 1221.320 1622.320 1221.580 ;
        RECT 1622.060 1207.720 1622.320 1207.980 ;
        RECT 1622.060 1207.040 1622.320 1207.300 ;
        RECT 1622.520 1207.040 1622.780 1207.300 ;
        RECT 1622.520 1079.880 1622.780 1080.140 ;
        RECT 1623.440 1079.880 1623.700 1080.140 ;
        RECT 1622.520 1007.120 1622.780 1007.380 ;
        RECT 1623.440 1007.120 1623.700 1007.380 ;
        RECT 1622.520 931.980 1622.780 932.240 ;
        RECT 1622.060 917.700 1622.320 917.960 ;
        RECT 1622.060 869.420 1622.320 869.680 ;
        RECT 1622.520 869.420 1622.780 869.680 ;
        RECT 1622.520 786.800 1622.780 787.060 ;
        RECT 1622.060 786.120 1622.320 786.380 ;
        RECT 1622.520 594.020 1622.780 594.280 ;
        RECT 1622.520 572.600 1622.780 572.860 ;
        RECT 1622.520 531.120 1622.780 531.380 ;
        RECT 1622.520 483.180 1622.780 483.440 ;
        RECT 1622.520 434.560 1622.780 434.820 ;
        RECT 1622.980 434.560 1623.240 434.820 ;
        RECT 1622.520 330.860 1622.780 331.120 ;
        RECT 1622.520 282.920 1622.780 283.180 ;
        RECT 1622.520 200.640 1622.780 200.900 ;
        RECT 1622.520 144.880 1622.780 145.140 ;
        RECT 1622.520 137.740 1622.780 138.000 ;
        RECT 1622.060 89.800 1622.320 90.060 ;
        RECT 930.220 46.280 930.480 46.540 ;
        RECT 1622.060 46.280 1622.320 46.540 ;
      LAYER met2 ;
        RECT 1627.500 1700.410 1627.780 1704.000 ;
        RECT 1625.340 1700.270 1627.780 1700.410 ;
        RECT 1625.340 1659.530 1625.480 1700.270 ;
        RECT 1627.500 1700.000 1627.780 1700.270 ;
        RECT 1622.060 1659.210 1622.320 1659.530 ;
        RECT 1625.280 1659.210 1625.540 1659.530 ;
        RECT 1622.120 1635.810 1622.260 1659.210 ;
        RECT 1622.120 1635.670 1622.720 1635.810 ;
        RECT 1622.580 1588.325 1622.720 1635.670 ;
        RECT 1622.510 1587.955 1622.790 1588.325 ;
        RECT 1622.050 1587.275 1622.330 1587.645 ;
        RECT 1622.120 1580.165 1622.260 1587.275 ;
        RECT 1622.050 1579.795 1622.330 1580.165 ;
        RECT 1623.430 1579.795 1623.710 1580.165 ;
        RECT 1623.500 1449.410 1623.640 1579.795 ;
        RECT 1622.520 1449.090 1622.780 1449.410 ;
        RECT 1623.440 1449.090 1623.700 1449.410 ;
        RECT 1622.580 1448.925 1622.720 1449.090 ;
        RECT 1622.510 1448.555 1622.790 1448.925 ;
        RECT 1623.430 1448.555 1623.710 1448.925 ;
        RECT 1623.500 1401.130 1623.640 1448.555 ;
        RECT 1622.060 1400.810 1622.320 1401.130 ;
        RECT 1623.440 1400.810 1623.700 1401.130 ;
        RECT 1622.120 1400.530 1622.260 1400.810 ;
        RECT 1622.120 1400.390 1622.720 1400.530 ;
        RECT 1622.580 1383.530 1622.720 1400.390 ;
        RECT 1622.120 1383.390 1622.720 1383.530 ;
        RECT 1622.120 1318.170 1622.260 1383.390 ;
        RECT 1622.060 1317.850 1622.320 1318.170 ;
        RECT 1622.060 1304.250 1622.320 1304.570 ;
        RECT 1622.120 1303.970 1622.260 1304.250 ;
        RECT 1622.120 1303.830 1622.720 1303.970 ;
        RECT 1622.580 1293.770 1622.720 1303.830 ;
        RECT 1622.120 1293.630 1622.720 1293.770 ;
        RECT 1622.120 1221.610 1622.260 1293.630 ;
        RECT 1622.060 1221.290 1622.320 1221.610 ;
        RECT 1622.060 1207.690 1622.320 1208.010 ;
        RECT 1622.120 1207.330 1622.260 1207.690 ;
        RECT 1622.060 1207.010 1622.320 1207.330 ;
        RECT 1622.520 1207.010 1622.780 1207.330 ;
        RECT 1622.580 1080.170 1622.720 1207.010 ;
        RECT 1622.520 1079.850 1622.780 1080.170 ;
        RECT 1623.440 1079.850 1623.700 1080.170 ;
        RECT 1623.500 1055.885 1623.640 1079.850 ;
        RECT 1622.510 1055.515 1622.790 1055.885 ;
        RECT 1623.430 1055.515 1623.710 1055.885 ;
        RECT 1622.580 1007.410 1622.720 1055.515 ;
        RECT 1622.520 1007.090 1622.780 1007.410 ;
        RECT 1623.440 1007.090 1623.700 1007.410 ;
        RECT 1623.500 959.325 1623.640 1007.090 ;
        RECT 1622.510 958.955 1622.790 959.325 ;
        RECT 1623.430 958.955 1623.710 959.325 ;
        RECT 1622.580 932.270 1622.720 958.955 ;
        RECT 1622.520 931.950 1622.780 932.270 ;
        RECT 1622.060 917.670 1622.320 917.990 ;
        RECT 1622.120 869.710 1622.260 917.670 ;
        RECT 1622.060 869.390 1622.320 869.710 ;
        RECT 1622.520 869.390 1622.780 869.710 ;
        RECT 1622.580 787.090 1622.720 869.390 ;
        RECT 1622.520 786.770 1622.780 787.090 ;
        RECT 1622.060 786.090 1622.320 786.410 ;
        RECT 1622.120 738.210 1622.260 786.090 ;
        RECT 1622.120 738.070 1622.720 738.210 ;
        RECT 1622.580 677.125 1622.720 738.070 ;
        RECT 1622.510 676.755 1622.790 677.125 ;
        RECT 1622.510 676.075 1622.790 676.445 ;
        RECT 1622.580 628.845 1622.720 676.075 ;
        RECT 1622.510 628.475 1622.790 628.845 ;
        RECT 1622.510 627.795 1622.790 628.165 ;
        RECT 1622.580 594.310 1622.720 627.795 ;
        RECT 1622.520 593.990 1622.780 594.310 ;
        RECT 1622.520 572.570 1622.780 572.890 ;
        RECT 1622.580 531.410 1622.720 572.570 ;
        RECT 1622.520 531.090 1622.780 531.410 ;
        RECT 1622.520 483.150 1622.780 483.470 ;
        RECT 1622.580 434.850 1622.720 483.150 ;
        RECT 1622.520 434.530 1622.780 434.850 ;
        RECT 1622.980 434.530 1623.240 434.850 ;
        RECT 1623.040 338.370 1623.180 434.530 ;
        RECT 1622.580 338.230 1623.180 338.370 ;
        RECT 1622.580 331.150 1622.720 338.230 ;
        RECT 1622.520 330.830 1622.780 331.150 ;
        RECT 1622.520 282.890 1622.780 283.210 ;
        RECT 1622.580 200.930 1622.720 282.890 ;
        RECT 1622.520 200.610 1622.780 200.930 ;
        RECT 1622.520 144.850 1622.780 145.170 ;
        RECT 1622.580 138.030 1622.720 144.850 ;
        RECT 1622.520 137.710 1622.780 138.030 ;
        RECT 1622.060 89.770 1622.320 90.090 ;
        RECT 1622.120 46.570 1622.260 89.770 ;
        RECT 930.220 46.250 930.480 46.570 ;
        RECT 1622.060 46.250 1622.320 46.570 ;
        RECT 930.280 2.400 930.420 46.250 ;
        RECT 930.070 -4.800 930.630 2.400 ;
      LAYER via2 ;
        RECT 1622.510 1588.000 1622.790 1588.280 ;
        RECT 1622.050 1587.320 1622.330 1587.600 ;
        RECT 1622.050 1579.840 1622.330 1580.120 ;
        RECT 1623.430 1579.840 1623.710 1580.120 ;
        RECT 1622.510 1448.600 1622.790 1448.880 ;
        RECT 1623.430 1448.600 1623.710 1448.880 ;
        RECT 1622.510 1055.560 1622.790 1055.840 ;
        RECT 1623.430 1055.560 1623.710 1055.840 ;
        RECT 1622.510 959.000 1622.790 959.280 ;
        RECT 1623.430 959.000 1623.710 959.280 ;
        RECT 1622.510 676.800 1622.790 677.080 ;
        RECT 1622.510 676.120 1622.790 676.400 ;
        RECT 1622.510 628.520 1622.790 628.800 ;
        RECT 1622.510 627.840 1622.790 628.120 ;
      LAYER met3 ;
        RECT 1622.485 1588.290 1622.815 1588.305 ;
        RECT 1621.350 1587.990 1622.815 1588.290 ;
        RECT 1621.350 1587.610 1621.650 1587.990 ;
        RECT 1622.485 1587.975 1622.815 1587.990 ;
        RECT 1622.025 1587.610 1622.355 1587.625 ;
        RECT 1621.350 1587.310 1622.355 1587.610 ;
        RECT 1622.025 1587.295 1622.355 1587.310 ;
        RECT 1622.025 1580.130 1622.355 1580.145 ;
        RECT 1623.405 1580.130 1623.735 1580.145 ;
        RECT 1622.025 1579.830 1623.735 1580.130 ;
        RECT 1622.025 1579.815 1622.355 1579.830 ;
        RECT 1623.405 1579.815 1623.735 1579.830 ;
        RECT 1622.485 1448.890 1622.815 1448.905 ;
        RECT 1623.405 1448.890 1623.735 1448.905 ;
        RECT 1622.485 1448.590 1623.735 1448.890 ;
        RECT 1622.485 1448.575 1622.815 1448.590 ;
        RECT 1623.405 1448.575 1623.735 1448.590 ;
        RECT 1622.485 1055.850 1622.815 1055.865 ;
        RECT 1623.405 1055.850 1623.735 1055.865 ;
        RECT 1622.485 1055.550 1623.735 1055.850 ;
        RECT 1622.485 1055.535 1622.815 1055.550 ;
        RECT 1623.405 1055.535 1623.735 1055.550 ;
        RECT 1622.485 959.290 1622.815 959.305 ;
        RECT 1623.405 959.290 1623.735 959.305 ;
        RECT 1622.485 958.990 1623.735 959.290 ;
        RECT 1622.485 958.975 1622.815 958.990 ;
        RECT 1623.405 958.975 1623.735 958.990 ;
        RECT 1622.485 677.090 1622.815 677.105 ;
        RECT 1622.270 676.775 1622.815 677.090 ;
        RECT 1622.270 676.425 1622.570 676.775 ;
        RECT 1622.270 676.110 1622.815 676.425 ;
        RECT 1622.485 676.095 1622.815 676.110 ;
        RECT 1622.485 628.495 1622.815 628.825 ;
        RECT 1622.500 628.145 1622.800 628.495 ;
        RECT 1622.485 627.815 1622.815 628.145 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 948.130 46.820 948.450 46.880 ;
        RECT 1635.370 46.820 1635.690 46.880 ;
        RECT 948.130 46.680 1635.690 46.820 ;
        RECT 948.130 46.620 948.450 46.680 ;
        RECT 1635.370 46.620 1635.690 46.680 ;
      LAYER via ;
        RECT 948.160 46.620 948.420 46.880 ;
        RECT 1635.400 46.620 1635.660 46.880 ;
      LAYER met2 ;
        RECT 1636.700 1700.410 1636.980 1704.000 ;
        RECT 1635.460 1700.270 1636.980 1700.410 ;
        RECT 1635.460 46.910 1635.600 1700.270 ;
        RECT 1636.700 1700.000 1636.980 1700.270 ;
        RECT 948.160 46.590 948.420 46.910 ;
        RECT 1635.400 46.590 1635.660 46.910 ;
        RECT 948.220 2.400 948.360 46.590 ;
        RECT 948.010 -4.800 948.570 2.400 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 966.070 47.160 966.390 47.220 ;
        RECT 1643.650 47.160 1643.970 47.220 ;
        RECT 966.070 47.020 1643.970 47.160 ;
        RECT 966.070 46.960 966.390 47.020 ;
        RECT 1643.650 46.960 1643.970 47.020 ;
      LAYER via ;
        RECT 966.100 46.960 966.360 47.220 ;
        RECT 1643.680 46.960 1643.940 47.220 ;
      LAYER met2 ;
        RECT 1645.900 1700.410 1646.180 1704.000 ;
        RECT 1643.740 1700.270 1646.180 1700.410 ;
        RECT 1643.740 47.250 1643.880 1700.270 ;
        RECT 1645.900 1700.000 1646.180 1700.270 ;
        RECT 966.100 46.930 966.360 47.250 ;
        RECT 1643.680 46.930 1643.940 47.250 ;
        RECT 966.160 2.400 966.300 46.930 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1650.165 531.505 1650.335 601.375 ;
        RECT 1649.705 234.685 1649.875 275.995 ;
        RECT 1650.165 131.325 1650.335 220.575 ;
        RECT 1650.625 47.345 1650.795 89.675 ;
      LAYER mcon ;
        RECT 1650.165 601.205 1650.335 601.375 ;
        RECT 1649.705 275.825 1649.875 275.995 ;
        RECT 1650.165 220.405 1650.335 220.575 ;
        RECT 1650.625 89.505 1650.795 89.675 ;
      LAYER met1 ;
        RECT 1650.090 1642.440 1650.410 1642.500 ;
        RECT 1652.850 1642.440 1653.170 1642.500 ;
        RECT 1650.090 1642.300 1653.170 1642.440 ;
        RECT 1650.090 1642.240 1650.410 1642.300 ;
        RECT 1652.850 1642.240 1653.170 1642.300 ;
        RECT 1650.090 1463.060 1650.410 1463.320 ;
        RECT 1650.180 1462.640 1650.320 1463.060 ;
        RECT 1650.090 1462.380 1650.410 1462.640 ;
        RECT 1650.090 1366.500 1650.410 1366.760 ;
        RECT 1650.180 1366.080 1650.320 1366.500 ;
        RECT 1650.090 1365.820 1650.410 1366.080 ;
        RECT 1650.090 1269.940 1650.410 1270.200 ;
        RECT 1650.180 1269.520 1650.320 1269.940 ;
        RECT 1650.090 1269.260 1650.410 1269.520 ;
        RECT 1650.550 1173.240 1650.870 1173.300 ;
        RECT 1650.180 1173.100 1650.870 1173.240 ;
        RECT 1650.180 1172.960 1650.320 1173.100 ;
        RECT 1650.550 1173.040 1650.870 1173.100 ;
        RECT 1650.090 1172.700 1650.410 1172.960 ;
        RECT 1650.550 1076.680 1650.870 1076.740 ;
        RECT 1650.180 1076.540 1650.870 1076.680 ;
        RECT 1650.180 1076.400 1650.320 1076.540 ;
        RECT 1650.550 1076.480 1650.870 1076.540 ;
        RECT 1650.090 1076.140 1650.410 1076.400 ;
        RECT 1650.090 965.980 1650.410 966.240 ;
        RECT 1650.180 965.840 1650.320 965.980 ;
        RECT 1650.550 965.840 1650.870 965.900 ;
        RECT 1650.180 965.700 1650.870 965.840 ;
        RECT 1650.550 965.640 1650.870 965.700 ;
        RECT 1649.630 917.900 1649.950 917.960 ;
        RECT 1650.550 917.900 1650.870 917.960 ;
        RECT 1649.630 917.760 1650.870 917.900 ;
        RECT 1649.630 917.700 1649.950 917.760 ;
        RECT 1650.550 917.700 1650.870 917.760 ;
        RECT 1649.630 883.360 1649.950 883.620 ;
        RECT 1649.720 882.880 1649.860 883.360 ;
        RECT 1650.090 882.880 1650.410 882.940 ;
        RECT 1649.720 882.740 1650.410 882.880 ;
        RECT 1650.090 882.680 1650.410 882.740 ;
        RECT 1649.630 821.000 1649.950 821.060 ;
        RECT 1650.550 821.000 1650.870 821.060 ;
        RECT 1649.630 820.860 1650.870 821.000 ;
        RECT 1649.630 820.800 1649.950 820.860 ;
        RECT 1650.550 820.800 1650.870 820.860 ;
        RECT 1650.090 642.160 1650.410 642.220 ;
        RECT 1649.720 642.020 1650.410 642.160 ;
        RECT 1649.720 641.540 1649.860 642.020 ;
        RECT 1650.090 641.960 1650.410 642.020 ;
        RECT 1649.630 641.280 1649.950 641.540 ;
        RECT 1649.630 601.360 1649.950 601.420 ;
        RECT 1650.105 601.360 1650.395 601.405 ;
        RECT 1649.630 601.220 1650.395 601.360 ;
        RECT 1649.630 601.160 1649.950 601.220 ;
        RECT 1650.105 601.175 1650.395 601.220 ;
        RECT 1650.090 531.660 1650.410 531.720 ;
        RECT 1649.895 531.520 1650.410 531.660 ;
        RECT 1650.090 531.460 1650.410 531.520 ;
        RECT 1649.630 282.780 1649.950 282.840 ;
        RECT 1650.090 282.780 1650.410 282.840 ;
        RECT 1649.630 282.640 1650.410 282.780 ;
        RECT 1649.630 282.580 1649.950 282.640 ;
        RECT 1650.090 282.580 1650.410 282.640 ;
        RECT 1649.630 275.980 1649.950 276.040 ;
        RECT 1649.435 275.840 1649.950 275.980 ;
        RECT 1649.630 275.780 1649.950 275.840 ;
        RECT 1649.645 234.840 1649.935 234.885 ;
        RECT 1650.090 234.840 1650.410 234.900 ;
        RECT 1649.645 234.700 1650.410 234.840 ;
        RECT 1649.645 234.655 1649.935 234.700 ;
        RECT 1650.090 234.640 1650.410 234.700 ;
        RECT 1650.090 220.560 1650.410 220.620 ;
        RECT 1649.895 220.420 1650.410 220.560 ;
        RECT 1650.090 220.360 1650.410 220.420 ;
        RECT 1650.105 131.480 1650.395 131.525 ;
        RECT 1650.550 131.480 1650.870 131.540 ;
        RECT 1650.105 131.340 1650.870 131.480 ;
        RECT 1650.105 131.295 1650.395 131.340 ;
        RECT 1650.550 131.280 1650.870 131.340 ;
        RECT 1650.550 89.660 1650.870 89.720 ;
        RECT 1650.355 89.520 1650.870 89.660 ;
        RECT 1650.550 89.460 1650.870 89.520 ;
        RECT 984.010 47.500 984.330 47.560 ;
        RECT 1650.565 47.500 1650.855 47.545 ;
        RECT 984.010 47.360 1650.855 47.500 ;
        RECT 984.010 47.300 984.330 47.360 ;
        RECT 1650.565 47.315 1650.855 47.360 ;
      LAYER via ;
        RECT 1650.120 1642.240 1650.380 1642.500 ;
        RECT 1652.880 1642.240 1653.140 1642.500 ;
        RECT 1650.120 1463.060 1650.380 1463.320 ;
        RECT 1650.120 1462.380 1650.380 1462.640 ;
        RECT 1650.120 1366.500 1650.380 1366.760 ;
        RECT 1650.120 1365.820 1650.380 1366.080 ;
        RECT 1650.120 1269.940 1650.380 1270.200 ;
        RECT 1650.120 1269.260 1650.380 1269.520 ;
        RECT 1650.580 1173.040 1650.840 1173.300 ;
        RECT 1650.120 1172.700 1650.380 1172.960 ;
        RECT 1650.580 1076.480 1650.840 1076.740 ;
        RECT 1650.120 1076.140 1650.380 1076.400 ;
        RECT 1650.120 965.980 1650.380 966.240 ;
        RECT 1650.580 965.640 1650.840 965.900 ;
        RECT 1649.660 917.700 1649.920 917.960 ;
        RECT 1650.580 917.700 1650.840 917.960 ;
        RECT 1649.660 883.360 1649.920 883.620 ;
        RECT 1650.120 882.680 1650.380 882.940 ;
        RECT 1649.660 820.800 1649.920 821.060 ;
        RECT 1650.580 820.800 1650.840 821.060 ;
        RECT 1650.120 641.960 1650.380 642.220 ;
        RECT 1649.660 641.280 1649.920 641.540 ;
        RECT 1649.660 601.160 1649.920 601.420 ;
        RECT 1650.120 531.460 1650.380 531.720 ;
        RECT 1649.660 282.580 1649.920 282.840 ;
        RECT 1650.120 282.580 1650.380 282.840 ;
        RECT 1649.660 275.780 1649.920 276.040 ;
        RECT 1650.120 234.640 1650.380 234.900 ;
        RECT 1650.120 220.360 1650.380 220.620 ;
        RECT 1650.580 131.280 1650.840 131.540 ;
        RECT 1650.580 89.460 1650.840 89.720 ;
        RECT 984.040 47.300 984.300 47.560 ;
      LAYER met2 ;
        RECT 1655.100 1700.410 1655.380 1704.000 ;
        RECT 1652.940 1700.270 1655.380 1700.410 ;
        RECT 1652.940 1642.530 1653.080 1700.270 ;
        RECT 1655.100 1700.000 1655.380 1700.270 ;
        RECT 1650.120 1642.210 1650.380 1642.530 ;
        RECT 1652.880 1642.210 1653.140 1642.530 ;
        RECT 1650.180 1463.350 1650.320 1642.210 ;
        RECT 1650.120 1463.030 1650.380 1463.350 ;
        RECT 1650.120 1462.350 1650.380 1462.670 ;
        RECT 1650.180 1366.790 1650.320 1462.350 ;
        RECT 1650.120 1366.470 1650.380 1366.790 ;
        RECT 1650.120 1365.790 1650.380 1366.110 ;
        RECT 1650.180 1270.230 1650.320 1365.790 ;
        RECT 1650.120 1269.910 1650.380 1270.230 ;
        RECT 1650.120 1269.230 1650.380 1269.550 ;
        RECT 1650.180 1207.410 1650.320 1269.230 ;
        RECT 1650.180 1207.270 1650.780 1207.410 ;
        RECT 1650.640 1173.330 1650.780 1207.270 ;
        RECT 1650.580 1173.010 1650.840 1173.330 ;
        RECT 1650.120 1172.670 1650.380 1172.990 ;
        RECT 1650.180 1110.850 1650.320 1172.670 ;
        RECT 1650.180 1110.710 1650.780 1110.850 ;
        RECT 1650.640 1076.770 1650.780 1110.710 ;
        RECT 1650.580 1076.450 1650.840 1076.770 ;
        RECT 1650.120 1076.110 1650.380 1076.430 ;
        RECT 1650.180 966.270 1650.320 1076.110 ;
        RECT 1650.120 965.950 1650.380 966.270 ;
        RECT 1650.580 965.610 1650.840 965.930 ;
        RECT 1650.640 917.990 1650.780 965.610 ;
        RECT 1649.660 917.670 1649.920 917.990 ;
        RECT 1650.580 917.670 1650.840 917.990 ;
        RECT 1649.720 883.650 1649.860 917.670 ;
        RECT 1649.660 883.330 1649.920 883.650 ;
        RECT 1650.120 882.650 1650.380 882.970 ;
        RECT 1650.180 846.330 1650.320 882.650 ;
        RECT 1650.180 846.190 1650.780 846.330 ;
        RECT 1650.640 821.285 1650.780 846.190 ;
        RECT 1649.650 820.915 1649.930 821.285 ;
        RECT 1650.570 820.915 1650.850 821.285 ;
        RECT 1649.660 820.770 1649.920 820.915 ;
        RECT 1650.580 820.770 1650.840 820.915 ;
        RECT 1650.640 725.405 1650.780 820.770 ;
        RECT 1650.570 725.035 1650.850 725.405 ;
        RECT 1650.110 724.355 1650.390 724.725 ;
        RECT 1650.180 642.250 1650.320 724.355 ;
        RECT 1650.120 641.930 1650.380 642.250 ;
        RECT 1649.660 641.250 1649.920 641.570 ;
        RECT 1649.720 601.450 1649.860 641.250 ;
        RECT 1649.660 601.130 1649.920 601.450 ;
        RECT 1650.120 531.430 1650.380 531.750 ;
        RECT 1650.180 497.490 1650.320 531.430 ;
        RECT 1650.180 497.350 1650.780 497.490 ;
        RECT 1650.640 496.130 1650.780 497.350 ;
        RECT 1650.180 495.990 1650.780 496.130 ;
        RECT 1650.180 303.690 1650.320 495.990 ;
        RECT 1649.720 303.550 1650.320 303.690 ;
        RECT 1649.720 303.010 1649.860 303.550 ;
        RECT 1649.720 302.870 1650.320 303.010 ;
        RECT 1650.180 282.870 1650.320 302.870 ;
        RECT 1649.660 282.550 1649.920 282.870 ;
        RECT 1650.120 282.550 1650.380 282.870 ;
        RECT 1649.720 276.070 1649.860 282.550 ;
        RECT 1649.660 275.750 1649.920 276.070 ;
        RECT 1650.120 234.610 1650.380 234.930 ;
        RECT 1650.180 220.650 1650.320 234.610 ;
        RECT 1650.120 220.330 1650.380 220.650 ;
        RECT 1650.580 131.250 1650.840 131.570 ;
        RECT 1650.640 89.750 1650.780 131.250 ;
        RECT 1650.580 89.430 1650.840 89.750 ;
        RECT 984.040 47.270 984.300 47.590 ;
        RECT 984.100 2.400 984.240 47.270 ;
        RECT 983.890 -4.800 984.450 2.400 ;
      LAYER via2 ;
        RECT 1649.650 820.960 1649.930 821.240 ;
        RECT 1650.570 820.960 1650.850 821.240 ;
        RECT 1650.570 725.080 1650.850 725.360 ;
        RECT 1650.110 724.400 1650.390 724.680 ;
      LAYER met3 ;
        RECT 1649.625 821.250 1649.955 821.265 ;
        RECT 1650.545 821.250 1650.875 821.265 ;
        RECT 1649.625 820.950 1650.875 821.250 ;
        RECT 1649.625 820.935 1649.955 820.950 ;
        RECT 1650.545 820.935 1650.875 820.950 ;
        RECT 1650.545 725.370 1650.875 725.385 ;
        RECT 1649.870 725.070 1650.875 725.370 ;
        RECT 1649.870 724.705 1650.170 725.070 ;
        RECT 1650.545 725.055 1650.875 725.070 ;
        RECT 1649.870 724.390 1650.415 724.705 ;
        RECT 1650.085 724.375 1650.415 724.390 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1484.030 1672.360 1484.350 1672.420 ;
        RECT 1487.710 1672.360 1488.030 1672.420 ;
        RECT 1484.030 1672.220 1488.030 1672.360 ;
        RECT 1484.030 1672.160 1484.350 1672.220 ;
        RECT 1487.710 1672.160 1488.030 1672.220 ;
        RECT 662.930 44.780 663.250 44.840 ;
        RECT 1484.030 44.780 1484.350 44.840 ;
        RECT 662.930 44.640 1484.350 44.780 ;
        RECT 662.930 44.580 663.250 44.640 ;
        RECT 1484.030 44.580 1484.350 44.640 ;
      LAYER via ;
        RECT 1484.060 1672.160 1484.320 1672.420 ;
        RECT 1487.740 1672.160 1488.000 1672.420 ;
        RECT 662.960 44.580 663.220 44.840 ;
        RECT 1484.060 44.580 1484.320 44.840 ;
      LAYER met2 ;
        RECT 1489.500 1700.410 1489.780 1704.000 ;
        RECT 1487.800 1700.270 1489.780 1700.410 ;
        RECT 1487.800 1672.450 1487.940 1700.270 ;
        RECT 1489.500 1700.000 1489.780 1700.270 ;
        RECT 1484.060 1672.130 1484.320 1672.450 ;
        RECT 1487.740 1672.130 1488.000 1672.450 ;
        RECT 1484.120 44.870 1484.260 1672.130 ;
        RECT 662.960 44.550 663.220 44.870 ;
        RECT 1484.060 44.550 1484.320 44.870 ;
        RECT 663.020 2.400 663.160 44.550 ;
        RECT 662.810 -4.800 663.370 2.400 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1001.950 47.840 1002.270 47.900 ;
        RECT 1662.970 47.840 1663.290 47.900 ;
        RECT 1001.950 47.700 1663.290 47.840 ;
        RECT 1001.950 47.640 1002.270 47.700 ;
        RECT 1662.970 47.640 1663.290 47.700 ;
      LAYER via ;
        RECT 1001.980 47.640 1002.240 47.900 ;
        RECT 1663.000 47.640 1663.260 47.900 ;
      LAYER met2 ;
        RECT 1664.300 1700.410 1664.580 1704.000 ;
        RECT 1663.060 1700.270 1664.580 1700.410 ;
        RECT 1663.060 47.930 1663.200 1700.270 ;
        RECT 1664.300 1700.000 1664.580 1700.270 ;
        RECT 1001.980 47.610 1002.240 47.930 ;
        RECT 1663.000 47.610 1663.260 47.930 ;
        RECT 1002.040 2.400 1002.180 47.610 ;
        RECT 1001.830 -4.800 1002.390 2.400 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1669.870 1658.080 1670.190 1658.140 ;
        RECT 1671.250 1658.080 1671.570 1658.140 ;
        RECT 1669.870 1657.940 1671.570 1658.080 ;
        RECT 1669.870 1657.880 1670.190 1657.940 ;
        RECT 1671.250 1657.880 1671.570 1657.940 ;
        RECT 1019.430 48.180 1019.750 48.240 ;
        RECT 1669.870 48.180 1670.190 48.240 ;
        RECT 1019.430 48.040 1670.190 48.180 ;
        RECT 1019.430 47.980 1019.750 48.040 ;
        RECT 1669.870 47.980 1670.190 48.040 ;
      LAYER via ;
        RECT 1669.900 1657.880 1670.160 1658.140 ;
        RECT 1671.280 1657.880 1671.540 1658.140 ;
        RECT 1019.460 47.980 1019.720 48.240 ;
        RECT 1669.900 47.980 1670.160 48.240 ;
      LAYER met2 ;
        RECT 1673.500 1700.410 1673.780 1704.000 ;
        RECT 1671.340 1700.270 1673.780 1700.410 ;
        RECT 1671.340 1658.170 1671.480 1700.270 ;
        RECT 1673.500 1700.000 1673.780 1700.270 ;
        RECT 1669.900 1657.850 1670.160 1658.170 ;
        RECT 1671.280 1657.850 1671.540 1658.170 ;
        RECT 1669.960 48.270 1670.100 1657.850 ;
        RECT 1019.460 47.950 1019.720 48.270 ;
        RECT 1669.900 47.950 1670.160 48.270 ;
        RECT 1019.520 2.400 1019.660 47.950 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1676.770 1678.140 1677.090 1678.200 ;
        RECT 1680.910 1678.140 1681.230 1678.200 ;
        RECT 1676.770 1678.000 1681.230 1678.140 ;
        RECT 1676.770 1677.940 1677.090 1678.000 ;
        RECT 1680.910 1677.940 1681.230 1678.000 ;
        RECT 1037.370 44.100 1037.690 44.160 ;
        RECT 1676.770 44.100 1677.090 44.160 ;
        RECT 1037.370 43.960 1677.090 44.100 ;
        RECT 1037.370 43.900 1037.690 43.960 ;
        RECT 1676.770 43.900 1677.090 43.960 ;
      LAYER via ;
        RECT 1676.800 1677.940 1677.060 1678.200 ;
        RECT 1680.940 1677.940 1681.200 1678.200 ;
        RECT 1037.400 43.900 1037.660 44.160 ;
        RECT 1676.800 43.900 1677.060 44.160 ;
      LAYER met2 ;
        RECT 1682.240 1700.410 1682.520 1704.000 ;
        RECT 1681.000 1700.270 1682.520 1700.410 ;
        RECT 1681.000 1678.230 1681.140 1700.270 ;
        RECT 1682.240 1700.000 1682.520 1700.270 ;
        RECT 1676.800 1677.910 1677.060 1678.230 ;
        RECT 1680.940 1677.910 1681.200 1678.230 ;
        RECT 1676.860 44.190 1677.000 1677.910 ;
        RECT 1037.400 43.870 1037.660 44.190 ;
        RECT 1676.800 43.870 1677.060 44.190 ;
        RECT 1037.460 2.400 1037.600 43.870 ;
        RECT 1037.250 -4.800 1037.810 2.400 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1054.850 44.440 1055.170 44.500 ;
        RECT 1691.030 44.440 1691.350 44.500 ;
        RECT 1054.850 44.300 1691.350 44.440 ;
        RECT 1054.850 44.240 1055.170 44.300 ;
        RECT 1691.030 44.240 1691.350 44.300 ;
      LAYER via ;
        RECT 1054.880 44.240 1055.140 44.500 ;
        RECT 1691.060 44.240 1691.320 44.500 ;
      LAYER met2 ;
        RECT 1691.440 1700.410 1691.720 1704.000 ;
        RECT 1691.120 1700.270 1691.720 1700.410 ;
        RECT 1691.120 44.530 1691.260 1700.270 ;
        RECT 1691.440 1700.000 1691.720 1700.270 ;
        RECT 1054.880 44.210 1055.140 44.530 ;
        RECT 1691.060 44.210 1691.320 44.530 ;
        RECT 1054.940 17.410 1055.080 44.210 ;
        RECT 1054.940 17.270 1055.540 17.410 ;
        RECT 1055.400 2.400 1055.540 17.270 ;
        RECT 1055.190 -4.800 1055.750 2.400 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1073.250 43.760 1073.570 43.820 ;
        RECT 1698.850 43.760 1699.170 43.820 ;
        RECT 1073.250 43.620 1699.170 43.760 ;
        RECT 1073.250 43.560 1073.570 43.620 ;
        RECT 1698.850 43.560 1699.170 43.620 ;
      LAYER via ;
        RECT 1073.280 43.560 1073.540 43.820 ;
        RECT 1698.880 43.560 1699.140 43.820 ;
      LAYER met2 ;
        RECT 1700.640 1700.410 1700.920 1704.000 ;
        RECT 1698.940 1700.270 1700.920 1700.410 ;
        RECT 1698.940 43.850 1699.080 1700.270 ;
        RECT 1700.640 1700.000 1700.920 1700.270 ;
        RECT 1073.280 43.530 1073.540 43.850 ;
        RECT 1698.880 43.530 1699.140 43.850 ;
        RECT 1073.340 2.400 1073.480 43.530 ;
        RECT 1073.130 -4.800 1073.690 2.400 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1704.370 1678.140 1704.690 1678.200 ;
        RECT 1708.510 1678.140 1708.830 1678.200 ;
        RECT 1704.370 1678.000 1708.830 1678.140 ;
        RECT 1704.370 1677.940 1704.690 1678.000 ;
        RECT 1708.510 1677.940 1708.830 1678.000 ;
        RECT 1090.730 43.080 1091.050 43.140 ;
        RECT 1704.370 43.080 1704.690 43.140 ;
        RECT 1090.730 42.940 1704.690 43.080 ;
        RECT 1090.730 42.880 1091.050 42.940 ;
        RECT 1704.370 42.880 1704.690 42.940 ;
      LAYER via ;
        RECT 1704.400 1677.940 1704.660 1678.200 ;
        RECT 1708.540 1677.940 1708.800 1678.200 ;
        RECT 1090.760 42.880 1091.020 43.140 ;
        RECT 1704.400 42.880 1704.660 43.140 ;
      LAYER met2 ;
        RECT 1709.840 1700.410 1710.120 1704.000 ;
        RECT 1708.600 1700.270 1710.120 1700.410 ;
        RECT 1708.600 1678.230 1708.740 1700.270 ;
        RECT 1709.840 1700.000 1710.120 1700.270 ;
        RECT 1704.400 1677.910 1704.660 1678.230 ;
        RECT 1708.540 1677.910 1708.800 1678.230 ;
        RECT 1704.460 43.170 1704.600 1677.910 ;
        RECT 1090.760 42.850 1091.020 43.170 ;
        RECT 1704.400 42.850 1704.660 43.170 ;
        RECT 1090.820 2.400 1090.960 42.850 ;
        RECT 1090.610 -4.800 1091.170 2.400 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1108.670 43.420 1108.990 43.480 ;
        RECT 1718.630 43.420 1718.950 43.480 ;
        RECT 1108.670 43.280 1718.950 43.420 ;
        RECT 1108.670 43.220 1108.990 43.280 ;
        RECT 1718.630 43.220 1718.950 43.280 ;
      LAYER via ;
        RECT 1108.700 43.220 1108.960 43.480 ;
        RECT 1718.660 43.220 1718.920 43.480 ;
      LAYER met2 ;
        RECT 1719.040 1700.410 1719.320 1704.000 ;
        RECT 1718.720 1700.270 1719.320 1700.410 ;
        RECT 1718.720 43.510 1718.860 1700.270 ;
        RECT 1719.040 1700.000 1719.320 1700.270 ;
        RECT 1108.700 43.190 1108.960 43.510 ;
        RECT 1718.660 43.190 1718.920 43.510 ;
        RECT 1108.760 2.400 1108.900 43.190 ;
        RECT 1108.550 -4.800 1109.110 2.400 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1126.610 42.740 1126.930 42.800 ;
        RECT 1725.990 42.740 1726.310 42.800 ;
        RECT 1126.610 42.600 1726.310 42.740 ;
        RECT 1126.610 42.540 1126.930 42.600 ;
        RECT 1725.990 42.540 1726.310 42.600 ;
      LAYER via ;
        RECT 1126.640 42.540 1126.900 42.800 ;
        RECT 1726.020 42.540 1726.280 42.800 ;
      LAYER met2 ;
        RECT 1728.240 1700.410 1728.520 1704.000 ;
        RECT 1726.080 1700.270 1728.520 1700.410 ;
        RECT 1726.080 42.830 1726.220 1700.270 ;
        RECT 1728.240 1700.000 1728.520 1700.270 ;
        RECT 1126.640 42.510 1126.900 42.830 ;
        RECT 1726.020 42.510 1726.280 42.830 ;
        RECT 1126.700 2.400 1126.840 42.510 ;
        RECT 1126.490 -4.800 1127.050 2.400 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1732.965 1545.725 1733.135 1559.155 ;
        RECT 1732.965 1449.165 1733.135 1497.275 ;
        RECT 1732.965 1352.605 1733.135 1400.715 ;
        RECT 1732.965 1256.045 1733.135 1304.155 ;
        RECT 1732.965 399.925 1733.135 434.775 ;
        RECT 1732.505 89.845 1732.675 137.955 ;
        RECT 1732.505 42.245 1732.675 48.195 ;
      LAYER mcon ;
        RECT 1732.965 1558.985 1733.135 1559.155 ;
        RECT 1732.965 1497.105 1733.135 1497.275 ;
        RECT 1732.965 1400.545 1733.135 1400.715 ;
        RECT 1732.965 1303.985 1733.135 1304.155 ;
        RECT 1732.965 434.605 1733.135 434.775 ;
        RECT 1732.505 137.785 1732.675 137.955 ;
        RECT 1732.505 48.025 1732.675 48.195 ;
      LAYER met1 ;
        RECT 1732.890 1559.140 1733.210 1559.200 ;
        RECT 1732.695 1559.000 1733.210 1559.140 ;
        RECT 1732.890 1558.940 1733.210 1559.000 ;
        RECT 1732.890 1545.880 1733.210 1545.940 ;
        RECT 1732.695 1545.740 1733.210 1545.880 ;
        RECT 1732.890 1545.680 1733.210 1545.740 ;
        RECT 1732.890 1497.260 1733.210 1497.320 ;
        RECT 1732.695 1497.120 1733.210 1497.260 ;
        RECT 1732.890 1497.060 1733.210 1497.120 ;
        RECT 1732.890 1449.320 1733.210 1449.380 ;
        RECT 1732.695 1449.180 1733.210 1449.320 ;
        RECT 1732.890 1449.120 1733.210 1449.180 ;
        RECT 1732.890 1400.700 1733.210 1400.760 ;
        RECT 1732.695 1400.560 1733.210 1400.700 ;
        RECT 1732.890 1400.500 1733.210 1400.560 ;
        RECT 1732.890 1352.760 1733.210 1352.820 ;
        RECT 1732.695 1352.620 1733.210 1352.760 ;
        RECT 1732.890 1352.560 1733.210 1352.620 ;
        RECT 1732.890 1304.140 1733.210 1304.200 ;
        RECT 1732.695 1304.000 1733.210 1304.140 ;
        RECT 1732.890 1303.940 1733.210 1304.000 ;
        RECT 1732.890 1256.200 1733.210 1256.260 ;
        RECT 1732.695 1256.060 1733.210 1256.200 ;
        RECT 1732.890 1256.000 1733.210 1256.060 ;
        RECT 1732.890 1159.300 1733.210 1159.360 ;
        RECT 1733.810 1159.300 1734.130 1159.360 ;
        RECT 1732.890 1159.160 1734.130 1159.300 ;
        RECT 1732.890 1159.100 1733.210 1159.160 ;
        RECT 1733.810 1159.100 1734.130 1159.160 ;
        RECT 1732.890 1062.740 1733.210 1062.800 ;
        RECT 1733.810 1062.740 1734.130 1062.800 ;
        RECT 1732.890 1062.600 1734.130 1062.740 ;
        RECT 1732.890 1062.540 1733.210 1062.600 ;
        RECT 1733.810 1062.540 1734.130 1062.600 ;
        RECT 1732.890 966.180 1733.210 966.240 ;
        RECT 1733.810 966.180 1734.130 966.240 ;
        RECT 1732.890 966.040 1734.130 966.180 ;
        RECT 1732.890 965.980 1733.210 966.040 ;
        RECT 1733.810 965.980 1734.130 966.040 ;
        RECT 1732.890 883.020 1733.210 883.280 ;
        RECT 1732.980 882.600 1733.120 883.020 ;
        RECT 1732.890 882.340 1733.210 882.600 ;
        RECT 1732.890 786.460 1733.210 786.720 ;
        RECT 1732.980 786.040 1733.120 786.460 ;
        RECT 1732.890 785.780 1733.210 786.040 ;
        RECT 1732.890 593.340 1733.210 593.600 ;
        RECT 1732.980 592.920 1733.120 593.340 ;
        RECT 1732.890 592.660 1733.210 592.920 ;
        RECT 1732.890 434.760 1733.210 434.820 ;
        RECT 1732.695 434.620 1733.210 434.760 ;
        RECT 1732.890 434.560 1733.210 434.620 ;
        RECT 1732.890 400.080 1733.210 400.140 ;
        RECT 1732.695 399.940 1733.210 400.080 ;
        RECT 1732.890 399.880 1733.210 399.940 ;
        RECT 1732.890 331.060 1733.210 331.120 ;
        RECT 1733.350 331.060 1733.670 331.120 ;
        RECT 1732.890 330.920 1733.670 331.060 ;
        RECT 1732.890 330.860 1733.210 330.920 ;
        RECT 1733.350 330.860 1733.670 330.920 ;
        RECT 1732.430 137.940 1732.750 138.000 ;
        RECT 1732.235 137.800 1732.750 137.940 ;
        RECT 1732.430 137.740 1732.750 137.800 ;
        RECT 1732.430 90.000 1732.750 90.060 ;
        RECT 1732.235 89.860 1732.750 90.000 ;
        RECT 1732.430 89.800 1732.750 89.860 ;
        RECT 1732.430 48.180 1732.750 48.240 ;
        RECT 1732.235 48.040 1732.750 48.180 ;
        RECT 1732.430 47.980 1732.750 48.040 ;
        RECT 1144.550 42.400 1144.870 42.460 ;
        RECT 1732.445 42.400 1732.735 42.445 ;
        RECT 1144.550 42.260 1732.735 42.400 ;
        RECT 1144.550 42.200 1144.870 42.260 ;
        RECT 1732.445 42.215 1732.735 42.260 ;
      LAYER via ;
        RECT 1732.920 1558.940 1733.180 1559.200 ;
        RECT 1732.920 1545.680 1733.180 1545.940 ;
        RECT 1732.920 1497.060 1733.180 1497.320 ;
        RECT 1732.920 1449.120 1733.180 1449.380 ;
        RECT 1732.920 1400.500 1733.180 1400.760 ;
        RECT 1732.920 1352.560 1733.180 1352.820 ;
        RECT 1732.920 1303.940 1733.180 1304.200 ;
        RECT 1732.920 1256.000 1733.180 1256.260 ;
        RECT 1732.920 1159.100 1733.180 1159.360 ;
        RECT 1733.840 1159.100 1734.100 1159.360 ;
        RECT 1732.920 1062.540 1733.180 1062.800 ;
        RECT 1733.840 1062.540 1734.100 1062.800 ;
        RECT 1732.920 965.980 1733.180 966.240 ;
        RECT 1733.840 965.980 1734.100 966.240 ;
        RECT 1732.920 883.020 1733.180 883.280 ;
        RECT 1732.920 882.340 1733.180 882.600 ;
        RECT 1732.920 786.460 1733.180 786.720 ;
        RECT 1732.920 785.780 1733.180 786.040 ;
        RECT 1732.920 593.340 1733.180 593.600 ;
        RECT 1732.920 592.660 1733.180 592.920 ;
        RECT 1732.920 434.560 1733.180 434.820 ;
        RECT 1732.920 399.880 1733.180 400.140 ;
        RECT 1732.920 330.860 1733.180 331.120 ;
        RECT 1733.380 330.860 1733.640 331.120 ;
        RECT 1732.460 137.740 1732.720 138.000 ;
        RECT 1732.460 89.800 1732.720 90.060 ;
        RECT 1732.460 47.980 1732.720 48.240 ;
        RECT 1144.580 42.200 1144.840 42.460 ;
      LAYER met2 ;
        RECT 1737.440 1700.410 1737.720 1704.000 ;
        RECT 1735.740 1700.270 1737.720 1700.410 ;
        RECT 1735.740 1656.210 1735.880 1700.270 ;
        RECT 1737.440 1700.000 1737.720 1700.270 ;
        RECT 1732.980 1656.070 1735.880 1656.210 ;
        RECT 1732.980 1559.230 1733.120 1656.070 ;
        RECT 1732.920 1558.910 1733.180 1559.230 ;
        RECT 1732.920 1545.650 1733.180 1545.970 ;
        RECT 1732.980 1497.350 1733.120 1545.650 ;
        RECT 1732.920 1497.030 1733.180 1497.350 ;
        RECT 1732.920 1449.090 1733.180 1449.410 ;
        RECT 1732.980 1400.790 1733.120 1449.090 ;
        RECT 1732.920 1400.470 1733.180 1400.790 ;
        RECT 1732.920 1352.530 1733.180 1352.850 ;
        RECT 1732.980 1304.230 1733.120 1352.530 ;
        RECT 1732.920 1303.910 1733.180 1304.230 ;
        RECT 1732.920 1255.970 1733.180 1256.290 ;
        RECT 1732.980 1207.525 1733.120 1255.970 ;
        RECT 1732.910 1207.155 1733.190 1207.525 ;
        RECT 1733.830 1207.155 1734.110 1207.525 ;
        RECT 1733.900 1159.390 1734.040 1207.155 ;
        RECT 1732.920 1159.070 1733.180 1159.390 ;
        RECT 1733.840 1159.070 1734.100 1159.390 ;
        RECT 1732.980 1110.965 1733.120 1159.070 ;
        RECT 1732.910 1110.595 1733.190 1110.965 ;
        RECT 1733.830 1110.595 1734.110 1110.965 ;
        RECT 1733.900 1062.830 1734.040 1110.595 ;
        RECT 1732.920 1062.510 1733.180 1062.830 ;
        RECT 1733.840 1062.510 1734.100 1062.830 ;
        RECT 1732.980 1014.405 1733.120 1062.510 ;
        RECT 1732.910 1014.035 1733.190 1014.405 ;
        RECT 1733.830 1014.035 1734.110 1014.405 ;
        RECT 1733.900 966.270 1734.040 1014.035 ;
        RECT 1732.920 965.950 1733.180 966.270 ;
        RECT 1733.840 965.950 1734.100 966.270 ;
        RECT 1732.980 883.310 1733.120 965.950 ;
        RECT 1732.920 882.990 1733.180 883.310 ;
        RECT 1732.920 882.310 1733.180 882.630 ;
        RECT 1732.980 786.750 1733.120 882.310 ;
        RECT 1732.920 786.430 1733.180 786.750 ;
        RECT 1732.920 785.750 1733.180 786.070 ;
        RECT 1732.980 690.610 1733.120 785.750 ;
        RECT 1732.520 690.470 1733.120 690.610 ;
        RECT 1732.520 689.930 1732.660 690.470 ;
        RECT 1732.520 689.790 1733.120 689.930 ;
        RECT 1732.980 593.630 1733.120 689.790 ;
        RECT 1732.920 593.310 1733.180 593.630 ;
        RECT 1732.920 592.630 1733.180 592.950 ;
        RECT 1732.980 497.490 1733.120 592.630 ;
        RECT 1732.520 497.350 1733.120 497.490 ;
        RECT 1732.520 496.810 1732.660 497.350 ;
        RECT 1732.520 496.670 1733.120 496.810 ;
        RECT 1732.980 434.850 1733.120 496.670 ;
        RECT 1732.920 434.530 1733.180 434.850 ;
        RECT 1732.920 399.850 1733.180 400.170 ;
        RECT 1732.980 331.150 1733.120 399.850 ;
        RECT 1732.920 330.830 1733.180 331.150 ;
        RECT 1733.380 330.830 1733.640 331.150 ;
        RECT 1733.440 303.520 1733.580 330.830 ;
        RECT 1732.980 303.380 1733.580 303.520 ;
        RECT 1732.980 169.050 1733.120 303.380 ;
        RECT 1732.520 168.910 1733.120 169.050 ;
        RECT 1732.520 138.030 1732.660 168.910 ;
        RECT 1732.460 137.710 1732.720 138.030 ;
        RECT 1732.460 89.770 1732.720 90.090 ;
        RECT 1732.520 48.270 1732.660 89.770 ;
        RECT 1732.460 47.950 1732.720 48.270 ;
        RECT 1144.580 42.170 1144.840 42.490 ;
        RECT 1144.640 2.400 1144.780 42.170 ;
        RECT 1144.430 -4.800 1144.990 2.400 ;
      LAYER via2 ;
        RECT 1732.910 1207.200 1733.190 1207.480 ;
        RECT 1733.830 1207.200 1734.110 1207.480 ;
        RECT 1732.910 1110.640 1733.190 1110.920 ;
        RECT 1733.830 1110.640 1734.110 1110.920 ;
        RECT 1732.910 1014.080 1733.190 1014.360 ;
        RECT 1733.830 1014.080 1734.110 1014.360 ;
      LAYER met3 ;
        RECT 1732.885 1207.490 1733.215 1207.505 ;
        RECT 1733.805 1207.490 1734.135 1207.505 ;
        RECT 1732.885 1207.190 1734.135 1207.490 ;
        RECT 1732.885 1207.175 1733.215 1207.190 ;
        RECT 1733.805 1207.175 1734.135 1207.190 ;
        RECT 1732.885 1110.930 1733.215 1110.945 ;
        RECT 1733.805 1110.930 1734.135 1110.945 ;
        RECT 1732.885 1110.630 1734.135 1110.930 ;
        RECT 1732.885 1110.615 1733.215 1110.630 ;
        RECT 1733.805 1110.615 1734.135 1110.630 ;
        RECT 1732.885 1014.370 1733.215 1014.385 ;
        RECT 1733.805 1014.370 1734.135 1014.385 ;
        RECT 1732.885 1014.070 1734.135 1014.370 ;
        RECT 1732.885 1014.055 1733.215 1014.070 ;
        RECT 1733.805 1014.055 1734.135 1014.070 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1162.490 42.060 1162.810 42.120 ;
        RECT 1746.230 42.060 1746.550 42.120 ;
        RECT 1162.490 41.920 1746.550 42.060 ;
        RECT 1162.490 41.860 1162.810 41.920 ;
        RECT 1746.230 41.860 1746.550 41.920 ;
      LAYER via ;
        RECT 1162.520 41.860 1162.780 42.120 ;
        RECT 1746.260 41.860 1746.520 42.120 ;
      LAYER met2 ;
        RECT 1746.640 1700.410 1746.920 1704.000 ;
        RECT 1746.320 1700.270 1746.920 1700.410 ;
        RECT 1746.320 42.150 1746.460 1700.270 ;
        RECT 1746.640 1700.000 1746.920 1700.270 ;
        RECT 1162.520 41.830 1162.780 42.150 ;
        RECT 1746.260 41.830 1746.520 42.150 ;
        RECT 1162.580 2.400 1162.720 41.830 ;
        RECT 1162.370 -4.800 1162.930 2.400 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1498.700 1700.410 1498.980 1704.000 ;
        RECT 1497.920 1700.270 1498.980 1700.410 ;
        RECT 1497.920 44.725 1498.060 1700.270 ;
        RECT 1498.700 1700.000 1498.980 1700.270 ;
        RECT 680.430 44.355 680.710 44.725 ;
        RECT 1497.850 44.355 1498.130 44.725 ;
        RECT 680.500 2.400 680.640 44.355 ;
        RECT 680.290 -4.800 680.850 2.400 ;
      LAYER via2 ;
        RECT 680.430 44.400 680.710 44.680 ;
        RECT 1497.850 44.400 1498.130 44.680 ;
      LAYER met3 ;
        RECT 680.405 44.690 680.735 44.705 ;
        RECT 1497.825 44.690 1498.155 44.705 ;
        RECT 680.405 44.390 1498.155 44.690 ;
        RECT 680.405 44.375 680.735 44.390 ;
        RECT 1497.825 44.375 1498.155 44.390 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1179.970 41.720 1180.290 41.780 ;
        RECT 1753.590 41.720 1753.910 41.780 ;
        RECT 1179.970 41.580 1753.910 41.720 ;
        RECT 1179.970 41.520 1180.290 41.580 ;
        RECT 1753.590 41.520 1753.910 41.580 ;
      LAYER via ;
        RECT 1180.000 41.520 1180.260 41.780 ;
        RECT 1753.620 41.520 1753.880 41.780 ;
      LAYER met2 ;
        RECT 1755.840 1700.410 1756.120 1704.000 ;
        RECT 1753.680 1700.270 1756.120 1700.410 ;
        RECT 1753.680 41.810 1753.820 1700.270 ;
        RECT 1755.840 1700.000 1756.120 1700.270 ;
        RECT 1180.000 41.490 1180.260 41.810 ;
        RECT 1753.620 41.490 1753.880 41.810 ;
        RECT 1180.060 2.400 1180.200 41.490 ;
        RECT 1179.850 -4.800 1180.410 2.400 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1760.565 1439.645 1760.735 1490.475 ;
        RECT 1760.565 965.685 1760.735 1007.335 ;
        RECT 1760.565 814.385 1760.735 903.975 ;
        RECT 1760.105 331.245 1760.275 386.835 ;
      LAYER mcon ;
        RECT 1760.565 1490.305 1760.735 1490.475 ;
        RECT 1760.565 1007.165 1760.735 1007.335 ;
        RECT 1760.565 903.805 1760.735 903.975 ;
        RECT 1760.105 386.665 1760.275 386.835 ;
      LAYER met1 ;
        RECT 1760.030 1666.580 1760.350 1666.640 ;
        RECT 1763.250 1666.580 1763.570 1666.640 ;
        RECT 1760.030 1666.440 1763.570 1666.580 ;
        RECT 1760.030 1666.380 1760.350 1666.440 ;
        RECT 1763.250 1666.380 1763.570 1666.440 ;
        RECT 1760.490 1580.220 1760.810 1580.280 ;
        RECT 1761.410 1580.220 1761.730 1580.280 ;
        RECT 1760.490 1580.080 1761.730 1580.220 ;
        RECT 1760.490 1580.020 1760.810 1580.080 ;
        RECT 1761.410 1580.020 1761.730 1580.080 ;
        RECT 1760.490 1531.940 1760.810 1532.000 ;
        RECT 1761.410 1531.940 1761.730 1532.000 ;
        RECT 1760.490 1531.800 1761.730 1531.940 ;
        RECT 1760.490 1531.740 1760.810 1531.800 ;
        RECT 1761.410 1531.740 1761.730 1531.800 ;
        RECT 1760.490 1490.460 1760.810 1490.520 ;
        RECT 1760.295 1490.320 1760.810 1490.460 ;
        RECT 1760.490 1490.260 1760.810 1490.320 ;
        RECT 1760.490 1439.800 1760.810 1439.860 ;
        RECT 1760.295 1439.660 1760.810 1439.800 ;
        RECT 1760.490 1439.600 1760.810 1439.660 ;
        RECT 1760.490 1400.700 1760.810 1400.760 ;
        RECT 1761.410 1400.700 1761.730 1400.760 ;
        RECT 1760.490 1400.560 1761.730 1400.700 ;
        RECT 1760.490 1400.500 1760.810 1400.560 ;
        RECT 1761.410 1400.500 1761.730 1400.560 ;
        RECT 1759.110 1297.340 1759.430 1297.400 ;
        RECT 1760.030 1297.340 1760.350 1297.400 ;
        RECT 1759.110 1297.200 1760.350 1297.340 ;
        RECT 1759.110 1297.140 1759.430 1297.200 ;
        RECT 1760.030 1297.140 1760.350 1297.200 ;
        RECT 1760.030 1256.200 1760.350 1256.260 ;
        RECT 1760.490 1256.200 1760.810 1256.260 ;
        RECT 1760.030 1256.060 1760.810 1256.200 ;
        RECT 1760.030 1256.000 1760.350 1256.060 ;
        RECT 1760.490 1256.000 1760.810 1256.060 ;
        RECT 1759.110 1172.560 1759.430 1172.620 ;
        RECT 1760.490 1172.560 1760.810 1172.620 ;
        RECT 1759.110 1172.420 1760.810 1172.560 ;
        RECT 1759.110 1172.360 1759.430 1172.420 ;
        RECT 1760.490 1172.360 1760.810 1172.420 ;
        RECT 1759.110 1104.220 1759.430 1104.280 ;
        RECT 1760.030 1104.220 1760.350 1104.280 ;
        RECT 1759.110 1104.080 1760.350 1104.220 ;
        RECT 1759.110 1104.020 1759.430 1104.080 ;
        RECT 1760.030 1104.020 1760.350 1104.080 ;
        RECT 1760.030 1062.740 1760.350 1062.800 ;
        RECT 1760.490 1062.740 1760.810 1062.800 ;
        RECT 1760.030 1062.600 1760.810 1062.740 ;
        RECT 1760.030 1062.540 1760.350 1062.600 ;
        RECT 1760.490 1062.540 1760.810 1062.600 ;
        RECT 1759.110 1055.600 1759.430 1055.660 ;
        RECT 1760.030 1055.600 1760.350 1055.660 ;
        RECT 1759.110 1055.460 1760.350 1055.600 ;
        RECT 1759.110 1055.400 1759.430 1055.460 ;
        RECT 1760.030 1055.400 1760.350 1055.460 ;
        RECT 1760.490 1007.320 1760.810 1007.380 ;
        RECT 1760.295 1007.180 1760.810 1007.320 ;
        RECT 1760.490 1007.120 1760.810 1007.180 ;
        RECT 1760.490 965.840 1760.810 965.900 ;
        RECT 1760.295 965.700 1760.810 965.840 ;
        RECT 1760.490 965.640 1760.810 965.700 ;
        RECT 1760.030 917.900 1760.350 917.960 ;
        RECT 1760.950 917.900 1761.270 917.960 ;
        RECT 1760.030 917.760 1761.270 917.900 ;
        RECT 1760.030 917.700 1760.350 917.760 ;
        RECT 1760.950 917.700 1761.270 917.760 ;
        RECT 1760.030 903.960 1760.350 904.020 ;
        RECT 1760.505 903.960 1760.795 904.005 ;
        RECT 1760.030 903.820 1760.795 903.960 ;
        RECT 1760.030 903.760 1760.350 903.820 ;
        RECT 1760.505 903.775 1760.795 903.820 ;
        RECT 1760.490 814.540 1760.810 814.600 ;
        RECT 1760.295 814.400 1760.810 814.540 ;
        RECT 1760.490 814.340 1760.810 814.400 ;
        RECT 1760.030 724.440 1760.350 724.500 ;
        RECT 1760.950 724.440 1761.270 724.500 ;
        RECT 1760.030 724.300 1761.270 724.440 ;
        RECT 1760.030 724.240 1760.350 724.300 ;
        RECT 1760.950 724.240 1761.270 724.300 ;
        RECT 1759.110 475.560 1759.430 475.620 ;
        RECT 1760.950 475.560 1761.270 475.620 ;
        RECT 1759.110 475.420 1761.270 475.560 ;
        RECT 1759.110 475.360 1759.430 475.420 ;
        RECT 1760.950 475.360 1761.270 475.420 ;
        RECT 1760.490 427.960 1760.810 428.020 ;
        RECT 1760.950 427.960 1761.270 428.020 ;
        RECT 1760.490 427.820 1761.270 427.960 ;
        RECT 1760.490 427.760 1760.810 427.820 ;
        RECT 1760.950 427.760 1761.270 427.820 ;
        RECT 1760.045 386.820 1760.335 386.865 ;
        RECT 1760.490 386.820 1760.810 386.880 ;
        RECT 1760.045 386.680 1760.810 386.820 ;
        RECT 1760.045 386.635 1760.335 386.680 ;
        RECT 1760.490 386.620 1760.810 386.680 ;
        RECT 1760.030 331.400 1760.350 331.460 ;
        RECT 1759.835 331.260 1760.350 331.400 ;
        RECT 1760.030 331.200 1760.350 331.260 ;
        RECT 1760.490 241.980 1760.810 242.040 ;
        RECT 1760.120 241.840 1760.810 241.980 ;
        RECT 1760.120 241.700 1760.260 241.840 ;
        RECT 1760.490 241.780 1760.810 241.840 ;
        RECT 1760.030 241.440 1760.350 241.700 ;
        RECT 1760.030 186.560 1760.350 186.620 ;
        RECT 1760.490 186.560 1760.810 186.620 ;
        RECT 1760.030 186.420 1760.810 186.560 ;
        RECT 1760.030 186.360 1760.350 186.420 ;
        RECT 1760.490 186.360 1760.810 186.420 ;
        RECT 1200.210 70.280 1200.530 70.340 ;
        RECT 1760.950 70.280 1761.270 70.340 ;
        RECT 1200.210 70.140 1761.270 70.280 ;
        RECT 1200.210 70.080 1200.530 70.140 ;
        RECT 1760.950 70.080 1761.270 70.140 ;
        RECT 1197.910 18.260 1198.230 18.320 ;
        RECT 1200.210 18.260 1200.530 18.320 ;
        RECT 1197.910 18.120 1200.530 18.260 ;
        RECT 1197.910 18.060 1198.230 18.120 ;
        RECT 1200.210 18.060 1200.530 18.120 ;
      LAYER via ;
        RECT 1760.060 1666.380 1760.320 1666.640 ;
        RECT 1763.280 1666.380 1763.540 1666.640 ;
        RECT 1760.520 1580.020 1760.780 1580.280 ;
        RECT 1761.440 1580.020 1761.700 1580.280 ;
        RECT 1760.520 1531.740 1760.780 1532.000 ;
        RECT 1761.440 1531.740 1761.700 1532.000 ;
        RECT 1760.520 1490.260 1760.780 1490.520 ;
        RECT 1760.520 1439.600 1760.780 1439.860 ;
        RECT 1760.520 1400.500 1760.780 1400.760 ;
        RECT 1761.440 1400.500 1761.700 1400.760 ;
        RECT 1759.140 1297.140 1759.400 1297.400 ;
        RECT 1760.060 1297.140 1760.320 1297.400 ;
        RECT 1760.060 1256.000 1760.320 1256.260 ;
        RECT 1760.520 1256.000 1760.780 1256.260 ;
        RECT 1759.140 1172.360 1759.400 1172.620 ;
        RECT 1760.520 1172.360 1760.780 1172.620 ;
        RECT 1759.140 1104.020 1759.400 1104.280 ;
        RECT 1760.060 1104.020 1760.320 1104.280 ;
        RECT 1760.060 1062.540 1760.320 1062.800 ;
        RECT 1760.520 1062.540 1760.780 1062.800 ;
        RECT 1759.140 1055.400 1759.400 1055.660 ;
        RECT 1760.060 1055.400 1760.320 1055.660 ;
        RECT 1760.520 1007.120 1760.780 1007.380 ;
        RECT 1760.520 965.640 1760.780 965.900 ;
        RECT 1760.060 917.700 1760.320 917.960 ;
        RECT 1760.980 917.700 1761.240 917.960 ;
        RECT 1760.060 903.760 1760.320 904.020 ;
        RECT 1760.520 814.340 1760.780 814.600 ;
        RECT 1760.060 724.240 1760.320 724.500 ;
        RECT 1760.980 724.240 1761.240 724.500 ;
        RECT 1759.140 475.360 1759.400 475.620 ;
        RECT 1760.980 475.360 1761.240 475.620 ;
        RECT 1760.520 427.760 1760.780 428.020 ;
        RECT 1760.980 427.760 1761.240 428.020 ;
        RECT 1760.520 386.620 1760.780 386.880 ;
        RECT 1760.060 331.200 1760.320 331.460 ;
        RECT 1760.520 241.780 1760.780 242.040 ;
        RECT 1760.060 241.440 1760.320 241.700 ;
        RECT 1760.060 186.360 1760.320 186.620 ;
        RECT 1760.520 186.360 1760.780 186.620 ;
        RECT 1200.240 70.080 1200.500 70.340 ;
        RECT 1760.980 70.080 1761.240 70.340 ;
        RECT 1197.940 18.060 1198.200 18.320 ;
        RECT 1200.240 18.060 1200.500 18.320 ;
      LAYER met2 ;
        RECT 1765.040 1700.410 1765.320 1704.000 ;
        RECT 1763.340 1700.270 1765.320 1700.410 ;
        RECT 1763.340 1666.670 1763.480 1700.270 ;
        RECT 1765.040 1700.000 1765.320 1700.270 ;
        RECT 1760.060 1666.350 1760.320 1666.670 ;
        RECT 1763.280 1666.350 1763.540 1666.670 ;
        RECT 1760.120 1642.610 1760.260 1666.350 ;
        RECT 1760.120 1642.470 1760.720 1642.610 ;
        RECT 1760.580 1628.445 1760.720 1642.470 ;
        RECT 1760.510 1628.075 1760.790 1628.445 ;
        RECT 1761.430 1628.075 1761.710 1628.445 ;
        RECT 1761.500 1580.310 1761.640 1628.075 ;
        RECT 1760.520 1580.165 1760.780 1580.310 ;
        RECT 1761.440 1580.165 1761.700 1580.310 ;
        RECT 1760.510 1579.795 1760.790 1580.165 ;
        RECT 1761.430 1579.795 1761.710 1580.165 ;
        RECT 1761.500 1532.030 1761.640 1579.795 ;
        RECT 1760.520 1531.710 1760.780 1532.030 ;
        RECT 1761.440 1531.710 1761.700 1532.030 ;
        RECT 1760.580 1490.550 1760.720 1531.710 ;
        RECT 1760.520 1490.230 1760.780 1490.550 ;
        RECT 1760.520 1439.570 1760.780 1439.890 ;
        RECT 1760.580 1435.325 1760.720 1439.570 ;
        RECT 1760.510 1434.955 1760.790 1435.325 ;
        RECT 1761.430 1434.955 1761.710 1435.325 ;
        RECT 1761.500 1400.790 1761.640 1434.955 ;
        RECT 1760.520 1400.470 1760.780 1400.790 ;
        RECT 1761.440 1400.470 1761.700 1400.790 ;
        RECT 1760.580 1345.565 1760.720 1400.470 ;
        RECT 1759.130 1345.195 1759.410 1345.565 ;
        RECT 1760.510 1345.195 1760.790 1345.565 ;
        RECT 1759.200 1297.430 1759.340 1345.195 ;
        RECT 1759.140 1297.110 1759.400 1297.430 ;
        RECT 1760.060 1297.110 1760.320 1297.430 ;
        RECT 1760.120 1256.290 1760.260 1297.110 ;
        RECT 1760.060 1255.970 1760.320 1256.290 ;
        RECT 1760.520 1255.970 1760.780 1256.290 ;
        RECT 1760.580 1231.890 1760.720 1255.970 ;
        RECT 1760.120 1231.750 1760.720 1231.890 ;
        RECT 1760.120 1200.725 1760.260 1231.750 ;
        RECT 1759.130 1200.355 1759.410 1200.725 ;
        RECT 1760.050 1200.355 1760.330 1200.725 ;
        RECT 1759.200 1172.650 1759.340 1200.355 ;
        RECT 1759.140 1172.330 1759.400 1172.650 ;
        RECT 1760.520 1172.330 1760.780 1172.650 ;
        RECT 1760.580 1152.445 1760.720 1172.330 ;
        RECT 1759.130 1152.075 1759.410 1152.445 ;
        RECT 1760.510 1152.075 1760.790 1152.445 ;
        RECT 1759.200 1104.310 1759.340 1152.075 ;
        RECT 1759.140 1103.990 1759.400 1104.310 ;
        RECT 1760.060 1103.990 1760.320 1104.310 ;
        RECT 1760.120 1062.830 1760.260 1103.990 ;
        RECT 1760.060 1062.570 1760.320 1062.830 ;
        RECT 1760.520 1062.570 1760.780 1062.830 ;
        RECT 1760.060 1062.510 1760.780 1062.570 ;
        RECT 1760.120 1062.430 1760.720 1062.510 ;
        RECT 1760.120 1055.690 1760.260 1062.430 ;
        RECT 1759.140 1055.370 1759.400 1055.690 ;
        RECT 1760.060 1055.370 1760.320 1055.690 ;
        RECT 1759.200 1007.605 1759.340 1055.370 ;
        RECT 1759.130 1007.235 1759.410 1007.605 ;
        RECT 1760.510 1007.235 1760.790 1007.605 ;
        RECT 1760.520 1007.090 1760.780 1007.235 ;
        RECT 1760.520 965.610 1760.780 965.930 ;
        RECT 1760.580 959.210 1760.720 965.610 ;
        RECT 1760.580 959.070 1761.180 959.210 ;
        RECT 1761.040 917.990 1761.180 959.070 ;
        RECT 1760.060 917.670 1760.320 917.990 ;
        RECT 1760.980 917.670 1761.240 917.990 ;
        RECT 1760.120 904.050 1760.260 917.670 ;
        RECT 1760.060 903.730 1760.320 904.050 ;
        RECT 1760.520 814.310 1760.780 814.630 ;
        RECT 1760.580 766.090 1760.720 814.310 ;
        RECT 1760.120 765.950 1760.720 766.090 ;
        RECT 1760.120 724.530 1760.260 765.950 ;
        RECT 1760.060 724.210 1760.320 724.530 ;
        RECT 1760.980 724.210 1761.240 724.530 ;
        RECT 1761.040 688.570 1761.180 724.210 ;
        RECT 1760.580 688.430 1761.180 688.570 ;
        RECT 1760.580 628.845 1760.720 688.430 ;
        RECT 1760.510 628.475 1760.790 628.845 ;
        RECT 1760.050 627.795 1760.330 628.165 ;
        RECT 1760.120 596.770 1760.260 627.795 ;
        RECT 1760.120 596.630 1760.720 596.770 ;
        RECT 1760.580 548.490 1760.720 596.630 ;
        RECT 1760.120 548.350 1760.720 548.490 ;
        RECT 1760.120 524.125 1760.260 548.350 ;
        RECT 1759.130 523.755 1759.410 524.125 ;
        RECT 1760.050 523.755 1760.330 524.125 ;
        RECT 1759.200 475.650 1759.340 523.755 ;
        RECT 1759.140 475.330 1759.400 475.650 ;
        RECT 1760.980 475.330 1761.240 475.650 ;
        RECT 1761.040 428.050 1761.180 475.330 ;
        RECT 1760.520 427.730 1760.780 428.050 ;
        RECT 1760.980 427.730 1761.240 428.050 ;
        RECT 1760.580 386.910 1760.720 427.730 ;
        RECT 1760.520 386.590 1760.780 386.910 ;
        RECT 1760.060 331.170 1760.320 331.490 ;
        RECT 1760.120 330.890 1760.260 331.170 ;
        RECT 1760.120 330.750 1760.720 330.890 ;
        RECT 1760.580 242.070 1760.720 330.750 ;
        RECT 1760.520 241.750 1760.780 242.070 ;
        RECT 1760.060 241.410 1760.320 241.730 ;
        RECT 1760.120 186.650 1760.260 241.410 ;
        RECT 1760.060 186.330 1760.320 186.650 ;
        RECT 1760.520 186.330 1760.780 186.650 ;
        RECT 1760.580 186.050 1760.720 186.330 ;
        RECT 1760.580 185.910 1761.640 186.050 ;
        RECT 1761.500 96.290 1761.640 185.910 ;
        RECT 1761.040 96.150 1761.640 96.290 ;
        RECT 1761.040 70.370 1761.180 96.150 ;
        RECT 1200.240 70.050 1200.500 70.370 ;
        RECT 1760.980 70.050 1761.240 70.370 ;
        RECT 1200.300 18.350 1200.440 70.050 ;
        RECT 1197.940 18.030 1198.200 18.350 ;
        RECT 1200.240 18.030 1200.500 18.350 ;
        RECT 1198.000 2.400 1198.140 18.030 ;
        RECT 1197.790 -4.800 1198.350 2.400 ;
      LAYER via2 ;
        RECT 1760.510 1628.120 1760.790 1628.400 ;
        RECT 1761.430 1628.120 1761.710 1628.400 ;
        RECT 1760.510 1579.840 1760.790 1580.120 ;
        RECT 1761.430 1579.840 1761.710 1580.120 ;
        RECT 1760.510 1435.000 1760.790 1435.280 ;
        RECT 1761.430 1435.000 1761.710 1435.280 ;
        RECT 1759.130 1345.240 1759.410 1345.520 ;
        RECT 1760.510 1345.240 1760.790 1345.520 ;
        RECT 1759.130 1200.400 1759.410 1200.680 ;
        RECT 1760.050 1200.400 1760.330 1200.680 ;
        RECT 1759.130 1152.120 1759.410 1152.400 ;
        RECT 1760.510 1152.120 1760.790 1152.400 ;
        RECT 1759.130 1007.280 1759.410 1007.560 ;
        RECT 1760.510 1007.280 1760.790 1007.560 ;
        RECT 1760.510 628.520 1760.790 628.800 ;
        RECT 1760.050 627.840 1760.330 628.120 ;
        RECT 1759.130 523.800 1759.410 524.080 ;
        RECT 1760.050 523.800 1760.330 524.080 ;
      LAYER met3 ;
        RECT 1760.485 1628.410 1760.815 1628.425 ;
        RECT 1761.405 1628.410 1761.735 1628.425 ;
        RECT 1760.485 1628.110 1761.735 1628.410 ;
        RECT 1760.485 1628.095 1760.815 1628.110 ;
        RECT 1761.405 1628.095 1761.735 1628.110 ;
        RECT 1760.485 1580.130 1760.815 1580.145 ;
        RECT 1761.405 1580.130 1761.735 1580.145 ;
        RECT 1760.485 1579.830 1761.735 1580.130 ;
        RECT 1760.485 1579.815 1760.815 1579.830 ;
        RECT 1761.405 1579.815 1761.735 1579.830 ;
        RECT 1760.485 1435.290 1760.815 1435.305 ;
        RECT 1761.405 1435.290 1761.735 1435.305 ;
        RECT 1760.485 1434.990 1761.735 1435.290 ;
        RECT 1760.485 1434.975 1760.815 1434.990 ;
        RECT 1761.405 1434.975 1761.735 1434.990 ;
        RECT 1759.105 1345.530 1759.435 1345.545 ;
        RECT 1760.485 1345.530 1760.815 1345.545 ;
        RECT 1759.105 1345.230 1760.815 1345.530 ;
        RECT 1759.105 1345.215 1759.435 1345.230 ;
        RECT 1760.485 1345.215 1760.815 1345.230 ;
        RECT 1759.105 1200.690 1759.435 1200.705 ;
        RECT 1760.025 1200.690 1760.355 1200.705 ;
        RECT 1759.105 1200.390 1760.355 1200.690 ;
        RECT 1759.105 1200.375 1759.435 1200.390 ;
        RECT 1760.025 1200.375 1760.355 1200.390 ;
        RECT 1759.105 1152.410 1759.435 1152.425 ;
        RECT 1760.485 1152.410 1760.815 1152.425 ;
        RECT 1759.105 1152.110 1760.815 1152.410 ;
        RECT 1759.105 1152.095 1759.435 1152.110 ;
        RECT 1760.485 1152.095 1760.815 1152.110 ;
        RECT 1759.105 1007.570 1759.435 1007.585 ;
        RECT 1760.485 1007.570 1760.815 1007.585 ;
        RECT 1759.105 1007.270 1760.815 1007.570 ;
        RECT 1759.105 1007.255 1759.435 1007.270 ;
        RECT 1760.485 1007.255 1760.815 1007.270 ;
        RECT 1760.485 628.810 1760.815 628.825 ;
        RECT 1760.270 628.495 1760.815 628.810 ;
        RECT 1760.270 628.145 1760.570 628.495 ;
        RECT 1760.025 627.830 1760.570 628.145 ;
        RECT 1760.025 627.815 1760.355 627.830 ;
        RECT 1759.105 524.090 1759.435 524.105 ;
        RECT 1760.025 524.090 1760.355 524.105 ;
        RECT 1759.105 523.790 1760.355 524.090 ;
        RECT 1759.105 523.775 1759.435 523.790 ;
        RECT 1760.025 523.775 1760.355 523.790 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1220.910 72.320 1221.230 72.380 ;
        RECT 1773.830 72.320 1774.150 72.380 ;
        RECT 1220.910 72.180 1774.150 72.320 ;
        RECT 1220.910 72.120 1221.230 72.180 ;
        RECT 1773.830 72.120 1774.150 72.180 ;
        RECT 1215.850 18.260 1216.170 18.320 ;
        RECT 1220.910 18.260 1221.230 18.320 ;
        RECT 1215.850 18.120 1221.230 18.260 ;
        RECT 1215.850 18.060 1216.170 18.120 ;
        RECT 1220.910 18.060 1221.230 18.120 ;
      LAYER via ;
        RECT 1220.940 72.120 1221.200 72.380 ;
        RECT 1773.860 72.120 1774.120 72.380 ;
        RECT 1215.880 18.060 1216.140 18.320 ;
        RECT 1220.940 18.060 1221.200 18.320 ;
      LAYER met2 ;
        RECT 1774.240 1700.410 1774.520 1704.000 ;
        RECT 1773.920 1700.270 1774.520 1700.410 ;
        RECT 1773.920 72.410 1774.060 1700.270 ;
        RECT 1774.240 1700.000 1774.520 1700.270 ;
        RECT 1220.940 72.090 1221.200 72.410 ;
        RECT 1773.860 72.090 1774.120 72.410 ;
        RECT 1221.000 18.350 1221.140 72.090 ;
        RECT 1215.880 18.030 1216.140 18.350 ;
        RECT 1220.940 18.030 1221.200 18.350 ;
        RECT 1215.940 2.400 1216.080 18.030 ;
        RECT 1215.730 -4.800 1216.290 2.400 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1233.790 49.540 1234.110 49.600 ;
        RECT 1781.190 49.540 1781.510 49.600 ;
        RECT 1233.790 49.400 1781.510 49.540 ;
        RECT 1233.790 49.340 1234.110 49.400 ;
        RECT 1781.190 49.340 1781.510 49.400 ;
      LAYER via ;
        RECT 1233.820 49.340 1234.080 49.600 ;
        RECT 1781.220 49.340 1781.480 49.600 ;
      LAYER met2 ;
        RECT 1783.440 1700.410 1783.720 1704.000 ;
        RECT 1781.280 1700.270 1783.720 1700.410 ;
        RECT 1781.280 49.630 1781.420 1700.270 ;
        RECT 1783.440 1700.000 1783.720 1700.270 ;
        RECT 1233.820 49.310 1234.080 49.630 ;
        RECT 1781.220 49.310 1781.480 49.630 ;
        RECT 1233.880 2.400 1234.020 49.310 ;
        RECT 1233.670 -4.800 1234.230 2.400 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1787.705 1587.205 1787.875 1635.315 ;
        RECT 1788.165 897.005 1788.335 932.195 ;
        RECT 1788.165 482.545 1788.335 531.335 ;
        RECT 1788.625 372.725 1788.795 420.835 ;
        RECT 1787.705 179.605 1787.875 207.315 ;
        RECT 1787.705 49.045 1787.875 131.155 ;
      LAYER mcon ;
        RECT 1787.705 1635.145 1787.875 1635.315 ;
        RECT 1788.165 932.025 1788.335 932.195 ;
        RECT 1788.165 531.165 1788.335 531.335 ;
        RECT 1788.625 420.665 1788.795 420.835 ;
        RECT 1787.705 207.145 1787.875 207.315 ;
        RECT 1787.705 130.985 1787.875 131.155 ;
      LAYER met1 ;
        RECT 1788.090 1678.140 1788.410 1678.200 ;
        RECT 1791.310 1678.140 1791.630 1678.200 ;
        RECT 1788.090 1678.000 1791.630 1678.140 ;
        RECT 1788.090 1677.940 1788.410 1678.000 ;
        RECT 1791.310 1677.940 1791.630 1678.000 ;
        RECT 1787.645 1635.300 1787.935 1635.345 ;
        RECT 1788.090 1635.300 1788.410 1635.360 ;
        RECT 1787.645 1635.160 1788.410 1635.300 ;
        RECT 1787.645 1635.115 1787.935 1635.160 ;
        RECT 1788.090 1635.100 1788.410 1635.160 ;
        RECT 1787.630 1587.360 1787.950 1587.420 ;
        RECT 1787.435 1587.220 1787.950 1587.360 ;
        RECT 1787.630 1587.160 1787.950 1587.220 ;
        RECT 1787.630 1531.940 1787.950 1532.000 ;
        RECT 1788.550 1531.940 1788.870 1532.000 ;
        RECT 1787.630 1531.800 1788.870 1531.940 ;
        RECT 1787.630 1531.740 1787.950 1531.800 ;
        RECT 1788.550 1531.740 1788.870 1531.800 ;
        RECT 1788.090 1393.900 1788.410 1393.960 ;
        RECT 1789.010 1393.900 1789.330 1393.960 ;
        RECT 1788.090 1393.760 1789.330 1393.900 ;
        RECT 1788.090 1393.700 1788.410 1393.760 ;
        RECT 1789.010 1393.700 1789.330 1393.760 ;
        RECT 1788.090 1366.500 1788.410 1366.760 ;
        RECT 1788.180 1366.080 1788.320 1366.500 ;
        RECT 1788.090 1365.820 1788.410 1366.080 ;
        RECT 1788.550 1173.240 1788.870 1173.300 ;
        RECT 1788.180 1173.100 1788.870 1173.240 ;
        RECT 1788.180 1172.960 1788.320 1173.100 ;
        RECT 1788.550 1173.040 1788.870 1173.100 ;
        RECT 1788.090 1172.700 1788.410 1172.960 ;
        RECT 1788.550 1076.680 1788.870 1076.740 ;
        RECT 1788.180 1076.540 1788.870 1076.680 ;
        RECT 1788.180 1076.400 1788.320 1076.540 ;
        RECT 1788.550 1076.480 1788.870 1076.540 ;
        RECT 1788.090 1076.140 1788.410 1076.400 ;
        RECT 1788.090 932.180 1788.410 932.240 ;
        RECT 1787.895 932.040 1788.410 932.180 ;
        RECT 1788.090 931.980 1788.410 932.040 ;
        RECT 1788.090 897.160 1788.410 897.220 ;
        RECT 1787.895 897.020 1788.410 897.160 ;
        RECT 1788.090 896.960 1788.410 897.020 ;
        RECT 1787.630 724.440 1787.950 724.500 ;
        RECT 1788.550 724.440 1788.870 724.500 ;
        RECT 1787.630 724.300 1788.870 724.440 ;
        RECT 1787.630 724.240 1787.950 724.300 ;
        RECT 1788.550 724.240 1788.870 724.300 ;
        RECT 1788.090 593.680 1788.410 593.940 ;
        RECT 1788.180 593.260 1788.320 593.680 ;
        RECT 1788.090 593.000 1788.410 593.260 ;
        RECT 1788.090 531.320 1788.410 531.380 ;
        RECT 1787.895 531.180 1788.410 531.320 ;
        RECT 1788.090 531.120 1788.410 531.180 ;
        RECT 1788.105 482.700 1788.395 482.745 ;
        RECT 1788.550 482.700 1788.870 482.760 ;
        RECT 1788.105 482.560 1788.870 482.700 ;
        RECT 1788.105 482.515 1788.395 482.560 ;
        RECT 1788.550 482.500 1788.870 482.560 ;
        RECT 1787.630 434.420 1787.950 434.480 ;
        RECT 1788.550 434.420 1788.870 434.480 ;
        RECT 1787.630 434.280 1788.870 434.420 ;
        RECT 1787.630 434.220 1787.950 434.280 ;
        RECT 1788.550 434.220 1788.870 434.280 ;
        RECT 1788.550 420.820 1788.870 420.880 ;
        RECT 1788.355 420.680 1788.870 420.820 ;
        RECT 1788.550 420.620 1788.870 420.680 ;
        RECT 1788.550 372.880 1788.870 372.940 ;
        RECT 1788.355 372.740 1788.870 372.880 ;
        RECT 1788.550 372.680 1788.870 372.740 ;
        RECT 1788.090 324.600 1788.410 324.660 ;
        RECT 1788.550 324.600 1788.870 324.660 ;
        RECT 1788.090 324.460 1788.870 324.600 ;
        RECT 1788.090 324.400 1788.410 324.460 ;
        RECT 1788.550 324.400 1788.870 324.460 ;
        RECT 1787.645 207.300 1787.935 207.345 ;
        RECT 1788.090 207.300 1788.410 207.360 ;
        RECT 1787.645 207.160 1788.410 207.300 ;
        RECT 1787.645 207.115 1787.935 207.160 ;
        RECT 1788.090 207.100 1788.410 207.160 ;
        RECT 1787.630 179.760 1787.950 179.820 ;
        RECT 1787.435 179.620 1787.950 179.760 ;
        RECT 1787.630 179.560 1787.950 179.620 ;
        RECT 1787.630 131.140 1787.950 131.200 ;
        RECT 1787.435 131.000 1787.950 131.140 ;
        RECT 1787.630 130.940 1787.950 131.000 ;
        RECT 1251.730 49.200 1252.050 49.260 ;
        RECT 1787.645 49.200 1787.935 49.245 ;
        RECT 1251.730 49.060 1787.935 49.200 ;
        RECT 1251.730 49.000 1252.050 49.060 ;
        RECT 1787.645 49.015 1787.935 49.060 ;
      LAYER via ;
        RECT 1788.120 1677.940 1788.380 1678.200 ;
        RECT 1791.340 1677.940 1791.600 1678.200 ;
        RECT 1788.120 1635.100 1788.380 1635.360 ;
        RECT 1787.660 1587.160 1787.920 1587.420 ;
        RECT 1787.660 1531.740 1787.920 1532.000 ;
        RECT 1788.580 1531.740 1788.840 1532.000 ;
        RECT 1788.120 1393.700 1788.380 1393.960 ;
        RECT 1789.040 1393.700 1789.300 1393.960 ;
        RECT 1788.120 1366.500 1788.380 1366.760 ;
        RECT 1788.120 1365.820 1788.380 1366.080 ;
        RECT 1788.580 1173.040 1788.840 1173.300 ;
        RECT 1788.120 1172.700 1788.380 1172.960 ;
        RECT 1788.580 1076.480 1788.840 1076.740 ;
        RECT 1788.120 1076.140 1788.380 1076.400 ;
        RECT 1788.120 931.980 1788.380 932.240 ;
        RECT 1788.120 896.960 1788.380 897.220 ;
        RECT 1787.660 724.240 1787.920 724.500 ;
        RECT 1788.580 724.240 1788.840 724.500 ;
        RECT 1788.120 593.680 1788.380 593.940 ;
        RECT 1788.120 593.000 1788.380 593.260 ;
        RECT 1788.120 531.120 1788.380 531.380 ;
        RECT 1788.580 482.500 1788.840 482.760 ;
        RECT 1787.660 434.220 1787.920 434.480 ;
        RECT 1788.580 434.220 1788.840 434.480 ;
        RECT 1788.580 420.620 1788.840 420.880 ;
        RECT 1788.580 372.680 1788.840 372.940 ;
        RECT 1788.120 324.400 1788.380 324.660 ;
        RECT 1788.580 324.400 1788.840 324.660 ;
        RECT 1788.120 207.100 1788.380 207.360 ;
        RECT 1787.660 179.560 1787.920 179.820 ;
        RECT 1787.660 130.940 1787.920 131.200 ;
        RECT 1251.760 49.000 1252.020 49.260 ;
      LAYER met2 ;
        RECT 1792.640 1700.410 1792.920 1704.000 ;
        RECT 1791.400 1700.270 1792.920 1700.410 ;
        RECT 1791.400 1678.230 1791.540 1700.270 ;
        RECT 1792.640 1700.000 1792.920 1700.270 ;
        RECT 1788.120 1677.910 1788.380 1678.230 ;
        RECT 1791.340 1677.910 1791.600 1678.230 ;
        RECT 1788.180 1635.390 1788.320 1677.910 ;
        RECT 1788.120 1635.070 1788.380 1635.390 ;
        RECT 1787.660 1587.130 1787.920 1587.450 ;
        RECT 1787.720 1580.165 1787.860 1587.130 ;
        RECT 1787.650 1579.795 1787.930 1580.165 ;
        RECT 1788.570 1579.795 1788.850 1580.165 ;
        RECT 1788.640 1532.030 1788.780 1579.795 ;
        RECT 1787.660 1531.710 1787.920 1532.030 ;
        RECT 1788.580 1531.710 1788.840 1532.030 ;
        RECT 1787.720 1496.410 1787.860 1531.710 ;
        RECT 1787.720 1496.270 1788.320 1496.410 ;
        RECT 1788.180 1490.290 1788.320 1496.270 ;
        RECT 1787.720 1490.150 1788.320 1490.290 ;
        RECT 1787.720 1483.605 1787.860 1490.150 ;
        RECT 1787.650 1483.235 1787.930 1483.605 ;
        RECT 1789.030 1483.235 1789.310 1483.605 ;
        RECT 1789.100 1393.990 1789.240 1483.235 ;
        RECT 1788.120 1393.670 1788.380 1393.990 ;
        RECT 1789.040 1393.670 1789.300 1393.990 ;
        RECT 1788.180 1366.790 1788.320 1393.670 ;
        RECT 1788.120 1366.470 1788.380 1366.790 ;
        RECT 1788.120 1365.790 1788.380 1366.110 ;
        RECT 1788.180 1269.970 1788.320 1365.790 ;
        RECT 1787.720 1269.830 1788.320 1269.970 ;
        RECT 1787.720 1269.290 1787.860 1269.830 ;
        RECT 1787.720 1269.150 1788.320 1269.290 ;
        RECT 1788.180 1207.410 1788.320 1269.150 ;
        RECT 1788.180 1207.270 1788.780 1207.410 ;
        RECT 1788.640 1173.330 1788.780 1207.270 ;
        RECT 1788.580 1173.010 1788.840 1173.330 ;
        RECT 1788.120 1172.670 1788.380 1172.990 ;
        RECT 1788.180 1110.850 1788.320 1172.670 ;
        RECT 1788.180 1110.710 1788.780 1110.850 ;
        RECT 1788.640 1076.770 1788.780 1110.710 ;
        RECT 1788.580 1076.450 1788.840 1076.770 ;
        RECT 1788.120 1076.110 1788.380 1076.430 ;
        RECT 1788.180 980.290 1788.320 1076.110 ;
        RECT 1787.720 980.150 1788.320 980.290 ;
        RECT 1787.720 979.610 1787.860 980.150 ;
        RECT 1787.720 979.470 1788.320 979.610 ;
        RECT 1788.180 932.270 1788.320 979.470 ;
        RECT 1788.120 931.950 1788.380 932.270 ;
        RECT 1788.120 896.930 1788.380 897.250 ;
        RECT 1788.180 896.650 1788.320 896.930 ;
        RECT 1788.180 896.510 1788.780 896.650 ;
        RECT 1788.640 724.725 1788.780 896.510 ;
        RECT 1787.650 724.355 1787.930 724.725 ;
        RECT 1788.570 724.355 1788.850 724.725 ;
        RECT 1787.660 724.210 1787.920 724.355 ;
        RECT 1788.580 724.210 1788.840 724.355 ;
        RECT 1788.640 688.570 1788.780 724.210 ;
        RECT 1788.180 688.430 1788.780 688.570 ;
        RECT 1788.180 628.845 1788.320 688.430 ;
        RECT 1788.110 628.475 1788.390 628.845 ;
        RECT 1788.110 627.795 1788.390 628.165 ;
        RECT 1788.180 593.970 1788.320 627.795 ;
        RECT 1788.120 593.650 1788.380 593.970 ;
        RECT 1788.120 592.970 1788.380 593.290 ;
        RECT 1788.180 531.410 1788.320 592.970 ;
        RECT 1788.120 531.090 1788.380 531.410 ;
        RECT 1788.580 482.470 1788.840 482.790 ;
        RECT 1788.640 435.045 1788.780 482.470 ;
        RECT 1787.650 434.675 1787.930 435.045 ;
        RECT 1788.570 434.675 1788.850 435.045 ;
        RECT 1787.720 434.510 1787.860 434.675 ;
        RECT 1787.660 434.190 1787.920 434.510 ;
        RECT 1788.580 434.190 1788.840 434.510 ;
        RECT 1788.640 420.910 1788.780 434.190 ;
        RECT 1788.580 420.590 1788.840 420.910 ;
        RECT 1788.580 372.650 1788.840 372.970 ;
        RECT 1788.640 324.690 1788.780 372.650 ;
        RECT 1788.120 324.370 1788.380 324.690 ;
        RECT 1788.580 324.370 1788.840 324.690 ;
        RECT 1788.180 207.390 1788.320 324.370 ;
        RECT 1788.120 207.070 1788.380 207.390 ;
        RECT 1787.660 179.530 1787.920 179.850 ;
        RECT 1787.720 131.230 1787.860 179.530 ;
        RECT 1787.660 130.910 1787.920 131.230 ;
        RECT 1251.760 48.970 1252.020 49.290 ;
        RECT 1251.820 2.400 1251.960 48.970 ;
        RECT 1251.610 -4.800 1252.170 2.400 ;
      LAYER via2 ;
        RECT 1787.650 1579.840 1787.930 1580.120 ;
        RECT 1788.570 1579.840 1788.850 1580.120 ;
        RECT 1787.650 1483.280 1787.930 1483.560 ;
        RECT 1789.030 1483.280 1789.310 1483.560 ;
        RECT 1787.650 724.400 1787.930 724.680 ;
        RECT 1788.570 724.400 1788.850 724.680 ;
        RECT 1788.110 628.520 1788.390 628.800 ;
        RECT 1788.110 627.840 1788.390 628.120 ;
        RECT 1787.650 434.720 1787.930 435.000 ;
        RECT 1788.570 434.720 1788.850 435.000 ;
      LAYER met3 ;
        RECT 1787.625 1580.130 1787.955 1580.145 ;
        RECT 1788.545 1580.130 1788.875 1580.145 ;
        RECT 1787.625 1579.830 1788.875 1580.130 ;
        RECT 1787.625 1579.815 1787.955 1579.830 ;
        RECT 1788.545 1579.815 1788.875 1579.830 ;
        RECT 1787.625 1483.570 1787.955 1483.585 ;
        RECT 1789.005 1483.570 1789.335 1483.585 ;
        RECT 1787.625 1483.270 1789.335 1483.570 ;
        RECT 1787.625 1483.255 1787.955 1483.270 ;
        RECT 1789.005 1483.255 1789.335 1483.270 ;
        RECT 1787.625 724.690 1787.955 724.705 ;
        RECT 1788.545 724.690 1788.875 724.705 ;
        RECT 1787.625 724.390 1788.875 724.690 ;
        RECT 1787.625 724.375 1787.955 724.390 ;
        RECT 1788.545 724.375 1788.875 724.390 ;
        RECT 1788.085 628.810 1788.415 628.825 ;
        RECT 1787.870 628.495 1788.415 628.810 ;
        RECT 1787.870 628.145 1788.170 628.495 ;
        RECT 1787.870 627.830 1788.415 628.145 ;
        RECT 1788.085 627.815 1788.415 627.830 ;
        RECT 1787.625 435.010 1787.955 435.025 ;
        RECT 1788.545 435.010 1788.875 435.025 ;
        RECT 1787.625 434.710 1788.875 435.010 ;
        RECT 1787.625 434.695 1787.955 434.710 ;
        RECT 1788.545 434.695 1788.875 434.710 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1269.210 48.860 1269.530 48.920 ;
        RECT 1801.430 48.860 1801.750 48.920 ;
        RECT 1269.210 48.720 1801.750 48.860 ;
        RECT 1269.210 48.660 1269.530 48.720 ;
        RECT 1801.430 48.660 1801.750 48.720 ;
      LAYER via ;
        RECT 1269.240 48.660 1269.500 48.920 ;
        RECT 1801.460 48.660 1801.720 48.920 ;
      LAYER met2 ;
        RECT 1801.840 1700.410 1802.120 1704.000 ;
        RECT 1801.520 1700.270 1802.120 1700.410 ;
        RECT 1801.520 48.950 1801.660 1700.270 ;
        RECT 1801.840 1700.000 1802.120 1700.270 ;
        RECT 1269.240 48.630 1269.500 48.950 ;
        RECT 1801.460 48.630 1801.720 48.950 ;
        RECT 1269.300 2.400 1269.440 48.630 ;
        RECT 1269.090 -4.800 1269.650 2.400 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1287.150 48.520 1287.470 48.580 ;
        RECT 1808.790 48.520 1809.110 48.580 ;
        RECT 1287.150 48.380 1809.110 48.520 ;
        RECT 1287.150 48.320 1287.470 48.380 ;
        RECT 1808.790 48.320 1809.110 48.380 ;
      LAYER via ;
        RECT 1287.180 48.320 1287.440 48.580 ;
        RECT 1808.820 48.320 1809.080 48.580 ;
      LAYER met2 ;
        RECT 1811.040 1700.410 1811.320 1704.000 ;
        RECT 1808.880 1700.270 1811.320 1700.410 ;
        RECT 1808.880 48.610 1809.020 1700.270 ;
        RECT 1811.040 1700.000 1811.320 1700.270 ;
        RECT 1287.180 48.290 1287.440 48.610 ;
        RECT 1808.820 48.290 1809.080 48.610 ;
        RECT 1287.240 2.400 1287.380 48.290 ;
        RECT 1287.030 -4.800 1287.590 2.400 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1814.770 1678.140 1815.090 1678.200 ;
        RECT 1818.910 1678.140 1819.230 1678.200 ;
        RECT 1814.770 1678.000 1819.230 1678.140 ;
        RECT 1814.770 1677.940 1815.090 1678.000 ;
        RECT 1818.910 1677.940 1819.230 1678.000 ;
        RECT 1780.270 23.020 1780.590 23.080 ;
        RECT 1814.770 23.020 1815.090 23.080 ;
        RECT 1780.270 22.880 1815.090 23.020 ;
        RECT 1780.270 22.820 1780.590 22.880 ;
        RECT 1814.770 22.820 1815.090 22.880 ;
        RECT 1305.090 17.240 1305.410 17.300 ;
        RECT 1780.270 17.240 1780.590 17.300 ;
        RECT 1305.090 17.100 1780.590 17.240 ;
        RECT 1305.090 17.040 1305.410 17.100 ;
        RECT 1780.270 17.040 1780.590 17.100 ;
      LAYER via ;
        RECT 1814.800 1677.940 1815.060 1678.200 ;
        RECT 1818.940 1677.940 1819.200 1678.200 ;
        RECT 1780.300 22.820 1780.560 23.080 ;
        RECT 1814.800 22.820 1815.060 23.080 ;
        RECT 1305.120 17.040 1305.380 17.300 ;
        RECT 1780.300 17.040 1780.560 17.300 ;
      LAYER met2 ;
        RECT 1820.240 1700.410 1820.520 1704.000 ;
        RECT 1819.000 1700.270 1820.520 1700.410 ;
        RECT 1819.000 1678.230 1819.140 1700.270 ;
        RECT 1820.240 1700.000 1820.520 1700.270 ;
        RECT 1814.800 1677.910 1815.060 1678.230 ;
        RECT 1818.940 1677.910 1819.200 1678.230 ;
        RECT 1814.860 23.110 1815.000 1677.910 ;
        RECT 1780.300 22.790 1780.560 23.110 ;
        RECT 1814.800 22.790 1815.060 23.110 ;
        RECT 1780.360 17.330 1780.500 22.790 ;
        RECT 1305.120 17.010 1305.380 17.330 ;
        RECT 1780.300 17.010 1780.560 17.330 ;
        RECT 1305.180 2.400 1305.320 17.010 ;
        RECT 1304.970 -4.800 1305.530 2.400 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1410.505 20.145 1411.595 20.315 ;
        RECT 1410.505 18.445 1410.675 20.145 ;
        RECT 1411.425 19.805 1411.595 20.145 ;
      LAYER met1 ;
        RECT 1417.790 1688.340 1418.110 1688.400 ;
        RECT 1829.490 1688.340 1829.810 1688.400 ;
        RECT 1417.790 1688.200 1829.810 1688.340 ;
        RECT 1417.790 1688.140 1418.110 1688.200 ;
        RECT 1829.490 1688.140 1829.810 1688.200 ;
        RECT 1411.365 19.960 1411.655 20.005 ;
        RECT 1417.330 19.960 1417.650 20.020 ;
        RECT 1411.365 19.820 1417.650 19.960 ;
        RECT 1411.365 19.775 1411.655 19.820 ;
        RECT 1417.330 19.760 1417.650 19.820 ;
        RECT 1323.030 18.600 1323.350 18.660 ;
        RECT 1410.445 18.600 1410.735 18.645 ;
        RECT 1323.030 18.460 1410.735 18.600 ;
        RECT 1323.030 18.400 1323.350 18.460 ;
        RECT 1410.445 18.415 1410.735 18.460 ;
      LAYER via ;
        RECT 1417.820 1688.140 1418.080 1688.400 ;
        RECT 1829.520 1688.140 1829.780 1688.400 ;
        RECT 1417.360 19.760 1417.620 20.020 ;
        RECT 1323.060 18.400 1323.320 18.660 ;
      LAYER met2 ;
        RECT 1829.440 1700.000 1829.720 1704.000 ;
        RECT 1829.580 1688.430 1829.720 1700.000 ;
        RECT 1417.820 1688.110 1418.080 1688.430 ;
        RECT 1829.520 1688.110 1829.780 1688.430 ;
        RECT 1417.880 40.530 1418.020 1688.110 ;
        RECT 1417.420 40.390 1418.020 40.530 ;
        RECT 1417.420 20.050 1417.560 40.390 ;
        RECT 1417.360 19.730 1417.620 20.050 ;
        RECT 1323.060 18.370 1323.320 18.690 ;
        RECT 1323.120 2.400 1323.260 18.370 ;
        RECT 1322.910 -4.800 1323.470 2.400 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1383.825 16.745 1383.995 17.935 ;
      LAYER mcon ;
        RECT 1383.825 17.765 1383.995 17.935 ;
      LAYER met1 ;
        RECT 1449.530 53.280 1449.850 53.340 ;
        RECT 1835.930 53.280 1836.250 53.340 ;
        RECT 1449.530 53.140 1836.250 53.280 ;
        RECT 1449.530 53.080 1449.850 53.140 ;
        RECT 1835.930 53.080 1836.250 53.140 ;
        RECT 1383.765 17.920 1384.055 17.965 ;
        RECT 1383.765 17.780 1438.720 17.920 ;
        RECT 1383.765 17.735 1384.055 17.780 ;
        RECT 1438.580 17.580 1438.720 17.780 ;
        RECT 1449.530 17.580 1449.850 17.640 ;
        RECT 1438.580 17.440 1449.850 17.580 ;
        RECT 1449.530 17.380 1449.850 17.440 ;
        RECT 1340.510 16.900 1340.830 16.960 ;
        RECT 1383.765 16.900 1384.055 16.945 ;
        RECT 1340.510 16.760 1384.055 16.900 ;
        RECT 1340.510 16.700 1340.830 16.760 ;
        RECT 1383.765 16.715 1384.055 16.760 ;
      LAYER via ;
        RECT 1449.560 53.080 1449.820 53.340 ;
        RECT 1835.960 53.080 1836.220 53.340 ;
        RECT 1449.560 17.380 1449.820 17.640 ;
        RECT 1340.540 16.700 1340.800 16.960 ;
      LAYER met2 ;
        RECT 1838.640 1700.410 1838.920 1704.000 ;
        RECT 1836.020 1700.270 1838.920 1700.410 ;
        RECT 1836.020 53.370 1836.160 1700.270 ;
        RECT 1838.640 1700.000 1838.920 1700.270 ;
        RECT 1449.560 53.050 1449.820 53.370 ;
        RECT 1835.960 53.050 1836.220 53.370 ;
        RECT 1449.620 17.670 1449.760 53.050 ;
        RECT 1449.560 17.350 1449.820 17.670 ;
        RECT 1340.540 16.670 1340.800 16.990 ;
        RECT 1340.600 2.400 1340.740 16.670 ;
        RECT 1340.390 -4.800 1340.950 2.400 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 703.410 54.640 703.730 54.700 ;
        RECT 1505.190 54.640 1505.510 54.700 ;
        RECT 703.410 54.500 1505.510 54.640 ;
        RECT 703.410 54.440 703.730 54.500 ;
        RECT 1505.190 54.440 1505.510 54.500 ;
        RECT 698.350 2.960 698.670 3.020 ;
        RECT 703.410 2.960 703.730 3.020 ;
        RECT 698.350 2.820 703.730 2.960 ;
        RECT 698.350 2.760 698.670 2.820 ;
        RECT 703.410 2.760 703.730 2.820 ;
      LAYER via ;
        RECT 703.440 54.440 703.700 54.700 ;
        RECT 1505.220 54.440 1505.480 54.700 ;
        RECT 698.380 2.760 698.640 3.020 ;
        RECT 703.440 2.760 703.700 3.020 ;
      LAYER met2 ;
        RECT 1507.900 1700.410 1508.180 1704.000 ;
        RECT 1505.280 1700.270 1508.180 1700.410 ;
        RECT 1505.280 54.730 1505.420 1700.270 ;
        RECT 1507.900 1700.000 1508.180 1700.270 ;
        RECT 703.440 54.410 703.700 54.730 ;
        RECT 1505.220 54.410 1505.480 54.730 ;
        RECT 703.500 3.050 703.640 54.410 ;
        RECT 698.380 2.730 698.640 3.050 ;
        RECT 703.440 2.730 703.700 3.050 ;
        RECT 698.440 2.400 698.580 2.730 ;
        RECT 698.230 -4.800 698.790 2.400 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1410.965 18.445 1411.135 19.975 ;
      LAYER mcon ;
        RECT 1410.965 19.805 1411.135 19.975 ;
      LAYER met1 ;
        RECT 1438.490 1688.680 1438.810 1688.740 ;
        RECT 1847.890 1688.680 1848.210 1688.740 ;
        RECT 1438.490 1688.540 1848.210 1688.680 ;
        RECT 1438.490 1688.480 1438.810 1688.540 ;
        RECT 1847.890 1688.480 1848.210 1688.540 ;
        RECT 1358.450 19.960 1358.770 20.020 ;
        RECT 1410.905 19.960 1411.195 20.005 ;
        RECT 1358.450 19.820 1411.195 19.960 ;
        RECT 1358.450 19.760 1358.770 19.820 ;
        RECT 1410.905 19.775 1411.195 19.820 ;
        RECT 1410.905 18.600 1411.195 18.645 ;
        RECT 1438.490 18.600 1438.810 18.660 ;
        RECT 1410.905 18.460 1438.810 18.600 ;
        RECT 1410.905 18.415 1411.195 18.460 ;
        RECT 1438.490 18.400 1438.810 18.460 ;
      LAYER via ;
        RECT 1438.520 1688.480 1438.780 1688.740 ;
        RECT 1847.920 1688.480 1848.180 1688.740 ;
        RECT 1358.480 19.760 1358.740 20.020 ;
        RECT 1438.520 18.400 1438.780 18.660 ;
      LAYER met2 ;
        RECT 1847.840 1700.000 1848.120 1704.000 ;
        RECT 1847.980 1688.770 1848.120 1700.000 ;
        RECT 1438.520 1688.450 1438.780 1688.770 ;
        RECT 1847.920 1688.450 1848.180 1688.770 ;
        RECT 1358.480 19.730 1358.740 20.050 ;
        RECT 1358.540 2.400 1358.680 19.730 ;
        RECT 1438.580 18.690 1438.720 1688.450 ;
        RECT 1438.520 18.370 1438.780 18.690 ;
        RECT 1358.330 -4.800 1358.890 2.400 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1383.290 1686.980 1383.610 1687.040 ;
        RECT 1857.090 1686.980 1857.410 1687.040 ;
        RECT 1383.290 1686.840 1857.410 1686.980 ;
        RECT 1383.290 1686.780 1383.610 1686.840 ;
        RECT 1857.090 1686.780 1857.410 1686.840 ;
        RECT 1376.390 17.920 1376.710 17.980 ;
        RECT 1383.290 17.920 1383.610 17.980 ;
        RECT 1376.390 17.780 1383.610 17.920 ;
        RECT 1376.390 17.720 1376.710 17.780 ;
        RECT 1383.290 17.720 1383.610 17.780 ;
      LAYER via ;
        RECT 1383.320 1686.780 1383.580 1687.040 ;
        RECT 1857.120 1686.780 1857.380 1687.040 ;
        RECT 1376.420 17.720 1376.680 17.980 ;
        RECT 1383.320 17.720 1383.580 17.980 ;
      LAYER met2 ;
        RECT 1857.040 1700.000 1857.320 1704.000 ;
        RECT 1857.180 1687.070 1857.320 1700.000 ;
        RECT 1383.320 1686.750 1383.580 1687.070 ;
        RECT 1857.120 1686.750 1857.380 1687.070 ;
        RECT 1383.380 18.010 1383.520 1686.750 ;
        RECT 1376.420 17.690 1376.680 18.010 ;
        RECT 1383.320 17.690 1383.580 18.010 ;
        RECT 1376.480 2.400 1376.620 17.690 ;
        RECT 1376.270 -4.800 1376.830 2.400 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1400.310 1687.320 1400.630 1687.380 ;
        RECT 1866.290 1687.320 1866.610 1687.380 ;
        RECT 1400.310 1687.180 1866.610 1687.320 ;
        RECT 1400.310 1687.120 1400.630 1687.180 ;
        RECT 1866.290 1687.120 1866.610 1687.180 ;
        RECT 1394.330 16.900 1394.650 16.960 ;
        RECT 1400.310 16.900 1400.630 16.960 ;
        RECT 1394.330 16.760 1400.630 16.900 ;
        RECT 1394.330 16.700 1394.650 16.760 ;
        RECT 1400.310 16.700 1400.630 16.760 ;
      LAYER via ;
        RECT 1400.340 1687.120 1400.600 1687.380 ;
        RECT 1866.320 1687.120 1866.580 1687.380 ;
        RECT 1394.360 16.700 1394.620 16.960 ;
        RECT 1400.340 16.700 1400.600 16.960 ;
      LAYER met2 ;
        RECT 1866.240 1700.000 1866.520 1704.000 ;
        RECT 1866.380 1687.410 1866.520 1700.000 ;
        RECT 1400.340 1687.090 1400.600 1687.410 ;
        RECT 1866.320 1687.090 1866.580 1687.410 ;
        RECT 1400.400 16.990 1400.540 1687.090 ;
        RECT 1394.360 16.670 1394.620 16.990 ;
        RECT 1400.340 16.670 1400.600 16.990 ;
        RECT 1394.420 2.400 1394.560 16.670 ;
        RECT 1394.210 -4.800 1394.770 2.400 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1472.990 1689.020 1473.310 1689.080 ;
        RECT 1875.490 1689.020 1875.810 1689.080 ;
        RECT 1472.990 1688.880 1875.810 1689.020 ;
        RECT 1472.990 1688.820 1473.310 1688.880 ;
        RECT 1875.490 1688.820 1875.810 1688.880 ;
        RECT 1412.270 16.900 1412.590 16.960 ;
        RECT 1472.990 16.900 1473.310 16.960 ;
        RECT 1412.270 16.760 1473.310 16.900 ;
        RECT 1412.270 16.700 1412.590 16.760 ;
        RECT 1472.990 16.700 1473.310 16.760 ;
      LAYER via ;
        RECT 1473.020 1688.820 1473.280 1689.080 ;
        RECT 1875.520 1688.820 1875.780 1689.080 ;
        RECT 1412.300 16.700 1412.560 16.960 ;
        RECT 1473.020 16.700 1473.280 16.960 ;
      LAYER met2 ;
        RECT 1875.440 1700.000 1875.720 1704.000 ;
        RECT 1875.580 1689.110 1875.720 1700.000 ;
        RECT 1473.020 1688.790 1473.280 1689.110 ;
        RECT 1875.520 1688.790 1875.780 1689.110 ;
        RECT 1473.080 16.990 1473.220 1688.790 ;
        RECT 1412.300 16.670 1412.560 16.990 ;
        RECT 1473.020 16.670 1473.280 16.990 ;
        RECT 1412.360 2.400 1412.500 16.670 ;
        RECT 1412.150 -4.800 1412.710 2.400 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1434.810 1687.660 1435.130 1687.720 ;
        RECT 1884.690 1687.660 1885.010 1687.720 ;
        RECT 1434.810 1687.520 1885.010 1687.660 ;
        RECT 1434.810 1687.460 1435.130 1687.520 ;
        RECT 1884.690 1687.460 1885.010 1687.520 ;
        RECT 1429.750 15.880 1430.070 15.940 ;
        RECT 1434.810 15.880 1435.130 15.940 ;
        RECT 1429.750 15.740 1435.130 15.880 ;
        RECT 1429.750 15.680 1430.070 15.740 ;
        RECT 1434.810 15.680 1435.130 15.740 ;
      LAYER via ;
        RECT 1434.840 1687.460 1435.100 1687.720 ;
        RECT 1884.720 1687.460 1884.980 1687.720 ;
        RECT 1429.780 15.680 1430.040 15.940 ;
        RECT 1434.840 15.680 1435.100 15.940 ;
      LAYER met2 ;
        RECT 1884.640 1700.000 1884.920 1704.000 ;
        RECT 1884.780 1687.750 1884.920 1700.000 ;
        RECT 1434.840 1687.430 1435.100 1687.750 ;
        RECT 1884.720 1687.430 1884.980 1687.750 ;
        RECT 1434.900 15.970 1435.040 1687.430 ;
        RECT 1429.780 15.650 1430.040 15.970 ;
        RECT 1434.840 15.650 1435.100 15.970 ;
        RECT 1429.840 2.400 1429.980 15.650 ;
        RECT 1429.630 -4.800 1430.190 2.400 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1462.945 16.405 1463.115 17.935 ;
        RECT 1510.785 16.405 1510.955 17.595 ;
        RECT 1864.065 17.425 1864.235 18.615 ;
      LAYER mcon ;
        RECT 1864.065 18.445 1864.235 18.615 ;
        RECT 1462.945 17.765 1463.115 17.935 ;
        RECT 1510.785 17.425 1510.955 17.595 ;
      LAYER met1 ;
        RECT 1864.005 18.600 1864.295 18.645 ;
        RECT 1892.050 18.600 1892.370 18.660 ;
        RECT 1864.005 18.460 1892.370 18.600 ;
        RECT 1864.005 18.415 1864.295 18.460 ;
        RECT 1892.050 18.400 1892.370 18.460 ;
        RECT 1447.690 17.920 1448.010 17.980 ;
        RECT 1462.885 17.920 1463.175 17.965 ;
        RECT 1447.690 17.780 1463.175 17.920 ;
        RECT 1447.690 17.720 1448.010 17.780 ;
        RECT 1462.885 17.735 1463.175 17.780 ;
        RECT 1510.725 17.580 1511.015 17.625 ;
        RECT 1864.005 17.580 1864.295 17.625 ;
        RECT 1510.725 17.440 1864.295 17.580 ;
        RECT 1510.725 17.395 1511.015 17.440 ;
        RECT 1864.005 17.395 1864.295 17.440 ;
        RECT 1462.885 16.560 1463.175 16.605 ;
        RECT 1510.725 16.560 1511.015 16.605 ;
        RECT 1462.885 16.420 1511.015 16.560 ;
        RECT 1462.885 16.375 1463.175 16.420 ;
        RECT 1510.725 16.375 1511.015 16.420 ;
      LAYER via ;
        RECT 1892.080 18.400 1892.340 18.660 ;
        RECT 1447.720 17.720 1447.980 17.980 ;
      LAYER met2 ;
        RECT 1893.840 1700.410 1894.120 1704.000 ;
        RECT 1892.140 1700.270 1894.120 1700.410 ;
        RECT 1892.140 18.690 1892.280 1700.270 ;
        RECT 1893.840 1700.000 1894.120 1700.270 ;
        RECT 1892.080 18.370 1892.340 18.690 ;
        RECT 1447.720 17.690 1447.980 18.010 ;
        RECT 1447.780 2.400 1447.920 17.690 ;
        RECT 1447.570 -4.800 1448.130 2.400 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1469.310 1688.000 1469.630 1688.060 ;
        RECT 1903.090 1688.000 1903.410 1688.060 ;
        RECT 1469.310 1687.860 1903.410 1688.000 ;
        RECT 1469.310 1687.800 1469.630 1687.860 ;
        RECT 1903.090 1687.800 1903.410 1687.860 ;
        RECT 1465.630 15.880 1465.950 15.940 ;
        RECT 1469.310 15.880 1469.630 15.940 ;
        RECT 1465.630 15.740 1469.630 15.880 ;
        RECT 1465.630 15.680 1465.950 15.740 ;
        RECT 1469.310 15.680 1469.630 15.740 ;
      LAYER via ;
        RECT 1469.340 1687.800 1469.600 1688.060 ;
        RECT 1903.120 1687.800 1903.380 1688.060 ;
        RECT 1465.660 15.680 1465.920 15.940 ;
        RECT 1469.340 15.680 1469.600 15.940 ;
      LAYER met2 ;
        RECT 1903.040 1700.000 1903.320 1704.000 ;
        RECT 1903.180 1688.090 1903.320 1700.000 ;
        RECT 1469.340 1687.770 1469.600 1688.090 ;
        RECT 1903.120 1687.770 1903.380 1688.090 ;
        RECT 1469.400 15.970 1469.540 1687.770 ;
        RECT 1465.660 15.650 1465.920 15.970 ;
        RECT 1469.340 15.650 1469.600 15.970 ;
        RECT 1465.720 2.400 1465.860 15.650 ;
        RECT 1465.510 -4.800 1466.070 2.400 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1907.690 1683.920 1908.010 1683.980 ;
        RECT 1912.290 1683.920 1912.610 1683.980 ;
        RECT 1907.690 1683.780 1912.610 1683.920 ;
        RECT 1907.690 1683.720 1908.010 1683.780 ;
        RECT 1912.290 1683.720 1912.610 1683.780 ;
        RECT 1483.570 17.920 1483.890 17.980 ;
        RECT 1907.690 17.920 1908.010 17.980 ;
        RECT 1483.570 17.780 1908.010 17.920 ;
        RECT 1483.570 17.720 1483.890 17.780 ;
        RECT 1907.690 17.720 1908.010 17.780 ;
      LAYER via ;
        RECT 1907.720 1683.720 1907.980 1683.980 ;
        RECT 1912.320 1683.720 1912.580 1683.980 ;
        RECT 1483.600 17.720 1483.860 17.980 ;
        RECT 1907.720 17.720 1907.980 17.980 ;
      LAYER met2 ;
        RECT 1912.240 1700.000 1912.520 1704.000 ;
        RECT 1912.380 1684.010 1912.520 1700.000 ;
        RECT 1907.720 1683.690 1907.980 1684.010 ;
        RECT 1912.320 1683.690 1912.580 1684.010 ;
        RECT 1907.780 18.010 1907.920 1683.690 ;
        RECT 1483.600 17.690 1483.860 18.010 ;
        RECT 1907.720 17.690 1907.980 18.010 ;
        RECT 1483.660 2.400 1483.800 17.690 ;
        RECT 1483.450 -4.800 1484.010 2.400 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1885.225 1683.765 1885.395 1687.675 ;
      LAYER mcon ;
        RECT 1885.225 1687.505 1885.395 1687.675 ;
      LAYER met1 ;
        RECT 1885.165 1687.660 1885.455 1687.705 ;
        RECT 1920.110 1687.660 1920.430 1687.720 ;
        RECT 1885.165 1687.520 1920.430 1687.660 ;
        RECT 1885.165 1687.475 1885.455 1687.520 ;
        RECT 1920.110 1687.460 1920.430 1687.520 ;
        RECT 1818.450 1683.920 1818.770 1683.980 ;
        RECT 1885.165 1683.920 1885.455 1683.965 ;
        RECT 1818.450 1683.780 1885.455 1683.920 ;
        RECT 1818.450 1683.720 1818.770 1683.780 ;
        RECT 1885.165 1683.735 1885.455 1683.780 ;
        RECT 1501.510 19.960 1501.830 20.020 ;
        RECT 1818.450 19.960 1818.770 20.020 ;
        RECT 1501.510 19.820 1818.770 19.960 ;
        RECT 1501.510 19.760 1501.830 19.820 ;
        RECT 1818.450 19.760 1818.770 19.820 ;
      LAYER via ;
        RECT 1920.140 1687.460 1920.400 1687.720 ;
        RECT 1818.480 1683.720 1818.740 1683.980 ;
        RECT 1501.540 19.760 1501.800 20.020 ;
        RECT 1818.480 19.760 1818.740 20.020 ;
      LAYER met2 ;
        RECT 1921.440 1700.410 1921.720 1704.000 ;
        RECT 1920.200 1700.270 1921.720 1700.410 ;
        RECT 1920.200 1687.750 1920.340 1700.270 ;
        RECT 1921.440 1700.000 1921.720 1700.270 ;
        RECT 1920.140 1687.430 1920.400 1687.750 ;
        RECT 1818.480 1683.690 1818.740 1684.010 ;
        RECT 1818.540 20.050 1818.680 1683.690 ;
        RECT 1501.540 19.730 1501.800 20.050 ;
        RECT 1818.480 19.730 1818.740 20.050 ;
        RECT 1501.600 2.400 1501.740 19.730 ;
        RECT 1501.390 -4.800 1501.950 2.400 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1914.590 1683.920 1914.910 1683.980 ;
        RECT 1930.690 1683.920 1931.010 1683.980 ;
        RECT 1914.590 1683.780 1931.010 1683.920 ;
        RECT 1914.590 1683.720 1914.910 1683.780 ;
        RECT 1930.690 1683.720 1931.010 1683.780 ;
        RECT 1518.990 18.260 1519.310 18.320 ;
        RECT 1914.590 18.260 1914.910 18.320 ;
        RECT 1518.990 18.120 1914.910 18.260 ;
        RECT 1518.990 18.060 1519.310 18.120 ;
        RECT 1914.590 18.060 1914.910 18.120 ;
      LAYER via ;
        RECT 1914.620 1683.720 1914.880 1683.980 ;
        RECT 1930.720 1683.720 1930.980 1683.980 ;
        RECT 1519.020 18.060 1519.280 18.320 ;
        RECT 1914.620 18.060 1914.880 18.320 ;
      LAYER met2 ;
        RECT 1930.640 1700.000 1930.920 1704.000 ;
        RECT 1930.780 1684.010 1930.920 1700.000 ;
        RECT 1914.620 1683.690 1914.880 1684.010 ;
        RECT 1930.720 1683.690 1930.980 1684.010 ;
        RECT 1914.680 18.350 1914.820 1683.690 ;
        RECT 1519.020 18.030 1519.280 18.350 ;
        RECT 1914.620 18.030 1914.880 18.350 ;
        RECT 1519.080 2.400 1519.220 18.030 ;
        RECT 1518.870 -4.800 1519.430 2.400 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1511.630 1678.140 1511.950 1678.200 ;
        RECT 1515.310 1678.140 1515.630 1678.200 ;
        RECT 1511.630 1678.000 1515.630 1678.140 ;
        RECT 1511.630 1677.940 1511.950 1678.000 ;
        RECT 1515.310 1677.940 1515.630 1678.000 ;
        RECT 717.210 54.980 717.530 55.040 ;
        RECT 1511.630 54.980 1511.950 55.040 ;
        RECT 717.210 54.840 1511.950 54.980 ;
        RECT 717.210 54.780 717.530 54.840 ;
        RECT 1511.630 54.780 1511.950 54.840 ;
      LAYER via ;
        RECT 1511.660 1677.940 1511.920 1678.200 ;
        RECT 1515.340 1677.940 1515.600 1678.200 ;
        RECT 717.240 54.780 717.500 55.040 ;
        RECT 1511.660 54.780 1511.920 55.040 ;
      LAYER met2 ;
        RECT 1517.100 1700.410 1517.380 1704.000 ;
        RECT 1515.400 1700.270 1517.380 1700.410 ;
        RECT 1515.400 1678.230 1515.540 1700.270 ;
        RECT 1517.100 1700.000 1517.380 1700.270 ;
        RECT 1511.660 1677.910 1511.920 1678.230 ;
        RECT 1515.340 1677.910 1515.600 1678.230 ;
        RECT 1511.720 55.070 1511.860 1677.910 ;
        RECT 717.240 54.750 717.500 55.070 ;
        RECT 1511.660 54.750 1511.920 55.070 ;
        RECT 717.300 16.730 717.440 54.750 ;
        RECT 716.380 16.590 717.440 16.730 ;
        RECT 716.380 2.400 716.520 16.590 ;
        RECT 716.170 -4.800 716.730 2.400 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1548.890 1689.700 1549.210 1689.760 ;
        RECT 1548.890 1689.560 1577.640 1689.700 ;
        RECT 1548.890 1689.500 1549.210 1689.560 ;
        RECT 1577.500 1689.360 1577.640 1689.560 ;
        RECT 1939.890 1689.360 1940.210 1689.420 ;
        RECT 1577.500 1689.220 1940.210 1689.360 ;
        RECT 1939.890 1689.160 1940.210 1689.220 ;
        RECT 1536.930 18.600 1537.250 18.660 ;
        RECT 1548.890 18.600 1549.210 18.660 ;
        RECT 1536.930 18.460 1549.210 18.600 ;
        RECT 1536.930 18.400 1537.250 18.460 ;
        RECT 1548.890 18.400 1549.210 18.460 ;
      LAYER via ;
        RECT 1548.920 1689.500 1549.180 1689.760 ;
        RECT 1939.920 1689.160 1940.180 1689.420 ;
        RECT 1536.960 18.400 1537.220 18.660 ;
        RECT 1548.920 18.400 1549.180 18.660 ;
      LAYER met2 ;
        RECT 1939.840 1700.000 1940.120 1704.000 ;
        RECT 1548.920 1689.470 1549.180 1689.790 ;
        RECT 1548.980 18.690 1549.120 1689.470 ;
        RECT 1939.980 1689.450 1940.120 1700.000 ;
        RECT 1939.920 1689.130 1940.180 1689.450 ;
        RECT 1536.960 18.370 1537.220 18.690 ;
        RECT 1548.920 18.370 1549.180 18.690 ;
        RECT 1537.020 2.400 1537.160 18.370 ;
        RECT 1536.810 -4.800 1537.370 2.400 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1928.390 1689.700 1928.710 1689.760 ;
        RECT 1948.630 1689.700 1948.950 1689.760 ;
        RECT 1928.390 1689.560 1948.950 1689.700 ;
        RECT 1928.390 1689.500 1928.710 1689.560 ;
        RECT 1948.630 1689.500 1948.950 1689.560 ;
        RECT 1554.870 14.180 1555.190 14.240 ;
        RECT 1928.390 14.180 1928.710 14.240 ;
        RECT 1554.870 14.040 1928.710 14.180 ;
        RECT 1554.870 13.980 1555.190 14.040 ;
        RECT 1928.390 13.980 1928.710 14.040 ;
      LAYER via ;
        RECT 1928.420 1689.500 1928.680 1689.760 ;
        RECT 1948.660 1689.500 1948.920 1689.760 ;
        RECT 1554.900 13.980 1555.160 14.240 ;
        RECT 1928.420 13.980 1928.680 14.240 ;
      LAYER met2 ;
        RECT 1948.580 1700.000 1948.860 1704.000 ;
        RECT 1948.720 1689.790 1948.860 1700.000 ;
        RECT 1928.420 1689.470 1928.680 1689.790 ;
        RECT 1948.660 1689.470 1948.920 1689.790 ;
        RECT 1928.480 14.270 1928.620 1689.470 ;
        RECT 1554.900 13.950 1555.160 14.270 ;
        RECT 1928.420 13.950 1928.680 14.270 ;
        RECT 1554.960 2.400 1555.100 13.950 ;
        RECT 1554.750 -4.800 1555.310 2.400 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1631.765 1685.805 1631.935 1689.715 ;
        RECT 1921.565 1687.845 1921.735 1689.715 ;
      LAYER mcon ;
        RECT 1631.765 1689.545 1631.935 1689.715 ;
        RECT 1921.565 1689.545 1921.735 1689.715 ;
      LAYER met1 ;
        RECT 1631.705 1689.700 1631.995 1689.745 ;
        RECT 1921.505 1689.700 1921.795 1689.745 ;
        RECT 1631.705 1689.560 1921.795 1689.700 ;
        RECT 1631.705 1689.515 1631.995 1689.560 ;
        RECT 1921.505 1689.515 1921.795 1689.560 ;
        RECT 1921.505 1688.000 1921.795 1688.045 ;
        RECT 1957.830 1688.000 1958.150 1688.060 ;
        RECT 1921.505 1687.860 1958.150 1688.000 ;
        RECT 1921.505 1687.815 1921.795 1687.860 ;
        RECT 1957.830 1687.800 1958.150 1687.860 ;
        RECT 1583.390 1685.960 1583.710 1686.020 ;
        RECT 1631.705 1685.960 1631.995 1686.005 ;
        RECT 1583.390 1685.820 1631.995 1685.960 ;
        RECT 1583.390 1685.760 1583.710 1685.820 ;
        RECT 1631.705 1685.775 1631.995 1685.820 ;
        RECT 1572.810 20.640 1573.130 20.700 ;
        RECT 1583.390 20.640 1583.710 20.700 ;
        RECT 1572.810 20.500 1583.710 20.640 ;
        RECT 1572.810 20.440 1573.130 20.500 ;
        RECT 1583.390 20.440 1583.710 20.500 ;
      LAYER via ;
        RECT 1957.860 1687.800 1958.120 1688.060 ;
        RECT 1583.420 1685.760 1583.680 1686.020 ;
        RECT 1572.840 20.440 1573.100 20.700 ;
        RECT 1583.420 20.440 1583.680 20.700 ;
      LAYER met2 ;
        RECT 1957.780 1700.000 1958.060 1704.000 ;
        RECT 1957.920 1688.090 1958.060 1700.000 ;
        RECT 1957.860 1687.770 1958.120 1688.090 ;
        RECT 1583.420 1685.730 1583.680 1686.050 ;
        RECT 1583.480 20.730 1583.620 1685.730 ;
        RECT 1572.840 20.410 1573.100 20.730 ;
        RECT 1583.420 20.410 1583.680 20.730 ;
        RECT 1572.900 2.400 1573.040 20.410 ;
        RECT 1572.690 -4.800 1573.250 2.400 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1949.550 1683.920 1949.870 1683.980 ;
        RECT 1967.030 1683.920 1967.350 1683.980 ;
        RECT 1949.550 1683.780 1967.350 1683.920 ;
        RECT 1949.550 1683.720 1949.870 1683.780 ;
        RECT 1967.030 1683.720 1967.350 1683.780 ;
        RECT 1590.290 18.940 1590.610 19.000 ;
        RECT 1949.090 18.940 1949.410 19.000 ;
        RECT 1590.290 18.800 1949.410 18.940 ;
        RECT 1590.290 18.740 1590.610 18.800 ;
        RECT 1949.090 18.740 1949.410 18.800 ;
      LAYER via ;
        RECT 1949.580 1683.720 1949.840 1683.980 ;
        RECT 1967.060 1683.720 1967.320 1683.980 ;
        RECT 1590.320 18.740 1590.580 19.000 ;
        RECT 1949.120 18.740 1949.380 19.000 ;
      LAYER met2 ;
        RECT 1966.980 1700.000 1967.260 1704.000 ;
        RECT 1967.120 1684.010 1967.260 1700.000 ;
        RECT 1949.580 1683.690 1949.840 1684.010 ;
        RECT 1967.060 1683.690 1967.320 1684.010 ;
        RECT 1949.640 1677.970 1949.780 1683.690 ;
        RECT 1949.180 1677.830 1949.780 1677.970 ;
        RECT 1949.180 19.030 1949.320 1677.830 ;
        RECT 1590.320 18.710 1590.580 19.030 ;
        RECT 1949.120 18.710 1949.380 19.030 ;
        RECT 1590.380 2.400 1590.520 18.710 ;
        RECT 1590.170 -4.800 1590.730 2.400 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1613.750 1690.040 1614.070 1690.100 ;
        RECT 1976.230 1690.040 1976.550 1690.100 ;
        RECT 1613.750 1689.900 1976.550 1690.040 ;
        RECT 1613.750 1689.840 1614.070 1689.900 ;
        RECT 1976.230 1689.840 1976.550 1689.900 ;
        RECT 1608.230 20.640 1608.550 20.700 ;
        RECT 1613.750 20.640 1614.070 20.700 ;
        RECT 1608.230 20.500 1614.070 20.640 ;
        RECT 1608.230 20.440 1608.550 20.500 ;
        RECT 1613.750 20.440 1614.070 20.500 ;
      LAYER via ;
        RECT 1613.780 1689.840 1614.040 1690.100 ;
        RECT 1976.260 1689.840 1976.520 1690.100 ;
        RECT 1608.260 20.440 1608.520 20.700 ;
        RECT 1613.780 20.440 1614.040 20.700 ;
      LAYER met2 ;
        RECT 1976.180 1700.000 1976.460 1704.000 ;
        RECT 1976.320 1690.130 1976.460 1700.000 ;
        RECT 1613.780 1689.810 1614.040 1690.130 ;
        RECT 1976.260 1689.810 1976.520 1690.130 ;
        RECT 1613.840 20.730 1613.980 1689.810 ;
        RECT 1608.260 20.410 1608.520 20.730 ;
        RECT 1613.780 20.410 1614.040 20.730 ;
        RECT 1608.320 2.400 1608.460 20.410 ;
        RECT 1608.110 -4.800 1608.670 2.400 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1955.990 1689.360 1956.310 1689.420 ;
        RECT 1985.430 1689.360 1985.750 1689.420 ;
        RECT 1955.990 1689.220 1985.750 1689.360 ;
        RECT 1955.990 1689.160 1956.310 1689.220 ;
        RECT 1985.430 1689.160 1985.750 1689.220 ;
        RECT 1626.170 19.620 1626.490 19.680 ;
        RECT 1955.990 19.620 1956.310 19.680 ;
        RECT 1626.170 19.480 1956.310 19.620 ;
        RECT 1626.170 19.420 1626.490 19.480 ;
        RECT 1955.990 19.420 1956.310 19.480 ;
      LAYER via ;
        RECT 1956.020 1689.160 1956.280 1689.420 ;
        RECT 1985.460 1689.160 1985.720 1689.420 ;
        RECT 1626.200 19.420 1626.460 19.680 ;
        RECT 1956.020 19.420 1956.280 19.680 ;
      LAYER met2 ;
        RECT 1985.380 1700.000 1985.660 1704.000 ;
        RECT 1985.520 1689.450 1985.660 1700.000 ;
        RECT 1956.020 1689.130 1956.280 1689.450 ;
        RECT 1985.460 1689.130 1985.720 1689.450 ;
        RECT 1956.080 19.710 1956.220 1689.130 ;
        RECT 1626.200 19.390 1626.460 19.710 ;
        RECT 1956.020 19.390 1956.280 19.710 ;
        RECT 1626.260 2.400 1626.400 19.390 ;
        RECT 1626.050 -4.800 1626.610 2.400 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1817.990 1684.260 1818.310 1684.320 ;
        RECT 1994.630 1684.260 1994.950 1684.320 ;
        RECT 1817.990 1684.120 1994.950 1684.260 ;
        RECT 1817.990 1684.060 1818.310 1684.120 ;
        RECT 1994.630 1684.060 1994.950 1684.120 ;
        RECT 1644.110 16.220 1644.430 16.280 ;
        RECT 1817.990 16.220 1818.310 16.280 ;
        RECT 1644.110 16.080 1818.310 16.220 ;
        RECT 1644.110 16.020 1644.430 16.080 ;
        RECT 1817.990 16.020 1818.310 16.080 ;
      LAYER via ;
        RECT 1818.020 1684.060 1818.280 1684.320 ;
        RECT 1994.660 1684.060 1994.920 1684.320 ;
        RECT 1644.140 16.020 1644.400 16.280 ;
        RECT 1818.020 16.020 1818.280 16.280 ;
      LAYER met2 ;
        RECT 1994.580 1700.000 1994.860 1704.000 ;
        RECT 1994.720 1684.350 1994.860 1700.000 ;
        RECT 1818.020 1684.030 1818.280 1684.350 ;
        RECT 1994.660 1684.030 1994.920 1684.350 ;
        RECT 1818.080 16.310 1818.220 1684.030 ;
        RECT 1644.140 15.990 1644.400 16.310 ;
        RECT 1818.020 15.990 1818.280 16.310 ;
        RECT 1644.200 2.400 1644.340 15.990 ;
        RECT 1643.990 -4.800 1644.550 2.400 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1977.150 1684.600 1977.470 1684.660 ;
        RECT 2003.830 1684.600 2004.150 1684.660 ;
        RECT 1977.150 1684.460 2004.150 1684.600 ;
        RECT 1977.150 1684.400 1977.470 1684.460 ;
        RECT 2003.830 1684.400 2004.150 1684.460 ;
        RECT 1662.050 19.280 1662.370 19.340 ;
        RECT 1662.050 19.140 1961.280 19.280 ;
        RECT 1662.050 19.080 1662.370 19.140 ;
        RECT 1961.140 18.940 1961.280 19.140 ;
        RECT 1976.690 18.940 1977.010 19.000 ;
        RECT 1961.140 18.800 1977.010 18.940 ;
        RECT 1976.690 18.740 1977.010 18.800 ;
      LAYER via ;
        RECT 1977.180 1684.400 1977.440 1684.660 ;
        RECT 2003.860 1684.400 2004.120 1684.660 ;
        RECT 1662.080 19.080 1662.340 19.340 ;
        RECT 1976.720 18.740 1976.980 19.000 ;
      LAYER met2 ;
        RECT 2003.780 1700.000 2004.060 1704.000 ;
        RECT 2003.920 1684.690 2004.060 1700.000 ;
        RECT 1977.180 1684.370 1977.440 1684.690 ;
        RECT 2003.860 1684.370 2004.120 1684.690 ;
        RECT 1977.240 1656.210 1977.380 1684.370 ;
        RECT 1976.780 1656.070 1977.380 1656.210 ;
        RECT 1662.080 19.050 1662.340 19.370 ;
        RECT 1662.140 2.400 1662.280 19.050 ;
        RECT 1976.780 19.030 1976.920 1656.070 ;
        RECT 1976.720 18.710 1976.980 19.030 ;
        RECT 1661.930 -4.800 1662.490 2.400 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1976.765 1684.445 1976.935 1690.055 ;
      LAYER mcon ;
        RECT 1976.765 1689.885 1976.935 1690.055 ;
      LAYER met1 ;
        RECT 1976.705 1690.040 1976.995 1690.085 ;
        RECT 2013.030 1690.040 2013.350 1690.100 ;
        RECT 1976.705 1689.900 2013.350 1690.040 ;
        RECT 1976.705 1689.855 1976.995 1689.900 ;
        RECT 2013.030 1689.840 2013.350 1689.900 ;
        RECT 1831.790 1684.600 1832.110 1684.660 ;
        RECT 1976.705 1684.600 1976.995 1684.645 ;
        RECT 1831.790 1684.460 1976.995 1684.600 ;
        RECT 1831.790 1684.400 1832.110 1684.460 ;
        RECT 1976.705 1684.415 1976.995 1684.460 ;
        RECT 1679.530 15.540 1679.850 15.600 ;
        RECT 1831.790 15.540 1832.110 15.600 ;
        RECT 1679.530 15.400 1832.110 15.540 ;
        RECT 1679.530 15.340 1679.850 15.400 ;
        RECT 1831.790 15.340 1832.110 15.400 ;
      LAYER via ;
        RECT 2013.060 1689.840 2013.320 1690.100 ;
        RECT 1831.820 1684.400 1832.080 1684.660 ;
        RECT 1679.560 15.340 1679.820 15.600 ;
        RECT 1831.820 15.340 1832.080 15.600 ;
      LAYER met2 ;
        RECT 2012.980 1700.000 2013.260 1704.000 ;
        RECT 2013.120 1690.130 2013.260 1700.000 ;
        RECT 2013.060 1689.810 2013.320 1690.130 ;
        RECT 1831.820 1684.370 1832.080 1684.690 ;
        RECT 1831.880 15.630 1832.020 1684.370 ;
        RECT 1679.560 15.310 1679.820 15.630 ;
        RECT 1831.820 15.310 1832.080 15.630 ;
        RECT 1679.620 2.400 1679.760 15.310 ;
        RECT 1679.410 -4.800 1679.970 2.400 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1964.805 19.465 1964.975 20.315 ;
      LAYER mcon ;
        RECT 1964.805 20.145 1964.975 20.315 ;
      LAYER met1 ;
        RECT 2022.230 1684.260 2022.550 1684.320 ;
        RECT 2004.380 1684.120 2022.550 1684.260 ;
        RECT 1983.590 1683.920 1983.910 1683.980 ;
        RECT 2004.380 1683.920 2004.520 1684.120 ;
        RECT 2022.230 1684.060 2022.550 1684.120 ;
        RECT 1983.590 1683.780 2004.520 1683.920 ;
        RECT 1983.590 1683.720 1983.910 1683.780 ;
        RECT 1697.470 20.300 1697.790 20.360 ;
        RECT 1964.745 20.300 1965.035 20.345 ;
        RECT 1697.470 20.160 1965.035 20.300 ;
        RECT 1697.470 20.100 1697.790 20.160 ;
        RECT 1964.745 20.115 1965.035 20.160 ;
        RECT 1964.745 19.620 1965.035 19.665 ;
        RECT 1983.590 19.620 1983.910 19.680 ;
        RECT 1964.745 19.480 1983.910 19.620 ;
        RECT 1964.745 19.435 1965.035 19.480 ;
        RECT 1983.590 19.420 1983.910 19.480 ;
      LAYER via ;
        RECT 1983.620 1683.720 1983.880 1683.980 ;
        RECT 2022.260 1684.060 2022.520 1684.320 ;
        RECT 1697.500 20.100 1697.760 20.360 ;
        RECT 1983.620 19.420 1983.880 19.680 ;
      LAYER met2 ;
        RECT 2022.180 1700.000 2022.460 1704.000 ;
        RECT 2022.320 1684.350 2022.460 1700.000 ;
        RECT 2022.260 1684.030 2022.520 1684.350 ;
        RECT 1983.620 1683.690 1983.880 1684.010 ;
        RECT 1697.500 20.070 1697.760 20.390 ;
        RECT 1697.560 2.400 1697.700 20.070 ;
        RECT 1983.680 19.710 1983.820 1683.690 ;
        RECT 1983.620 19.390 1983.880 19.710 ;
        RECT 1697.350 -4.800 1697.910 2.400 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 737.910 51.240 738.230 51.300 ;
        RECT 1524.970 51.240 1525.290 51.300 ;
        RECT 737.910 51.100 1525.290 51.240 ;
        RECT 737.910 51.040 738.230 51.100 ;
        RECT 1524.970 51.040 1525.290 51.100 ;
      LAYER via ;
        RECT 737.940 51.040 738.200 51.300 ;
        RECT 1525.000 51.040 1525.260 51.300 ;
      LAYER met2 ;
        RECT 1526.300 1700.410 1526.580 1704.000 ;
        RECT 1525.060 1700.270 1526.580 1700.410 ;
        RECT 1525.060 51.330 1525.200 1700.270 ;
        RECT 1526.300 1700.000 1526.580 1700.270 ;
        RECT 737.940 51.010 738.200 51.330 ;
        RECT 1525.000 51.010 1525.260 51.330 ;
        RECT 738.000 16.730 738.140 51.010 ;
        RECT 734.320 16.590 738.140 16.730 ;
        RECT 734.320 2.400 734.460 16.590 ;
        RECT 734.110 -4.800 734.670 2.400 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1864.525 15.725 1864.695 17.595 ;
      LAYER mcon ;
        RECT 1864.525 17.425 1864.695 17.595 ;
      LAYER met1 ;
        RECT 1880.090 1689.020 1880.410 1689.080 ;
        RECT 2031.430 1689.020 2031.750 1689.080 ;
        RECT 1880.090 1688.880 2031.750 1689.020 ;
        RECT 1880.090 1688.820 1880.410 1688.880 ;
        RECT 2031.430 1688.820 2031.750 1688.880 ;
        RECT 1864.465 17.580 1864.755 17.625 ;
        RECT 1880.090 17.580 1880.410 17.640 ;
        RECT 1864.465 17.440 1880.410 17.580 ;
        RECT 1864.465 17.395 1864.755 17.440 ;
        RECT 1880.090 17.380 1880.410 17.440 ;
        RECT 1715.410 15.880 1715.730 15.940 ;
        RECT 1864.465 15.880 1864.755 15.925 ;
        RECT 1715.410 15.740 1864.755 15.880 ;
        RECT 1715.410 15.680 1715.730 15.740 ;
        RECT 1864.465 15.695 1864.755 15.740 ;
      LAYER via ;
        RECT 1880.120 1688.820 1880.380 1689.080 ;
        RECT 2031.460 1688.820 2031.720 1689.080 ;
        RECT 1880.120 17.380 1880.380 17.640 ;
        RECT 1715.440 15.680 1715.700 15.940 ;
      LAYER met2 ;
        RECT 2031.380 1700.000 2031.660 1704.000 ;
        RECT 2031.520 1689.110 2031.660 1700.000 ;
        RECT 1880.120 1688.790 1880.380 1689.110 ;
        RECT 2031.460 1688.790 2031.720 1689.110 ;
        RECT 1880.180 17.670 1880.320 1688.790 ;
        RECT 1880.120 17.350 1880.380 17.670 ;
        RECT 1715.440 15.650 1715.700 15.970 ;
        RECT 1715.500 2.400 1715.640 15.650 ;
        RECT 1715.290 -4.800 1715.850 2.400 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1969.865 19.125 1970.035 20.655 ;
      LAYER mcon ;
        RECT 1969.865 20.485 1970.035 20.655 ;
      LAYER met1 ;
        RECT 2005.210 1683.920 2005.530 1683.980 ;
        RECT 2040.630 1683.920 2040.950 1683.980 ;
        RECT 2005.210 1683.780 2040.950 1683.920 ;
        RECT 2005.210 1683.720 2005.530 1683.780 ;
        RECT 2040.630 1683.720 2040.950 1683.780 ;
        RECT 1733.350 20.640 1733.670 20.700 ;
        RECT 1969.805 20.640 1970.095 20.685 ;
        RECT 1733.350 20.500 1970.095 20.640 ;
        RECT 1733.350 20.440 1733.670 20.500 ;
        RECT 1969.805 20.455 1970.095 20.500 ;
        RECT 1969.805 19.280 1970.095 19.325 ;
        RECT 2004.290 19.280 2004.610 19.340 ;
        RECT 1969.805 19.140 2004.610 19.280 ;
        RECT 1969.805 19.095 1970.095 19.140 ;
        RECT 2004.290 19.080 2004.610 19.140 ;
      LAYER via ;
        RECT 2005.240 1683.720 2005.500 1683.980 ;
        RECT 2040.660 1683.720 2040.920 1683.980 ;
        RECT 1733.380 20.440 1733.640 20.700 ;
        RECT 2004.320 19.080 2004.580 19.340 ;
      LAYER met2 ;
        RECT 2040.580 1700.000 2040.860 1704.000 ;
        RECT 2040.720 1684.010 2040.860 1700.000 ;
        RECT 2005.240 1683.690 2005.500 1684.010 ;
        RECT 2040.660 1683.690 2040.920 1684.010 ;
        RECT 2005.300 1656.210 2005.440 1683.690 ;
        RECT 2004.380 1656.070 2005.440 1656.210 ;
        RECT 1733.380 20.410 1733.640 20.730 ;
        RECT 1733.440 2.400 1733.580 20.410 ;
        RECT 2004.380 19.370 2004.520 1656.070 ;
        RECT 2004.320 19.050 2004.580 19.370 ;
        RECT 1733.230 -4.800 1733.790 2.400 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1873.190 1688.680 1873.510 1688.740 ;
        RECT 2049.830 1688.680 2050.150 1688.740 ;
        RECT 1873.190 1688.540 2050.150 1688.680 ;
        RECT 1873.190 1688.480 1873.510 1688.540 ;
        RECT 2049.830 1688.480 2050.150 1688.540 ;
        RECT 1751.290 15.200 1751.610 15.260 ;
        RECT 1872.730 15.200 1873.050 15.260 ;
        RECT 1751.290 15.060 1873.050 15.200 ;
        RECT 1751.290 15.000 1751.610 15.060 ;
        RECT 1872.730 15.000 1873.050 15.060 ;
      LAYER via ;
        RECT 1873.220 1688.480 1873.480 1688.740 ;
        RECT 2049.860 1688.480 2050.120 1688.740 ;
        RECT 1751.320 15.000 1751.580 15.260 ;
        RECT 1872.760 15.000 1873.020 15.260 ;
      LAYER met2 ;
        RECT 2049.780 1700.000 2050.060 1704.000 ;
        RECT 2049.920 1688.770 2050.060 1700.000 ;
        RECT 1873.220 1688.450 1873.480 1688.770 ;
        RECT 2049.860 1688.450 2050.120 1688.770 ;
        RECT 1873.280 15.370 1873.420 1688.450 ;
        RECT 1872.820 15.290 1873.420 15.370 ;
        RECT 1751.320 14.970 1751.580 15.290 ;
        RECT 1872.760 15.230 1873.420 15.290 ;
        RECT 1872.760 14.970 1873.020 15.230 ;
        RECT 1751.380 2.400 1751.520 14.970 ;
        RECT 1751.170 -4.800 1751.730 2.400 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1969.405 16.745 1969.575 20.315 ;
      LAYER mcon ;
        RECT 1969.405 20.145 1969.575 20.315 ;
      LAYER met1 ;
        RECT 2024.990 1689.360 2025.310 1689.420 ;
        RECT 2059.030 1689.360 2059.350 1689.420 ;
        RECT 2024.990 1689.220 2059.350 1689.360 ;
        RECT 2024.990 1689.160 2025.310 1689.220 ;
        RECT 2059.030 1689.160 2059.350 1689.220 ;
        RECT 2024.990 20.980 2025.310 21.040 ;
        RECT 2017.260 20.840 2025.310 20.980 ;
        RECT 1969.345 20.300 1969.635 20.345 ;
        RECT 2017.260 20.300 2017.400 20.840 ;
        RECT 2024.990 20.780 2025.310 20.840 ;
        RECT 1969.345 20.160 2017.400 20.300 ;
        RECT 1969.345 20.115 1969.635 20.160 ;
        RECT 1768.770 16.900 1769.090 16.960 ;
        RECT 1969.345 16.900 1969.635 16.945 ;
        RECT 1768.770 16.760 1969.635 16.900 ;
        RECT 1768.770 16.700 1769.090 16.760 ;
        RECT 1969.345 16.715 1969.635 16.760 ;
      LAYER via ;
        RECT 2025.020 1689.160 2025.280 1689.420 ;
        RECT 2059.060 1689.160 2059.320 1689.420 ;
        RECT 2025.020 20.780 2025.280 21.040 ;
        RECT 1768.800 16.700 1769.060 16.960 ;
      LAYER met2 ;
        RECT 2058.980 1700.000 2059.260 1704.000 ;
        RECT 2059.120 1689.450 2059.260 1700.000 ;
        RECT 2025.020 1689.130 2025.280 1689.450 ;
        RECT 2059.060 1689.130 2059.320 1689.450 ;
        RECT 2025.080 21.070 2025.220 1689.130 ;
        RECT 2025.020 20.750 2025.280 21.070 ;
        RECT 1768.800 16.670 1769.060 16.990 ;
        RECT 1768.860 2.400 1769.000 16.670 ;
        RECT 1768.650 -4.800 1769.210 2.400 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1786.710 1685.620 1787.030 1685.680 ;
        RECT 2068.230 1685.620 2068.550 1685.680 ;
        RECT 1786.710 1685.480 2068.550 1685.620 ;
        RECT 1786.710 1685.420 1787.030 1685.480 ;
        RECT 2068.230 1685.420 2068.550 1685.480 ;
      LAYER via ;
        RECT 1786.740 1685.420 1787.000 1685.680 ;
        RECT 2068.260 1685.420 2068.520 1685.680 ;
      LAYER met2 ;
        RECT 2068.180 1700.000 2068.460 1704.000 ;
        RECT 2068.320 1685.710 2068.460 1700.000 ;
        RECT 1786.740 1685.390 1787.000 1685.710 ;
        RECT 2068.260 1685.390 2068.520 1685.710 ;
        RECT 1786.800 2.400 1786.940 1685.390 ;
        RECT 1786.590 -4.800 1787.150 2.400 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2038.865 572.645 2039.035 620.755 ;
        RECT 2038.865 434.945 2039.035 524.195 ;
        RECT 2038.865 379.525 2039.035 427.635 ;
        RECT 2038.865 282.965 2039.035 331.075 ;
        RECT 2038.865 186.405 2039.035 234.515 ;
        RECT 2038.865 48.365 2039.035 137.955 ;
        RECT 2031.505 16.745 2031.675 21.335 ;
        RECT 2019.545 16.235 2019.715 16.575 ;
        RECT 2018.625 16.065 2019.715 16.235 ;
      LAYER mcon ;
        RECT 2038.865 620.585 2039.035 620.755 ;
        RECT 2038.865 524.025 2039.035 524.195 ;
        RECT 2038.865 427.465 2039.035 427.635 ;
        RECT 2038.865 330.905 2039.035 331.075 ;
        RECT 2038.865 234.345 2039.035 234.515 ;
        RECT 2038.865 137.785 2039.035 137.955 ;
        RECT 2031.505 21.165 2031.675 21.335 ;
        RECT 2019.545 16.405 2019.715 16.575 ;
      LAYER met1 ;
        RECT 2038.790 1689.700 2039.110 1689.760 ;
        RECT 2077.430 1689.700 2077.750 1689.760 ;
        RECT 2038.790 1689.560 2077.750 1689.700 ;
        RECT 2038.790 1689.500 2039.110 1689.560 ;
        RECT 2077.430 1689.500 2077.750 1689.560 ;
        RECT 2038.330 1255.860 2038.650 1255.920 ;
        RECT 2038.790 1255.860 2039.110 1255.920 ;
        RECT 2038.330 1255.720 2039.110 1255.860 ;
        RECT 2038.330 1255.660 2038.650 1255.720 ;
        RECT 2038.790 1255.660 2039.110 1255.720 ;
        RECT 2037.410 1200.780 2037.730 1200.840 ;
        RECT 2038.790 1200.780 2039.110 1200.840 ;
        RECT 2037.410 1200.640 2039.110 1200.780 ;
        RECT 2037.410 1200.580 2037.730 1200.640 ;
        RECT 2038.790 1200.580 2039.110 1200.640 ;
        RECT 2038.790 620.740 2039.110 620.800 ;
        RECT 2038.595 620.600 2039.110 620.740 ;
        RECT 2038.790 620.540 2039.110 620.600 ;
        RECT 2038.790 572.800 2039.110 572.860 ;
        RECT 2038.595 572.660 2039.110 572.800 ;
        RECT 2038.790 572.600 2039.110 572.660 ;
        RECT 2038.790 524.180 2039.110 524.240 ;
        RECT 2038.595 524.040 2039.110 524.180 ;
        RECT 2038.790 523.980 2039.110 524.040 ;
        RECT 2038.805 435.100 2039.095 435.145 ;
        RECT 2039.250 435.100 2039.570 435.160 ;
        RECT 2038.805 434.960 2039.570 435.100 ;
        RECT 2038.805 434.915 2039.095 434.960 ;
        RECT 2039.250 434.900 2039.570 434.960 ;
        RECT 2038.790 427.620 2039.110 427.680 ;
        RECT 2038.595 427.480 2039.110 427.620 ;
        RECT 2038.790 427.420 2039.110 427.480 ;
        RECT 2038.790 379.680 2039.110 379.740 ;
        RECT 2038.595 379.540 2039.110 379.680 ;
        RECT 2038.790 379.480 2039.110 379.540 ;
        RECT 2038.790 331.060 2039.110 331.120 ;
        RECT 2038.595 330.920 2039.110 331.060 ;
        RECT 2038.790 330.860 2039.110 330.920 ;
        RECT 2038.790 283.120 2039.110 283.180 ;
        RECT 2038.595 282.980 2039.110 283.120 ;
        RECT 2038.790 282.920 2039.110 282.980 ;
        RECT 2038.790 234.500 2039.110 234.560 ;
        RECT 2038.595 234.360 2039.110 234.500 ;
        RECT 2038.790 234.300 2039.110 234.360 ;
        RECT 2038.790 186.560 2039.110 186.620 ;
        RECT 2038.595 186.420 2039.110 186.560 ;
        RECT 2038.790 186.360 2039.110 186.420 ;
        RECT 2038.790 137.940 2039.110 138.000 ;
        RECT 2038.595 137.800 2039.110 137.940 ;
        RECT 2038.790 137.740 2039.110 137.800 ;
        RECT 2038.805 48.520 2039.095 48.565 ;
        RECT 2039.250 48.520 2039.570 48.580 ;
        RECT 2038.805 48.380 2039.570 48.520 ;
        RECT 2038.805 48.335 2039.095 48.380 ;
        RECT 2039.250 48.320 2039.570 48.380 ;
        RECT 2031.445 21.320 2031.735 21.365 ;
        RECT 2039.250 21.320 2039.570 21.380 ;
        RECT 2031.445 21.180 2039.570 21.320 ;
        RECT 2031.445 21.135 2031.735 21.180 ;
        RECT 2039.250 21.120 2039.570 21.180 ;
        RECT 2031.445 16.900 2031.735 16.945 ;
        RECT 2020.020 16.760 2031.735 16.900 ;
        RECT 1804.650 16.560 1804.970 16.620 ;
        RECT 2019.485 16.560 2019.775 16.605 ;
        RECT 2020.020 16.560 2020.160 16.760 ;
        RECT 2031.445 16.715 2031.735 16.760 ;
        RECT 1804.650 16.420 2018.780 16.560 ;
        RECT 1804.650 16.360 1804.970 16.420 ;
        RECT 2018.640 16.265 2018.780 16.420 ;
        RECT 2019.485 16.420 2020.160 16.560 ;
        RECT 2019.485 16.375 2019.775 16.420 ;
        RECT 2018.565 16.035 2018.855 16.265 ;
      LAYER via ;
        RECT 2038.820 1689.500 2039.080 1689.760 ;
        RECT 2077.460 1689.500 2077.720 1689.760 ;
        RECT 2038.360 1255.660 2038.620 1255.920 ;
        RECT 2038.820 1255.660 2039.080 1255.920 ;
        RECT 2037.440 1200.580 2037.700 1200.840 ;
        RECT 2038.820 1200.580 2039.080 1200.840 ;
        RECT 2038.820 620.540 2039.080 620.800 ;
        RECT 2038.820 572.600 2039.080 572.860 ;
        RECT 2038.820 523.980 2039.080 524.240 ;
        RECT 2039.280 434.900 2039.540 435.160 ;
        RECT 2038.820 427.420 2039.080 427.680 ;
        RECT 2038.820 379.480 2039.080 379.740 ;
        RECT 2038.820 330.860 2039.080 331.120 ;
        RECT 2038.820 282.920 2039.080 283.180 ;
        RECT 2038.820 234.300 2039.080 234.560 ;
        RECT 2038.820 186.360 2039.080 186.620 ;
        RECT 2038.820 137.740 2039.080 138.000 ;
        RECT 2039.280 48.320 2039.540 48.580 ;
        RECT 2039.280 21.120 2039.540 21.380 ;
        RECT 1804.680 16.360 1804.940 16.620 ;
      LAYER met2 ;
        RECT 2077.380 1700.000 2077.660 1704.000 ;
        RECT 2077.520 1689.790 2077.660 1700.000 ;
        RECT 2038.820 1689.470 2039.080 1689.790 ;
        RECT 2077.460 1689.470 2077.720 1689.790 ;
        RECT 2038.880 1255.950 2039.020 1689.470 ;
        RECT 2038.360 1255.630 2038.620 1255.950 ;
        RECT 2038.820 1255.630 2039.080 1255.950 ;
        RECT 2038.420 1249.005 2038.560 1255.630 ;
        RECT 2037.430 1248.635 2037.710 1249.005 ;
        RECT 2038.350 1248.635 2038.630 1249.005 ;
        RECT 2037.500 1200.870 2037.640 1248.635 ;
        RECT 2037.440 1200.550 2037.700 1200.870 ;
        RECT 2038.820 1200.550 2039.080 1200.870 ;
        RECT 2038.880 620.830 2039.020 1200.550 ;
        RECT 2038.820 620.510 2039.080 620.830 ;
        RECT 2038.820 572.570 2039.080 572.890 ;
        RECT 2038.880 524.270 2039.020 572.570 ;
        RECT 2038.820 523.950 2039.080 524.270 ;
        RECT 2039.280 434.930 2039.540 435.190 ;
        RECT 2038.880 434.870 2039.540 434.930 ;
        RECT 2038.880 434.790 2039.480 434.870 ;
        RECT 2038.880 427.710 2039.020 434.790 ;
        RECT 2038.820 427.390 2039.080 427.710 ;
        RECT 2038.820 379.450 2039.080 379.770 ;
        RECT 2038.880 331.150 2039.020 379.450 ;
        RECT 2038.820 330.830 2039.080 331.150 ;
        RECT 2038.820 282.890 2039.080 283.210 ;
        RECT 2038.880 234.590 2039.020 282.890 ;
        RECT 2038.820 234.270 2039.080 234.590 ;
        RECT 2038.820 186.330 2039.080 186.650 ;
        RECT 2038.880 138.030 2039.020 186.330 ;
        RECT 2038.820 137.710 2039.080 138.030 ;
        RECT 2039.280 48.290 2039.540 48.610 ;
        RECT 2039.340 21.410 2039.480 48.290 ;
        RECT 2039.280 21.090 2039.540 21.410 ;
        RECT 1804.680 16.330 1804.940 16.650 ;
        RECT 1804.740 2.400 1804.880 16.330 ;
        RECT 1804.530 -4.800 1805.090 2.400 ;
      LAYER via2 ;
        RECT 2037.430 1248.680 2037.710 1248.960 ;
        RECT 2038.350 1248.680 2038.630 1248.960 ;
      LAYER met3 ;
        RECT 2037.405 1248.970 2037.735 1248.985 ;
        RECT 2038.325 1248.970 2038.655 1248.985 ;
        RECT 2037.405 1248.670 2038.655 1248.970 ;
        RECT 2037.405 1248.655 2037.735 1248.670 ;
        RECT 2038.325 1248.655 2038.655 1248.670 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1832.250 1684.940 1832.570 1685.000 ;
        RECT 2086.630 1684.940 2086.950 1685.000 ;
        RECT 1832.250 1684.800 2086.950 1684.940 ;
        RECT 1832.250 1684.740 1832.570 1684.800 ;
        RECT 2086.630 1684.740 2086.950 1684.800 ;
        RECT 1822.590 19.960 1822.910 20.020 ;
        RECT 1832.250 19.960 1832.570 20.020 ;
        RECT 1822.590 19.820 1832.570 19.960 ;
        RECT 1822.590 19.760 1822.910 19.820 ;
        RECT 1832.250 19.760 1832.570 19.820 ;
      LAYER via ;
        RECT 1832.280 1684.740 1832.540 1685.000 ;
        RECT 2086.660 1684.740 2086.920 1685.000 ;
        RECT 1822.620 19.760 1822.880 20.020 ;
        RECT 1832.280 19.760 1832.540 20.020 ;
      LAYER met2 ;
        RECT 2086.580 1700.000 2086.860 1704.000 ;
        RECT 2086.720 1685.030 2086.860 1700.000 ;
        RECT 1832.280 1684.710 1832.540 1685.030 ;
        RECT 2086.660 1684.710 2086.920 1685.030 ;
        RECT 1832.340 20.050 1832.480 1684.710 ;
        RECT 1822.620 19.730 1822.880 20.050 ;
        RECT 1832.280 19.730 1832.540 20.050 ;
        RECT 1822.680 2.400 1822.820 19.730 ;
        RECT 1822.470 -4.800 1823.030 2.400 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2041.625 20.145 2042.255 20.315 ;
        RECT 1873.265 15.385 1873.435 19.975 ;
        RECT 2042.085 18.105 2042.255 20.145 ;
        RECT 2042.545 18.105 2043.175 18.275 ;
        RECT 2043.005 16.065 2043.175 18.105 ;
      LAYER mcon ;
        RECT 1873.265 19.805 1873.435 19.975 ;
      LAYER met1 ;
        RECT 2060.410 1690.380 2060.730 1690.440 ;
        RECT 2095.830 1690.380 2096.150 1690.440 ;
        RECT 2060.410 1690.240 2096.150 1690.380 ;
        RECT 2060.410 1690.180 2060.730 1690.240 ;
        RECT 2095.830 1690.180 2096.150 1690.240 ;
        RECT 2041.565 20.300 2041.855 20.345 ;
        RECT 2017.720 20.160 2041.855 20.300 ;
        RECT 1873.205 19.960 1873.495 20.005 ;
        RECT 2017.720 19.960 2017.860 20.160 ;
        RECT 2041.565 20.115 2041.855 20.160 ;
        RECT 1873.205 19.820 2017.860 19.960 ;
        RECT 1873.205 19.775 1873.495 19.820 ;
        RECT 2042.025 18.260 2042.315 18.305 ;
        RECT 2042.485 18.260 2042.775 18.305 ;
        RECT 2042.025 18.120 2042.775 18.260 ;
        RECT 2042.025 18.075 2042.315 18.120 ;
        RECT 2042.485 18.075 2042.775 18.120 ;
        RECT 2042.945 16.220 2043.235 16.265 ;
        RECT 2059.490 16.220 2059.810 16.280 ;
        RECT 2042.945 16.080 2059.810 16.220 ;
        RECT 2042.945 16.035 2043.235 16.080 ;
        RECT 2059.490 16.020 2059.810 16.080 ;
        RECT 1840.070 15.540 1840.390 15.600 ;
        RECT 1873.205 15.540 1873.495 15.585 ;
        RECT 1840.070 15.400 1873.495 15.540 ;
        RECT 1840.070 15.340 1840.390 15.400 ;
        RECT 1873.205 15.355 1873.495 15.400 ;
      LAYER via ;
        RECT 2060.440 1690.180 2060.700 1690.440 ;
        RECT 2095.860 1690.180 2096.120 1690.440 ;
        RECT 2059.520 16.020 2059.780 16.280 ;
        RECT 1840.100 15.340 1840.360 15.600 ;
      LAYER met2 ;
        RECT 2095.780 1700.000 2096.060 1704.000 ;
        RECT 2095.920 1690.470 2096.060 1700.000 ;
        RECT 2060.440 1690.150 2060.700 1690.470 ;
        RECT 2095.860 1690.150 2096.120 1690.470 ;
        RECT 2060.500 1656.210 2060.640 1690.150 ;
        RECT 2059.580 1656.070 2060.640 1656.210 ;
        RECT 2059.580 16.310 2059.720 1656.070 ;
        RECT 2059.520 15.990 2059.780 16.310 ;
        RECT 1840.100 15.310 1840.360 15.630 ;
        RECT 1840.160 2.400 1840.300 15.310 ;
        RECT 1839.950 -4.800 1840.510 2.400 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1862.610 1686.980 1862.930 1687.040 ;
        RECT 2105.030 1686.980 2105.350 1687.040 ;
        RECT 1862.610 1686.840 2105.350 1686.980 ;
        RECT 1862.610 1686.780 1862.930 1686.840 ;
        RECT 2105.030 1686.780 2105.350 1686.840 ;
        RECT 1858.010 14.860 1858.330 14.920 ;
        RECT 1862.610 14.860 1862.930 14.920 ;
        RECT 1858.010 14.720 1862.930 14.860 ;
        RECT 1858.010 14.660 1858.330 14.720 ;
        RECT 1862.610 14.660 1862.930 14.720 ;
      LAYER via ;
        RECT 1862.640 1686.780 1862.900 1687.040 ;
        RECT 2105.060 1686.780 2105.320 1687.040 ;
        RECT 1858.040 14.660 1858.300 14.920 ;
        RECT 1862.640 14.660 1862.900 14.920 ;
      LAYER met2 ;
        RECT 2104.980 1700.000 2105.260 1704.000 ;
        RECT 2105.120 1687.070 2105.260 1700.000 ;
        RECT 1862.640 1686.750 1862.900 1687.070 ;
        RECT 2105.060 1686.750 2105.320 1687.070 ;
        RECT 1862.700 14.950 1862.840 1686.750 ;
        RECT 1858.040 14.630 1858.300 14.950 ;
        RECT 1862.640 14.630 1862.900 14.950 ;
        RECT 1858.100 2.400 1858.240 14.630 ;
        RECT 1857.890 -4.800 1858.450 2.400 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2019.085 16.575 2019.255 17.255 ;
        RECT 2017.705 16.405 2019.255 16.575 ;
        RECT 2017.705 15.385 2017.875 16.405 ;
      LAYER mcon ;
        RECT 2019.085 17.085 2019.255 17.255 ;
      LAYER met1 ;
        RECT 2073.290 1685.620 2073.610 1685.680 ;
        RECT 2114.230 1685.620 2114.550 1685.680 ;
        RECT 2073.290 1685.480 2114.550 1685.620 ;
        RECT 2073.290 1685.420 2073.610 1685.480 ;
        RECT 2114.230 1685.420 2114.550 1685.480 ;
        RECT 2060.040 20.840 2063.400 20.980 ;
        RECT 2060.040 20.640 2060.180 20.840 ;
        RECT 2054.060 20.500 2060.180 20.640 ;
        RECT 2063.260 20.640 2063.400 20.840 ;
        RECT 2073.290 20.640 2073.610 20.700 ;
        RECT 2063.260 20.500 2073.610 20.640 ;
        RECT 2042.010 20.300 2042.330 20.360 ;
        RECT 2054.060 20.300 2054.200 20.500 ;
        RECT 2073.290 20.440 2073.610 20.500 ;
        RECT 2042.010 20.160 2054.200 20.300 ;
        RECT 2042.010 20.100 2042.330 20.160 ;
        RECT 2019.025 17.240 2019.315 17.285 ;
        RECT 2042.010 17.240 2042.330 17.300 ;
        RECT 2019.025 17.100 2042.330 17.240 ;
        RECT 2019.025 17.055 2019.315 17.100 ;
        RECT 2042.010 17.040 2042.330 17.100 ;
        RECT 1875.950 15.540 1876.270 15.600 ;
        RECT 2017.645 15.540 2017.935 15.585 ;
        RECT 1875.950 15.400 2017.935 15.540 ;
        RECT 1875.950 15.340 1876.270 15.400 ;
        RECT 2017.645 15.355 2017.935 15.400 ;
      LAYER via ;
        RECT 2073.320 1685.420 2073.580 1685.680 ;
        RECT 2114.260 1685.420 2114.520 1685.680 ;
        RECT 2042.040 20.100 2042.300 20.360 ;
        RECT 2073.320 20.440 2073.580 20.700 ;
        RECT 2042.040 17.040 2042.300 17.300 ;
        RECT 1875.980 15.340 1876.240 15.600 ;
      LAYER met2 ;
        RECT 2114.180 1700.000 2114.460 1704.000 ;
        RECT 2114.320 1685.710 2114.460 1700.000 ;
        RECT 2073.320 1685.390 2073.580 1685.710 ;
        RECT 2114.260 1685.390 2114.520 1685.710 ;
        RECT 2073.380 20.730 2073.520 1685.390 ;
        RECT 2073.320 20.410 2073.580 20.730 ;
        RECT 2042.040 20.070 2042.300 20.390 ;
        RECT 2042.100 17.330 2042.240 20.070 ;
        RECT 2042.040 17.010 2042.300 17.330 ;
        RECT 1875.980 15.310 1876.240 15.630 ;
        RECT 1876.040 2.400 1876.180 15.310 ;
        RECT 1875.830 -4.800 1876.390 2.400 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1531.870 1659.780 1532.190 1659.840 ;
        RECT 1533.710 1659.780 1534.030 1659.840 ;
        RECT 1531.870 1659.640 1534.030 1659.780 ;
        RECT 1531.870 1659.580 1532.190 1659.640 ;
        RECT 1533.710 1659.580 1534.030 1659.640 ;
        RECT 758.150 50.900 758.470 50.960 ;
        RECT 1531.870 50.900 1532.190 50.960 ;
        RECT 758.150 50.760 1532.190 50.900 ;
        RECT 758.150 50.700 758.470 50.760 ;
        RECT 1531.870 50.700 1532.190 50.760 ;
        RECT 752.170 20.980 752.490 21.040 ;
        RECT 758.150 20.980 758.470 21.040 ;
        RECT 752.170 20.840 758.470 20.980 ;
        RECT 752.170 20.780 752.490 20.840 ;
        RECT 758.150 20.780 758.470 20.840 ;
      LAYER via ;
        RECT 1531.900 1659.580 1532.160 1659.840 ;
        RECT 1533.740 1659.580 1534.000 1659.840 ;
        RECT 758.180 50.700 758.440 50.960 ;
        RECT 1531.900 50.700 1532.160 50.960 ;
        RECT 752.200 20.780 752.460 21.040 ;
        RECT 758.180 20.780 758.440 21.040 ;
      LAYER met2 ;
        RECT 1535.500 1700.410 1535.780 1704.000 ;
        RECT 1533.800 1700.270 1535.780 1700.410 ;
        RECT 1533.800 1659.870 1533.940 1700.270 ;
        RECT 1535.500 1700.000 1535.780 1700.270 ;
        RECT 1531.900 1659.550 1532.160 1659.870 ;
        RECT 1533.740 1659.550 1534.000 1659.870 ;
        RECT 1531.960 50.990 1532.100 1659.550 ;
        RECT 758.180 50.670 758.440 50.990 ;
        RECT 1531.900 50.670 1532.160 50.990 ;
        RECT 758.240 21.070 758.380 50.670 ;
        RECT 752.200 20.750 752.460 21.070 ;
        RECT 758.180 20.750 758.440 21.070 ;
        RECT 752.260 2.400 752.400 20.750 ;
        RECT 752.050 -4.800 752.610 2.400 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2080.190 1683.920 2080.510 1683.980 ;
        RECT 2121.130 1683.920 2121.450 1683.980 ;
        RECT 2080.190 1683.780 2121.450 1683.920 ;
        RECT 2080.190 1683.720 2080.510 1683.780 ;
        RECT 2121.130 1683.720 2121.450 1683.780 ;
        RECT 1893.890 15.200 1894.210 15.260 ;
        RECT 2042.930 15.200 2043.250 15.260 ;
        RECT 1893.890 15.060 2043.250 15.200 ;
        RECT 1893.890 15.000 1894.210 15.060 ;
        RECT 2042.930 15.000 2043.250 15.060 ;
        RECT 2042.930 14.520 2043.250 14.580 ;
        RECT 2080.190 14.520 2080.510 14.580 ;
        RECT 2042.930 14.380 2080.510 14.520 ;
        RECT 2042.930 14.320 2043.250 14.380 ;
        RECT 2080.190 14.320 2080.510 14.380 ;
      LAYER via ;
        RECT 2080.220 1683.720 2080.480 1683.980 ;
        RECT 2121.160 1683.720 2121.420 1683.980 ;
        RECT 1893.920 15.000 1894.180 15.260 ;
        RECT 2042.960 15.000 2043.220 15.260 ;
        RECT 2042.960 14.320 2043.220 14.580 ;
        RECT 2080.220 14.320 2080.480 14.580 ;
      LAYER met2 ;
        RECT 2123.380 1700.410 2123.660 1704.000 ;
        RECT 2121.220 1700.270 2123.660 1700.410 ;
        RECT 2121.220 1684.010 2121.360 1700.270 ;
        RECT 2123.380 1700.000 2123.660 1700.270 ;
        RECT 2080.220 1683.690 2080.480 1684.010 ;
        RECT 2121.160 1683.690 2121.420 1684.010 ;
        RECT 1893.920 14.970 1894.180 15.290 ;
        RECT 2042.960 14.970 2043.220 15.290 ;
        RECT 1893.980 2.400 1894.120 14.970 ;
        RECT 2043.020 14.610 2043.160 14.970 ;
        RECT 2080.280 14.610 2080.420 1683.690 ;
        RECT 2042.960 14.290 2043.220 14.610 ;
        RECT 2080.220 14.290 2080.480 14.610 ;
        RECT 1893.770 -4.800 1894.330 2.400 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2118.905 17.425 2119.075 18.275 ;
      LAYER mcon ;
        RECT 2118.905 18.105 2119.075 18.275 ;
      LAYER met1 ;
        RECT 2118.845 18.260 2119.135 18.305 ;
        RECT 2133.090 18.260 2133.410 18.320 ;
        RECT 2118.845 18.120 2133.410 18.260 ;
        RECT 2118.845 18.075 2119.135 18.120 ;
        RECT 2133.090 18.060 2133.410 18.120 ;
        RECT 1911.830 17.580 1912.150 17.640 ;
        RECT 2118.845 17.580 2119.135 17.625 ;
        RECT 1911.830 17.440 2119.135 17.580 ;
        RECT 1911.830 17.380 1912.150 17.440 ;
        RECT 2118.845 17.395 2119.135 17.440 ;
      LAYER via ;
        RECT 2133.120 18.060 2133.380 18.320 ;
        RECT 1911.860 17.380 1912.120 17.640 ;
      LAYER met2 ;
        RECT 2132.580 1700.410 2132.860 1704.000 ;
        RECT 2132.580 1700.270 2133.320 1700.410 ;
        RECT 2132.580 1700.000 2132.860 1700.270 ;
        RECT 2133.180 18.350 2133.320 1700.270 ;
        RECT 2133.120 18.030 2133.380 18.350 ;
        RECT 1911.860 17.350 1912.120 17.670 ;
        RECT 1911.920 2.400 1912.060 17.350 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2018.165 18.445 2018.335 19.975 ;
      LAYER mcon ;
        RECT 2018.165 19.805 2018.335 19.975 ;
      LAYER met1 ;
        RECT 2141.830 1686.640 2142.150 1686.700 ;
        RECT 2056.360 1686.500 2142.150 1686.640 ;
        RECT 2045.690 1686.300 2046.010 1686.360 ;
        RECT 2056.360 1686.300 2056.500 1686.500 ;
        RECT 2141.830 1686.440 2142.150 1686.500 ;
        RECT 2045.690 1686.160 2056.500 1686.300 ;
        RECT 2045.690 1686.100 2046.010 1686.160 ;
        RECT 2018.105 19.960 2018.395 20.005 ;
        RECT 2045.690 19.960 2046.010 20.020 ;
        RECT 2018.105 19.820 2046.010 19.960 ;
        RECT 2018.105 19.775 2018.395 19.820 ;
        RECT 2045.690 19.760 2046.010 19.820 ;
        RECT 1929.310 18.600 1929.630 18.660 ;
        RECT 2018.105 18.600 2018.395 18.645 ;
        RECT 1929.310 18.460 2018.395 18.600 ;
        RECT 1929.310 18.400 1929.630 18.460 ;
        RECT 2018.105 18.415 2018.395 18.460 ;
      LAYER via ;
        RECT 2045.720 1686.100 2045.980 1686.360 ;
        RECT 2141.860 1686.440 2142.120 1686.700 ;
        RECT 2045.720 19.760 2045.980 20.020 ;
        RECT 1929.340 18.400 1929.600 18.660 ;
      LAYER met2 ;
        RECT 2141.780 1700.000 2142.060 1704.000 ;
        RECT 2141.920 1686.730 2142.060 1700.000 ;
        RECT 2141.860 1686.410 2142.120 1686.730 ;
        RECT 2045.720 1686.070 2045.980 1686.390 ;
        RECT 2045.780 20.050 2045.920 1686.070 ;
        RECT 2045.720 19.730 2045.980 20.050 ;
        RECT 1929.340 18.370 1929.600 18.690 ;
        RECT 1929.400 2.400 1929.540 18.370 ;
        RECT 1929.190 -4.800 1929.750 2.400 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2090.845 14.365 2091.015 17.935 ;
        RECT 2133.625 14.365 2133.795 18.275 ;
      LAYER mcon ;
        RECT 2133.625 18.105 2133.795 18.275 ;
        RECT 2090.845 17.765 2091.015 17.935 ;
      LAYER met1 ;
        RECT 2133.565 18.260 2133.855 18.305 ;
        RECT 2146.430 18.260 2146.750 18.320 ;
        RECT 2133.565 18.120 2146.750 18.260 ;
        RECT 2133.565 18.075 2133.855 18.120 ;
        RECT 2146.430 18.060 2146.750 18.120 ;
        RECT 1947.250 17.920 1947.570 17.980 ;
        RECT 2090.785 17.920 2091.075 17.965 ;
        RECT 1947.250 17.780 2091.075 17.920 ;
        RECT 1947.250 17.720 1947.570 17.780 ;
        RECT 2090.785 17.735 2091.075 17.780 ;
        RECT 2090.785 14.520 2091.075 14.565 ;
        RECT 2133.565 14.520 2133.855 14.565 ;
        RECT 2090.785 14.380 2133.855 14.520 ;
        RECT 2090.785 14.335 2091.075 14.380 ;
        RECT 2133.565 14.335 2133.855 14.380 ;
      LAYER via ;
        RECT 2146.460 18.060 2146.720 18.320 ;
        RECT 1947.280 17.720 1947.540 17.980 ;
      LAYER met2 ;
        RECT 2150.980 1700.410 2151.260 1704.000 ;
        RECT 2148.820 1700.270 2151.260 1700.410 ;
        RECT 2148.820 1656.210 2148.960 1700.270 ;
        RECT 2150.980 1700.000 2151.260 1700.270 ;
        RECT 2146.520 1656.070 2148.960 1656.210 ;
        RECT 2146.520 18.350 2146.660 1656.070 ;
        RECT 2146.460 18.030 2146.720 18.350 ;
        RECT 1947.280 17.690 1947.540 18.010 ;
        RECT 1947.340 2.400 1947.480 17.690 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1966.185 1594.005 1966.355 1642.115 ;
        RECT 1966.185 724.965 1966.355 814.215 ;
        RECT 1966.185 669.545 1966.355 717.655 ;
        RECT 1965.725 493.425 1965.895 524.195 ;
        RECT 1966.185 89.845 1966.355 137.955 ;
        RECT 1965.265 2.805 1965.435 48.195 ;
      LAYER mcon ;
        RECT 1966.185 1641.945 1966.355 1642.115 ;
        RECT 1966.185 814.045 1966.355 814.215 ;
        RECT 1966.185 717.485 1966.355 717.655 ;
        RECT 1965.725 524.025 1965.895 524.195 ;
        RECT 1966.185 137.785 1966.355 137.955 ;
        RECT 1965.265 48.025 1965.435 48.195 ;
      LAYER met1 ;
        RECT 1966.110 1688.000 1966.430 1688.060 ;
        RECT 2160.230 1688.000 2160.550 1688.060 ;
        RECT 1966.110 1687.860 2160.550 1688.000 ;
        RECT 1966.110 1687.800 1966.430 1687.860 ;
        RECT 2160.230 1687.800 2160.550 1687.860 ;
        RECT 1966.110 1642.100 1966.430 1642.160 ;
        RECT 1965.915 1641.960 1966.430 1642.100 ;
        RECT 1966.110 1641.900 1966.430 1641.960 ;
        RECT 1966.110 1594.160 1966.430 1594.220 ;
        RECT 1965.915 1594.020 1966.430 1594.160 ;
        RECT 1966.110 1593.960 1966.430 1594.020 ;
        RECT 1966.110 1345.620 1966.430 1345.680 ;
        RECT 1967.030 1345.620 1967.350 1345.680 ;
        RECT 1966.110 1345.480 1967.350 1345.620 ;
        RECT 1966.110 1345.420 1966.430 1345.480 ;
        RECT 1967.030 1345.420 1967.350 1345.480 ;
        RECT 1966.110 1297.340 1966.430 1297.400 ;
        RECT 1967.030 1297.340 1967.350 1297.400 ;
        RECT 1966.110 1297.200 1967.350 1297.340 ;
        RECT 1966.110 1297.140 1966.430 1297.200 ;
        RECT 1967.030 1297.140 1967.350 1297.200 ;
        RECT 1966.110 1256.540 1966.430 1256.600 ;
        RECT 1965.740 1256.400 1966.430 1256.540 ;
        RECT 1965.740 1255.580 1965.880 1256.400 ;
        RECT 1966.110 1256.340 1966.430 1256.400 ;
        RECT 1965.650 1255.320 1965.970 1255.580 ;
        RECT 1964.730 1200.780 1965.050 1200.840 ;
        RECT 1966.110 1200.780 1966.430 1200.840 ;
        RECT 1964.730 1200.640 1966.430 1200.780 ;
        RECT 1964.730 1200.580 1965.050 1200.640 ;
        RECT 1966.110 1200.580 1966.430 1200.640 ;
        RECT 1966.110 821.140 1966.430 821.400 ;
        RECT 1966.200 820.720 1966.340 821.140 ;
        RECT 1966.110 820.460 1966.430 820.720 ;
        RECT 1966.110 814.200 1966.430 814.260 ;
        RECT 1965.915 814.060 1966.430 814.200 ;
        RECT 1966.110 814.000 1966.430 814.060 ;
        RECT 1966.110 725.120 1966.430 725.180 ;
        RECT 1965.915 724.980 1966.430 725.120 ;
        RECT 1966.110 724.920 1966.430 724.980 ;
        RECT 1966.110 717.640 1966.430 717.700 ;
        RECT 1965.915 717.500 1966.430 717.640 ;
        RECT 1966.110 717.440 1966.430 717.500 ;
        RECT 1966.110 669.700 1966.430 669.760 ;
        RECT 1965.915 669.560 1966.430 669.700 ;
        RECT 1966.110 669.500 1966.430 669.560 ;
        RECT 1966.110 573.280 1966.430 573.540 ;
        RECT 1966.200 572.860 1966.340 573.280 ;
        RECT 1966.110 572.600 1966.430 572.860 ;
        RECT 1965.665 524.180 1965.955 524.225 ;
        RECT 1966.110 524.180 1966.430 524.240 ;
        RECT 1965.665 524.040 1966.430 524.180 ;
        RECT 1965.665 523.995 1965.955 524.040 ;
        RECT 1966.110 523.980 1966.430 524.040 ;
        RECT 1965.650 493.580 1965.970 493.640 ;
        RECT 1965.455 493.440 1965.970 493.580 ;
        RECT 1965.650 493.380 1965.970 493.440 ;
        RECT 1966.110 331.060 1966.430 331.120 ;
        RECT 1965.740 330.920 1966.430 331.060 ;
        RECT 1965.740 330.780 1965.880 330.920 ;
        RECT 1966.110 330.860 1966.430 330.920 ;
        RECT 1965.650 330.520 1965.970 330.780 ;
        RECT 1965.650 241.640 1965.970 241.700 ;
        RECT 1966.110 241.640 1966.430 241.700 ;
        RECT 1965.650 241.500 1966.430 241.640 ;
        RECT 1965.650 241.440 1965.970 241.500 ;
        RECT 1966.110 241.440 1966.430 241.500 ;
        RECT 1965.650 145.080 1965.970 145.140 ;
        RECT 1966.110 145.080 1966.430 145.140 ;
        RECT 1965.650 144.940 1966.430 145.080 ;
        RECT 1965.650 144.880 1965.970 144.940 ;
        RECT 1966.110 144.880 1966.430 144.940 ;
        RECT 1966.110 137.940 1966.430 138.000 ;
        RECT 1965.915 137.800 1966.430 137.940 ;
        RECT 1966.110 137.740 1966.430 137.800 ;
        RECT 1966.110 90.000 1966.430 90.060 ;
        RECT 1965.915 89.860 1966.430 90.000 ;
        RECT 1966.110 89.800 1966.430 89.860 ;
        RECT 1966.110 62.460 1966.430 62.520 ;
        RECT 1965.280 62.320 1966.430 62.460 ;
        RECT 1965.280 62.180 1965.420 62.320 ;
        RECT 1966.110 62.260 1966.430 62.320 ;
        RECT 1965.190 61.920 1965.510 62.180 ;
        RECT 1965.190 48.180 1965.510 48.240 ;
        RECT 1964.995 48.040 1965.510 48.180 ;
        RECT 1965.190 47.980 1965.510 48.040 ;
        RECT 1965.190 2.960 1965.510 3.020 ;
        RECT 1964.995 2.820 1965.510 2.960 ;
        RECT 1965.190 2.760 1965.510 2.820 ;
      LAYER via ;
        RECT 1966.140 1687.800 1966.400 1688.060 ;
        RECT 2160.260 1687.800 2160.520 1688.060 ;
        RECT 1966.140 1641.900 1966.400 1642.160 ;
        RECT 1966.140 1593.960 1966.400 1594.220 ;
        RECT 1966.140 1345.420 1966.400 1345.680 ;
        RECT 1967.060 1345.420 1967.320 1345.680 ;
        RECT 1966.140 1297.140 1966.400 1297.400 ;
        RECT 1967.060 1297.140 1967.320 1297.400 ;
        RECT 1966.140 1256.340 1966.400 1256.600 ;
        RECT 1965.680 1255.320 1965.940 1255.580 ;
        RECT 1964.760 1200.580 1965.020 1200.840 ;
        RECT 1966.140 1200.580 1966.400 1200.840 ;
        RECT 1966.140 821.140 1966.400 821.400 ;
        RECT 1966.140 820.460 1966.400 820.720 ;
        RECT 1966.140 814.000 1966.400 814.260 ;
        RECT 1966.140 724.920 1966.400 725.180 ;
        RECT 1966.140 717.440 1966.400 717.700 ;
        RECT 1966.140 669.500 1966.400 669.760 ;
        RECT 1966.140 573.280 1966.400 573.540 ;
        RECT 1966.140 572.600 1966.400 572.860 ;
        RECT 1966.140 523.980 1966.400 524.240 ;
        RECT 1965.680 493.380 1965.940 493.640 ;
        RECT 1966.140 330.860 1966.400 331.120 ;
        RECT 1965.680 330.520 1965.940 330.780 ;
        RECT 1965.680 241.440 1965.940 241.700 ;
        RECT 1966.140 241.440 1966.400 241.700 ;
        RECT 1965.680 144.880 1965.940 145.140 ;
        RECT 1966.140 144.880 1966.400 145.140 ;
        RECT 1966.140 137.740 1966.400 138.000 ;
        RECT 1966.140 89.800 1966.400 90.060 ;
        RECT 1966.140 62.260 1966.400 62.520 ;
        RECT 1965.220 61.920 1965.480 62.180 ;
        RECT 1965.220 47.980 1965.480 48.240 ;
        RECT 1965.220 2.760 1965.480 3.020 ;
      LAYER met2 ;
        RECT 2160.180 1700.000 2160.460 1704.000 ;
        RECT 2160.320 1688.090 2160.460 1700.000 ;
        RECT 1966.140 1687.770 1966.400 1688.090 ;
        RECT 2160.260 1687.770 2160.520 1688.090 ;
        RECT 1966.200 1642.190 1966.340 1687.770 ;
        RECT 1966.140 1641.870 1966.400 1642.190 ;
        RECT 1966.140 1593.930 1966.400 1594.250 ;
        RECT 1966.200 1393.845 1966.340 1593.930 ;
        RECT 1966.130 1393.475 1966.410 1393.845 ;
        RECT 1967.050 1393.475 1967.330 1393.845 ;
        RECT 1967.120 1345.710 1967.260 1393.475 ;
        RECT 1966.140 1345.565 1966.400 1345.710 ;
        RECT 1967.060 1345.565 1967.320 1345.710 ;
        RECT 1966.130 1345.195 1966.410 1345.565 ;
        RECT 1967.050 1345.195 1967.330 1345.565 ;
        RECT 1967.120 1297.430 1967.260 1345.195 ;
        RECT 1966.140 1297.110 1966.400 1297.430 ;
        RECT 1967.060 1297.110 1967.320 1297.430 ;
        RECT 1966.200 1256.630 1966.340 1297.110 ;
        RECT 1966.140 1256.310 1966.400 1256.630 ;
        RECT 1965.680 1255.290 1965.940 1255.610 ;
        RECT 1965.740 1249.005 1965.880 1255.290 ;
        RECT 1964.750 1248.635 1965.030 1249.005 ;
        RECT 1965.670 1248.635 1965.950 1249.005 ;
        RECT 1964.820 1200.870 1964.960 1248.635 ;
        RECT 1964.760 1200.550 1965.020 1200.870 ;
        RECT 1966.140 1200.550 1966.400 1200.870 ;
        RECT 1966.200 821.430 1966.340 1200.550 ;
        RECT 1966.140 821.110 1966.400 821.430 ;
        RECT 1966.140 820.430 1966.400 820.750 ;
        RECT 1966.200 814.290 1966.340 820.430 ;
        RECT 1966.140 813.970 1966.400 814.290 ;
        RECT 1966.140 724.890 1966.400 725.210 ;
        RECT 1966.200 717.730 1966.340 724.890 ;
        RECT 1966.140 717.410 1966.400 717.730 ;
        RECT 1966.140 669.470 1966.400 669.790 ;
        RECT 1966.200 628.845 1966.340 669.470 ;
        RECT 1966.130 628.475 1966.410 628.845 ;
        RECT 1966.130 627.795 1966.410 628.165 ;
        RECT 1966.200 573.570 1966.340 627.795 ;
        RECT 1966.140 573.250 1966.400 573.570 ;
        RECT 1966.140 572.570 1966.400 572.890 ;
        RECT 1966.200 524.270 1966.340 572.570 ;
        RECT 1966.140 523.950 1966.400 524.270 ;
        RECT 1965.680 493.350 1965.940 493.670 ;
        RECT 1965.740 434.250 1965.880 493.350 ;
        RECT 1965.740 434.110 1966.340 434.250 ;
        RECT 1966.200 331.150 1966.340 434.110 ;
        RECT 1966.140 330.830 1966.400 331.150 ;
        RECT 1965.680 330.490 1965.940 330.810 ;
        RECT 1965.740 241.730 1965.880 330.490 ;
        RECT 1965.680 241.410 1965.940 241.730 ;
        RECT 1966.140 241.410 1966.400 241.730 ;
        RECT 1966.200 195.570 1966.340 241.410 ;
        RECT 1965.740 195.430 1966.340 195.570 ;
        RECT 1965.740 145.170 1965.880 195.430 ;
        RECT 1965.680 144.850 1965.940 145.170 ;
        RECT 1966.140 144.850 1966.400 145.170 ;
        RECT 1966.200 138.030 1966.340 144.850 ;
        RECT 1966.140 137.710 1966.400 138.030 ;
        RECT 1966.140 89.770 1966.400 90.090 ;
        RECT 1966.200 62.550 1966.340 89.770 ;
        RECT 1966.140 62.230 1966.400 62.550 ;
        RECT 1965.220 61.890 1965.480 62.210 ;
        RECT 1965.280 48.270 1965.420 61.890 ;
        RECT 1965.220 47.950 1965.480 48.270 ;
        RECT 1965.220 2.730 1965.480 3.050 ;
        RECT 1965.280 2.400 1965.420 2.730 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
      LAYER via2 ;
        RECT 1966.130 1393.520 1966.410 1393.800 ;
        RECT 1967.050 1393.520 1967.330 1393.800 ;
        RECT 1966.130 1345.240 1966.410 1345.520 ;
        RECT 1967.050 1345.240 1967.330 1345.520 ;
        RECT 1964.750 1248.680 1965.030 1248.960 ;
        RECT 1965.670 1248.680 1965.950 1248.960 ;
        RECT 1966.130 628.520 1966.410 628.800 ;
        RECT 1966.130 627.840 1966.410 628.120 ;
      LAYER met3 ;
        RECT 1966.105 1393.810 1966.435 1393.825 ;
        RECT 1967.025 1393.810 1967.355 1393.825 ;
        RECT 1966.105 1393.510 1967.355 1393.810 ;
        RECT 1966.105 1393.495 1966.435 1393.510 ;
        RECT 1967.025 1393.495 1967.355 1393.510 ;
        RECT 1966.105 1345.530 1966.435 1345.545 ;
        RECT 1967.025 1345.530 1967.355 1345.545 ;
        RECT 1966.105 1345.230 1967.355 1345.530 ;
        RECT 1966.105 1345.215 1966.435 1345.230 ;
        RECT 1967.025 1345.215 1967.355 1345.230 ;
        RECT 1964.725 1248.970 1965.055 1248.985 ;
        RECT 1965.645 1248.970 1965.975 1248.985 ;
        RECT 1964.725 1248.670 1965.975 1248.970 ;
        RECT 1964.725 1248.655 1965.055 1248.670 ;
        RECT 1965.645 1248.655 1965.975 1248.670 ;
        RECT 1966.105 628.810 1966.435 628.825 ;
        RECT 1966.105 628.495 1966.650 628.810 ;
        RECT 1966.350 628.145 1966.650 628.495 ;
        RECT 1966.105 627.830 1966.650 628.145 ;
        RECT 1966.105 627.815 1966.435 627.830 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2018.625 16.915 2018.795 18.615 ;
        RECT 2018.165 16.745 2018.795 16.915 ;
      LAYER mcon ;
        RECT 2018.625 18.445 2018.795 18.615 ;
      LAYER met1 ;
        RECT 2018.565 18.600 2018.855 18.645 ;
        RECT 2166.670 18.600 2166.990 18.660 ;
        RECT 2018.565 18.460 2166.990 18.600 ;
        RECT 2018.565 18.415 2018.855 18.460 ;
        RECT 2166.670 18.400 2166.990 18.460 ;
        RECT 1983.130 16.900 1983.450 16.960 ;
        RECT 2018.105 16.900 2018.395 16.945 ;
        RECT 1983.130 16.760 2018.395 16.900 ;
        RECT 1983.130 16.700 1983.450 16.760 ;
        RECT 2018.105 16.715 2018.395 16.760 ;
      LAYER via ;
        RECT 2166.700 18.400 2166.960 18.660 ;
        RECT 1983.160 16.700 1983.420 16.960 ;
      LAYER met2 ;
        RECT 2169.380 1700.410 2169.660 1704.000 ;
        RECT 2166.760 1700.270 2169.660 1700.410 ;
        RECT 2166.760 18.690 2166.900 1700.270 ;
        RECT 2169.380 1700.000 2169.660 1700.270 ;
        RECT 2166.700 18.370 2166.960 18.690 ;
        RECT 1983.160 16.670 1983.420 16.990 ;
        RECT 1983.220 2.400 1983.360 16.670 ;
        RECT 1983.010 -4.800 1983.570 2.400 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2162.990 1687.660 2163.310 1687.720 ;
        RECT 2178.630 1687.660 2178.950 1687.720 ;
        RECT 2162.990 1687.520 2178.950 1687.660 ;
        RECT 2162.990 1687.460 2163.310 1687.520 ;
        RECT 2178.630 1687.460 2178.950 1687.520 ;
        RECT 2001.070 19.620 2001.390 19.680 ;
        RECT 2162.070 19.620 2162.390 19.680 ;
        RECT 2001.070 19.480 2162.390 19.620 ;
        RECT 2001.070 19.420 2001.390 19.480 ;
        RECT 2162.070 19.420 2162.390 19.480 ;
      LAYER via ;
        RECT 2163.020 1687.460 2163.280 1687.720 ;
        RECT 2178.660 1687.460 2178.920 1687.720 ;
        RECT 2001.100 19.420 2001.360 19.680 ;
        RECT 2162.100 19.420 2162.360 19.680 ;
      LAYER met2 ;
        RECT 2178.580 1700.000 2178.860 1704.000 ;
        RECT 2178.720 1687.750 2178.860 1700.000 ;
        RECT 2163.020 1687.430 2163.280 1687.750 ;
        RECT 2178.660 1687.430 2178.920 1687.750 ;
        RECT 2001.100 19.390 2001.360 19.710 ;
        RECT 2162.100 19.450 2162.360 19.710 ;
        RECT 2163.080 19.450 2163.220 1687.430 ;
        RECT 2162.100 19.390 2163.220 19.450 ;
        RECT 2001.160 2.400 2001.300 19.390 ;
        RECT 2162.160 19.310 2163.220 19.390 ;
        RECT 2000.950 -4.800 2001.510 2.400 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2018.550 19.280 2018.870 19.340 ;
        RECT 2188.290 19.280 2188.610 19.340 ;
        RECT 2018.550 19.140 2188.610 19.280 ;
        RECT 2018.550 19.080 2018.870 19.140 ;
        RECT 2188.290 19.080 2188.610 19.140 ;
      LAYER via ;
        RECT 2018.580 19.080 2018.840 19.340 ;
        RECT 2188.320 19.080 2188.580 19.340 ;
      LAYER met2 ;
        RECT 2187.780 1700.410 2188.060 1704.000 ;
        RECT 2187.780 1700.270 2188.520 1700.410 ;
        RECT 2187.780 1700.000 2188.060 1700.270 ;
        RECT 2188.380 19.370 2188.520 1700.270 ;
        RECT 2018.580 19.050 2018.840 19.370 ;
        RECT 2188.320 19.050 2188.580 19.370 ;
        RECT 2018.640 2.400 2018.780 19.050 ;
        RECT 2018.430 -4.800 2018.990 2.400 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2048.065 17.085 2049.615 17.255 ;
        RECT 2081.185 17.085 2081.355 20.315 ;
        RECT 2048.065 16.745 2048.235 17.085 ;
      LAYER mcon ;
        RECT 2081.185 20.145 2081.355 20.315 ;
        RECT 2049.445 17.085 2049.615 17.255 ;
      LAYER met1 ;
        RECT 2081.125 20.300 2081.415 20.345 ;
        RECT 2194.730 20.300 2195.050 20.360 ;
        RECT 2081.125 20.160 2195.050 20.300 ;
        RECT 2081.125 20.115 2081.415 20.160 ;
        RECT 2194.730 20.100 2195.050 20.160 ;
        RECT 2049.385 17.240 2049.675 17.285 ;
        RECT 2081.125 17.240 2081.415 17.285 ;
        RECT 2049.385 17.100 2081.415 17.240 ;
        RECT 2049.385 17.055 2049.675 17.100 ;
        RECT 2081.125 17.055 2081.415 17.100 ;
        RECT 2036.490 16.900 2036.810 16.960 ;
        RECT 2048.005 16.900 2048.295 16.945 ;
        RECT 2036.490 16.760 2048.295 16.900 ;
        RECT 2036.490 16.700 2036.810 16.760 ;
        RECT 2048.005 16.715 2048.295 16.760 ;
      LAYER via ;
        RECT 2194.760 20.100 2195.020 20.360 ;
        RECT 2036.520 16.700 2036.780 16.960 ;
      LAYER met2 ;
        RECT 2196.980 1700.410 2197.260 1704.000 ;
        RECT 2194.820 1700.270 2197.260 1700.410 ;
        RECT 2194.820 20.390 2194.960 1700.270 ;
        RECT 2196.980 1700.000 2197.260 1700.270 ;
        RECT 2194.760 20.070 2195.020 20.390 ;
        RECT 2036.520 16.670 2036.780 16.990 ;
        RECT 2036.580 2.400 2036.720 16.670 ;
        RECT 2036.370 -4.800 2036.930 2.400 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2114.765 1684.445 2114.935 1689.715 ;
        RECT 2162.605 1687.845 2162.775 1689.715 ;
      LAYER mcon ;
        RECT 2114.765 1689.545 2114.935 1689.715 ;
        RECT 2162.605 1689.545 2162.775 1689.715 ;
      LAYER met1 ;
        RECT 2114.705 1689.700 2114.995 1689.745 ;
        RECT 2162.545 1689.700 2162.835 1689.745 ;
        RECT 2114.705 1689.560 2162.835 1689.700 ;
        RECT 2114.705 1689.515 2114.995 1689.560 ;
        RECT 2162.545 1689.515 2162.835 1689.560 ;
        RECT 2162.545 1688.000 2162.835 1688.045 ;
        RECT 2206.230 1688.000 2206.550 1688.060 ;
        RECT 2162.545 1687.860 2206.550 1688.000 ;
        RECT 2162.545 1687.815 2162.835 1687.860 ;
        RECT 2206.230 1687.800 2206.550 1687.860 ;
        RECT 2066.850 1684.600 2067.170 1684.660 ;
        RECT 2114.705 1684.600 2114.995 1684.645 ;
        RECT 2066.850 1684.460 2114.995 1684.600 ;
        RECT 2066.850 1684.400 2067.170 1684.460 ;
        RECT 2114.705 1684.415 2114.995 1684.460 ;
        RECT 2054.430 20.300 2054.750 20.360 ;
        RECT 2066.850 20.300 2067.170 20.360 ;
        RECT 2054.430 20.160 2067.170 20.300 ;
        RECT 2054.430 20.100 2054.750 20.160 ;
        RECT 2066.850 20.100 2067.170 20.160 ;
      LAYER via ;
        RECT 2206.260 1687.800 2206.520 1688.060 ;
        RECT 2066.880 1684.400 2067.140 1684.660 ;
        RECT 2054.460 20.100 2054.720 20.360 ;
        RECT 2066.880 20.100 2067.140 20.360 ;
      LAYER met2 ;
        RECT 2206.180 1700.000 2206.460 1704.000 ;
        RECT 2206.320 1688.090 2206.460 1700.000 ;
        RECT 2206.260 1687.770 2206.520 1688.090 ;
        RECT 2066.880 1684.370 2067.140 1684.690 ;
        RECT 2066.940 20.390 2067.080 1684.370 ;
        RECT 2054.460 20.070 2054.720 20.390 ;
        RECT 2066.880 20.070 2067.140 20.390 ;
        RECT 2054.520 2.400 2054.660 20.070 ;
        RECT 2054.310 -4.800 2054.870 2.400 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1540.685 483.225 1540.855 496.995 ;
        RECT 1540.685 386.325 1540.855 434.775 ;
        RECT 1540.225 50.405 1540.395 96.475 ;
      LAYER mcon ;
        RECT 1540.685 496.825 1540.855 496.995 ;
        RECT 1540.685 434.605 1540.855 434.775 ;
        RECT 1540.225 96.305 1540.395 96.475 ;
      LAYER met1 ;
        RECT 1540.610 1062.740 1540.930 1062.800 ;
        RECT 1541.530 1062.740 1541.850 1062.800 ;
        RECT 1540.610 1062.600 1541.850 1062.740 ;
        RECT 1540.610 1062.540 1540.930 1062.600 ;
        RECT 1541.530 1062.540 1541.850 1062.600 ;
        RECT 1540.610 966.180 1540.930 966.240 ;
        RECT 1541.530 966.180 1541.850 966.240 ;
        RECT 1540.610 966.040 1541.850 966.180 ;
        RECT 1540.610 965.980 1540.930 966.040 ;
        RECT 1541.530 965.980 1541.850 966.040 ;
        RECT 1540.610 869.620 1540.930 869.680 ;
        RECT 1541.070 869.620 1541.390 869.680 ;
        RECT 1540.610 869.480 1541.390 869.620 ;
        RECT 1540.610 869.420 1540.930 869.480 ;
        RECT 1541.070 869.420 1541.390 869.480 ;
        RECT 1540.150 821.000 1540.470 821.060 ;
        RECT 1541.070 821.000 1541.390 821.060 ;
        RECT 1540.150 820.860 1541.390 821.000 ;
        RECT 1540.150 820.800 1540.470 820.860 ;
        RECT 1541.070 820.800 1541.390 820.860 ;
        RECT 1541.070 814.200 1541.390 814.260 ;
        RECT 1541.990 814.200 1542.310 814.260 ;
        RECT 1541.070 814.060 1542.310 814.200 ;
        RECT 1541.070 814.000 1541.390 814.060 ;
        RECT 1541.990 814.000 1542.310 814.060 ;
        RECT 1540.610 724.780 1540.930 724.840 ;
        RECT 1541.070 724.780 1541.390 724.840 ;
        RECT 1540.610 724.640 1541.390 724.780 ;
        RECT 1540.610 724.580 1540.930 724.640 ;
        RECT 1541.070 724.580 1541.390 724.640 ;
        RECT 1540.610 593.340 1540.930 593.600 ;
        RECT 1540.700 592.920 1540.840 593.340 ;
        RECT 1540.610 592.660 1540.930 592.920 ;
        RECT 1540.610 496.980 1540.930 497.040 ;
        RECT 1540.415 496.840 1540.930 496.980 ;
        RECT 1540.610 496.780 1540.930 496.840 ;
        RECT 1540.610 483.380 1540.930 483.440 ;
        RECT 1540.415 483.240 1540.930 483.380 ;
        RECT 1540.610 483.180 1540.930 483.240 ;
        RECT 1540.610 434.760 1540.930 434.820 ;
        RECT 1540.415 434.620 1540.930 434.760 ;
        RECT 1540.610 434.560 1540.930 434.620 ;
        RECT 1540.610 386.480 1540.930 386.540 ;
        RECT 1540.415 386.340 1540.930 386.480 ;
        RECT 1540.610 386.280 1540.930 386.340 ;
        RECT 1540.150 289.920 1540.470 289.980 ;
        RECT 1540.610 289.920 1540.930 289.980 ;
        RECT 1540.150 289.780 1540.930 289.920 ;
        RECT 1540.150 289.720 1540.470 289.780 ;
        RECT 1540.610 289.720 1540.930 289.780 ;
        RECT 1540.150 96.460 1540.470 96.520 ;
        RECT 1539.955 96.320 1540.470 96.460 ;
        RECT 1540.150 96.260 1540.470 96.320 ;
        RECT 772.410 50.560 772.730 50.620 ;
        RECT 1540.165 50.560 1540.455 50.605 ;
        RECT 772.410 50.420 1540.455 50.560 ;
        RECT 772.410 50.360 772.730 50.420 ;
        RECT 1540.165 50.375 1540.455 50.420 ;
      LAYER via ;
        RECT 1540.640 1062.540 1540.900 1062.800 ;
        RECT 1541.560 1062.540 1541.820 1062.800 ;
        RECT 1540.640 965.980 1540.900 966.240 ;
        RECT 1541.560 965.980 1541.820 966.240 ;
        RECT 1540.640 869.420 1540.900 869.680 ;
        RECT 1541.100 869.420 1541.360 869.680 ;
        RECT 1540.180 820.800 1540.440 821.060 ;
        RECT 1541.100 820.800 1541.360 821.060 ;
        RECT 1541.100 814.000 1541.360 814.260 ;
        RECT 1542.020 814.000 1542.280 814.260 ;
        RECT 1540.640 724.580 1540.900 724.840 ;
        RECT 1541.100 724.580 1541.360 724.840 ;
        RECT 1540.640 593.340 1540.900 593.600 ;
        RECT 1540.640 592.660 1540.900 592.920 ;
        RECT 1540.640 496.780 1540.900 497.040 ;
        RECT 1540.640 483.180 1540.900 483.440 ;
        RECT 1540.640 434.560 1540.900 434.820 ;
        RECT 1540.640 386.280 1540.900 386.540 ;
        RECT 1540.180 289.720 1540.440 289.980 ;
        RECT 1540.640 289.720 1540.900 289.980 ;
        RECT 1540.180 96.260 1540.440 96.520 ;
        RECT 772.440 50.360 772.700 50.620 ;
      LAYER met2 ;
        RECT 1544.700 1700.410 1544.980 1704.000 ;
        RECT 1542.540 1700.270 1544.980 1700.410 ;
        RECT 1542.540 1656.210 1542.680 1700.270 ;
        RECT 1544.700 1700.000 1544.980 1700.270 ;
        RECT 1540.240 1656.070 1542.680 1656.210 ;
        RECT 1540.240 1110.965 1540.380 1656.070 ;
        RECT 1540.170 1110.595 1540.450 1110.965 ;
        RECT 1541.550 1110.595 1541.830 1110.965 ;
        RECT 1541.620 1062.830 1541.760 1110.595 ;
        RECT 1540.640 1062.510 1540.900 1062.830 ;
        RECT 1541.560 1062.510 1541.820 1062.830 ;
        RECT 1540.700 1014.405 1540.840 1062.510 ;
        RECT 1540.630 1014.035 1540.910 1014.405 ;
        RECT 1541.550 1014.035 1541.830 1014.405 ;
        RECT 1541.620 966.270 1541.760 1014.035 ;
        RECT 1540.640 965.950 1540.900 966.270 ;
        RECT 1541.560 965.950 1541.820 966.270 ;
        RECT 1540.700 883.050 1540.840 965.950 ;
        RECT 1540.700 882.910 1541.300 883.050 ;
        RECT 1541.160 869.710 1541.300 882.910 ;
        RECT 1540.640 869.390 1540.900 869.710 ;
        RECT 1541.100 869.390 1541.360 869.710 ;
        RECT 1540.700 845.650 1540.840 869.390 ;
        RECT 1540.240 845.510 1540.840 845.650 ;
        RECT 1540.240 821.090 1540.380 845.510 ;
        RECT 1540.180 820.770 1540.440 821.090 ;
        RECT 1541.100 820.770 1541.360 821.090 ;
        RECT 1541.160 814.290 1541.300 820.770 ;
        RECT 1541.100 813.970 1541.360 814.290 ;
        RECT 1542.020 813.970 1542.280 814.290 ;
        RECT 1542.080 766.205 1542.220 813.970 ;
        RECT 1541.090 765.835 1541.370 766.205 ;
        RECT 1542.010 765.835 1542.290 766.205 ;
        RECT 1541.160 724.870 1541.300 765.835 ;
        RECT 1540.640 724.550 1540.900 724.870 ;
        RECT 1541.100 724.550 1541.360 724.870 ;
        RECT 1540.700 690.610 1540.840 724.550 ;
        RECT 1540.240 690.470 1540.840 690.610 ;
        RECT 1540.240 689.930 1540.380 690.470 ;
        RECT 1540.240 689.790 1540.840 689.930 ;
        RECT 1540.700 593.630 1540.840 689.790 ;
        RECT 1540.640 593.310 1540.900 593.630 ;
        RECT 1540.640 592.630 1540.900 592.950 ;
        RECT 1540.700 497.070 1540.840 592.630 ;
        RECT 1540.640 496.750 1540.900 497.070 ;
        RECT 1540.640 483.150 1540.900 483.470 ;
        RECT 1540.700 434.850 1540.840 483.150 ;
        RECT 1540.640 434.530 1540.900 434.850 ;
        RECT 1540.640 386.250 1540.900 386.570 ;
        RECT 1540.700 290.010 1540.840 386.250 ;
        RECT 1540.180 289.690 1540.440 290.010 ;
        RECT 1540.640 289.690 1540.900 290.010 ;
        RECT 1540.240 254.730 1540.380 289.690 ;
        RECT 1540.240 254.590 1540.840 254.730 ;
        RECT 1540.700 109.890 1540.840 254.590 ;
        RECT 1540.240 109.750 1540.840 109.890 ;
        RECT 1540.240 96.550 1540.380 109.750 ;
        RECT 1540.180 96.230 1540.440 96.550 ;
        RECT 772.440 50.330 772.700 50.650 ;
        RECT 772.500 16.730 772.640 50.330 ;
        RECT 769.740 16.590 772.640 16.730 ;
        RECT 769.740 2.400 769.880 16.590 ;
        RECT 769.530 -4.800 770.090 2.400 ;
      LAYER via2 ;
        RECT 1540.170 1110.640 1540.450 1110.920 ;
        RECT 1541.550 1110.640 1541.830 1110.920 ;
        RECT 1540.630 1014.080 1540.910 1014.360 ;
        RECT 1541.550 1014.080 1541.830 1014.360 ;
        RECT 1541.090 765.880 1541.370 766.160 ;
        RECT 1542.010 765.880 1542.290 766.160 ;
      LAYER met3 ;
        RECT 1540.145 1110.930 1540.475 1110.945 ;
        RECT 1541.525 1110.930 1541.855 1110.945 ;
        RECT 1540.145 1110.630 1541.855 1110.930 ;
        RECT 1540.145 1110.615 1540.475 1110.630 ;
        RECT 1541.525 1110.615 1541.855 1110.630 ;
        RECT 1540.605 1014.370 1540.935 1014.385 ;
        RECT 1541.525 1014.370 1541.855 1014.385 ;
        RECT 1540.605 1014.070 1541.855 1014.370 ;
        RECT 1540.605 1014.055 1540.935 1014.070 ;
        RECT 1541.525 1014.055 1541.855 1014.070 ;
        RECT 1541.065 766.170 1541.395 766.185 ;
        RECT 1541.985 766.170 1542.315 766.185 ;
        RECT 1541.065 765.870 1542.315 766.170 ;
        RECT 1541.065 765.855 1541.395 765.870 ;
        RECT 1541.985 765.855 1542.315 765.870 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2080.650 1689.360 2080.970 1689.420 ;
        RECT 2214.970 1689.360 2215.290 1689.420 ;
        RECT 2080.650 1689.220 2215.290 1689.360 ;
        RECT 2080.650 1689.160 2080.970 1689.220 ;
        RECT 2214.970 1689.160 2215.290 1689.220 ;
        RECT 2072.370 20.300 2072.690 20.360 ;
        RECT 2080.650 20.300 2080.970 20.360 ;
        RECT 2072.370 20.160 2080.970 20.300 ;
        RECT 2072.370 20.100 2072.690 20.160 ;
        RECT 2080.650 20.100 2080.970 20.160 ;
      LAYER via ;
        RECT 2080.680 1689.160 2080.940 1689.420 ;
        RECT 2215.000 1689.160 2215.260 1689.420 ;
        RECT 2072.400 20.100 2072.660 20.360 ;
        RECT 2080.680 20.100 2080.940 20.360 ;
      LAYER met2 ;
        RECT 2214.920 1700.000 2215.200 1704.000 ;
        RECT 2215.060 1689.450 2215.200 1700.000 ;
        RECT 2080.680 1689.130 2080.940 1689.450 ;
        RECT 2215.000 1689.130 2215.260 1689.450 ;
        RECT 2080.740 20.390 2080.880 1689.130 ;
        RECT 2072.400 20.070 2072.660 20.390 ;
        RECT 2080.680 20.070 2080.940 20.390 ;
        RECT 2072.460 2.400 2072.600 20.070 ;
        RECT 2072.250 -4.800 2072.810 2.400 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2222.790 17.240 2223.110 17.300 ;
        RECT 2110.180 17.100 2223.110 17.240 ;
        RECT 2089.850 16.560 2090.170 16.620 ;
        RECT 2110.180 16.560 2110.320 17.100 ;
        RECT 2222.790 17.040 2223.110 17.100 ;
        RECT 2089.850 16.420 2110.320 16.560 ;
        RECT 2089.850 16.360 2090.170 16.420 ;
      LAYER via ;
        RECT 2089.880 16.360 2090.140 16.620 ;
        RECT 2222.820 17.040 2223.080 17.300 ;
      LAYER met2 ;
        RECT 2224.120 1700.410 2224.400 1704.000 ;
        RECT 2222.880 1700.270 2224.400 1700.410 ;
        RECT 2222.880 17.330 2223.020 1700.270 ;
        RECT 2224.120 1700.000 2224.400 1700.270 ;
        RECT 2222.820 17.010 2223.080 17.330 ;
        RECT 2089.880 16.330 2090.140 16.650 ;
        RECT 2089.940 2.400 2090.080 16.330 ;
        RECT 2089.730 -4.800 2090.290 2.400 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2115.225 1686.145 2115.395 1687.335 ;
      LAYER mcon ;
        RECT 2115.225 1687.165 2115.395 1687.335 ;
      LAYER met1 ;
        RECT 2115.165 1687.320 2115.455 1687.365 ;
        RECT 2231.990 1687.320 2232.310 1687.380 ;
        RECT 2115.165 1687.180 2232.310 1687.320 ;
        RECT 2115.165 1687.135 2115.455 1687.180 ;
        RECT 2231.990 1687.120 2232.310 1687.180 ;
        RECT 2111.010 1686.300 2111.330 1686.360 ;
        RECT 2115.165 1686.300 2115.455 1686.345 ;
        RECT 2111.010 1686.160 2115.455 1686.300 ;
        RECT 2111.010 1686.100 2111.330 1686.160 ;
        RECT 2115.165 1686.115 2115.455 1686.160 ;
        RECT 2107.790 20.640 2108.110 20.700 ;
        RECT 2111.010 20.640 2111.330 20.700 ;
        RECT 2107.790 20.500 2111.330 20.640 ;
        RECT 2107.790 20.440 2108.110 20.500 ;
        RECT 2111.010 20.440 2111.330 20.500 ;
      LAYER via ;
        RECT 2232.020 1687.120 2232.280 1687.380 ;
        RECT 2111.040 1686.100 2111.300 1686.360 ;
        RECT 2107.820 20.440 2108.080 20.700 ;
        RECT 2111.040 20.440 2111.300 20.700 ;
      LAYER met2 ;
        RECT 2233.320 1700.410 2233.600 1704.000 ;
        RECT 2232.080 1700.270 2233.600 1700.410 ;
        RECT 2232.080 1687.410 2232.220 1700.270 ;
        RECT 2233.320 1700.000 2233.600 1700.270 ;
        RECT 2232.020 1687.090 2232.280 1687.410 ;
        RECT 2111.040 1686.070 2111.300 1686.390 ;
        RECT 2111.100 20.730 2111.240 1686.070 ;
        RECT 2107.820 20.410 2108.080 20.730 ;
        RECT 2111.040 20.410 2111.300 20.730 ;
        RECT 2107.880 2.400 2108.020 20.410 ;
        RECT 2107.670 -4.800 2108.230 2.400 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2163.525 16.405 2163.695 19.975 ;
      LAYER mcon ;
        RECT 2163.525 19.805 2163.695 19.975 ;
      LAYER met1 ;
        RECT 2163.465 19.960 2163.755 20.005 ;
        RECT 2242.570 19.960 2242.890 20.020 ;
        RECT 2163.465 19.820 2242.890 19.960 ;
        RECT 2163.465 19.775 2163.755 19.820 ;
        RECT 2242.570 19.760 2242.890 19.820 ;
        RECT 2125.730 16.900 2126.050 16.960 ;
        RECT 2125.730 16.760 2161.380 16.900 ;
        RECT 2125.730 16.700 2126.050 16.760 ;
        RECT 2161.240 16.560 2161.380 16.760 ;
        RECT 2163.465 16.560 2163.755 16.605 ;
        RECT 2161.240 16.420 2163.755 16.560 ;
        RECT 2163.465 16.375 2163.755 16.420 ;
      LAYER via ;
        RECT 2242.600 19.760 2242.860 20.020 ;
        RECT 2125.760 16.700 2126.020 16.960 ;
      LAYER met2 ;
        RECT 2242.520 1700.000 2242.800 1704.000 ;
        RECT 2242.660 20.050 2242.800 1700.000 ;
        RECT 2242.600 19.730 2242.860 20.050 ;
        RECT 2125.760 16.670 2126.020 16.990 ;
        RECT 2125.820 2.400 2125.960 16.670 ;
        RECT 2125.610 -4.800 2126.170 2.400 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2167.205 1684.105 2167.375 1686.655 ;
      LAYER mcon ;
        RECT 2167.205 1686.485 2167.375 1686.655 ;
      LAYER met1 ;
        RECT 2167.145 1686.640 2167.435 1686.685 ;
        RECT 2251.770 1686.640 2252.090 1686.700 ;
        RECT 2167.145 1686.500 2252.090 1686.640 ;
        RECT 2167.145 1686.455 2167.435 1686.500 ;
        RECT 2251.770 1686.440 2252.090 1686.500 ;
        RECT 2145.510 1684.260 2145.830 1684.320 ;
        RECT 2167.145 1684.260 2167.435 1684.305 ;
        RECT 2145.510 1684.120 2167.435 1684.260 ;
        RECT 2145.510 1684.060 2145.830 1684.120 ;
        RECT 2167.145 1684.075 2167.435 1684.120 ;
      LAYER via ;
        RECT 2251.800 1686.440 2252.060 1686.700 ;
        RECT 2145.540 1684.060 2145.800 1684.320 ;
      LAYER met2 ;
        RECT 2251.720 1700.000 2252.000 1704.000 ;
        RECT 2251.860 1686.730 2252.000 1700.000 ;
        RECT 2251.800 1686.410 2252.060 1686.730 ;
        RECT 2145.540 1684.030 2145.800 1684.350 ;
        RECT 2145.600 3.130 2145.740 1684.030 ;
        RECT 2143.760 2.990 2145.740 3.130 ;
        RECT 2143.760 2.400 2143.900 2.990 ;
        RECT 2143.550 -4.800 2144.110 2.400 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2257.825 1510.365 2257.995 1579.895 ;
        RECT 2257.825 1317.245 2257.995 1368.755 ;
        RECT 2257.825 1220.685 2257.995 1297.015 ;
        RECT 2256.445 1110.865 2256.615 1124.975 ;
        RECT 2257.825 737.885 2257.995 814.215 ;
        RECT 2238.045 16.065 2238.215 16.915 ;
      LAYER mcon ;
        RECT 2257.825 1579.725 2257.995 1579.895 ;
        RECT 2257.825 1368.585 2257.995 1368.755 ;
        RECT 2257.825 1296.845 2257.995 1297.015 ;
        RECT 2256.445 1124.805 2256.615 1124.975 ;
        RECT 2257.825 814.045 2257.995 814.215 ;
        RECT 2238.045 16.745 2238.215 16.915 ;
      LAYER met1 ;
        RECT 2256.830 1628.500 2257.150 1628.560 ;
        RECT 2257.750 1628.500 2258.070 1628.560 ;
        RECT 2256.830 1628.360 2258.070 1628.500 ;
        RECT 2256.830 1628.300 2257.150 1628.360 ;
        RECT 2257.750 1628.300 2258.070 1628.360 ;
        RECT 2257.750 1580.560 2258.070 1580.620 ;
        RECT 2258.670 1580.560 2258.990 1580.620 ;
        RECT 2257.750 1580.420 2258.990 1580.560 ;
        RECT 2257.750 1580.360 2258.070 1580.420 ;
        RECT 2258.670 1580.360 2258.990 1580.420 ;
        RECT 2257.750 1579.880 2258.070 1579.940 ;
        RECT 2257.555 1579.740 2258.070 1579.880 ;
        RECT 2257.750 1579.680 2258.070 1579.740 ;
        RECT 2257.750 1510.520 2258.070 1510.580 ;
        RECT 2257.555 1510.380 2258.070 1510.520 ;
        RECT 2257.750 1510.320 2258.070 1510.380 ;
        RECT 2257.750 1463.260 2258.070 1463.320 ;
        RECT 2257.380 1463.120 2258.070 1463.260 ;
        RECT 2257.380 1462.640 2257.520 1463.120 ;
        RECT 2257.750 1463.060 2258.070 1463.120 ;
        RECT 2257.290 1462.380 2257.610 1462.640 ;
        RECT 2256.370 1393.900 2256.690 1393.960 ;
        RECT 2257.750 1393.900 2258.070 1393.960 ;
        RECT 2256.370 1393.760 2258.070 1393.900 ;
        RECT 2256.370 1393.700 2256.690 1393.760 ;
        RECT 2257.750 1393.700 2258.070 1393.760 ;
        RECT 2257.750 1368.740 2258.070 1368.800 ;
        RECT 2257.555 1368.600 2258.070 1368.740 ;
        RECT 2257.750 1368.540 2258.070 1368.600 ;
        RECT 2257.750 1317.400 2258.070 1317.460 ;
        RECT 2257.555 1317.260 2258.070 1317.400 ;
        RECT 2257.750 1317.200 2258.070 1317.260 ;
        RECT 2257.750 1297.000 2258.070 1297.060 ;
        RECT 2257.555 1296.860 2258.070 1297.000 ;
        RECT 2257.750 1296.800 2258.070 1296.860 ;
        RECT 2257.750 1220.840 2258.070 1220.900 ;
        RECT 2257.555 1220.700 2258.070 1220.840 ;
        RECT 2257.750 1220.640 2258.070 1220.700 ;
        RECT 2257.750 1173.580 2258.070 1173.640 ;
        RECT 2257.380 1173.440 2258.070 1173.580 ;
        RECT 2257.380 1172.960 2257.520 1173.440 ;
        RECT 2257.750 1173.380 2258.070 1173.440 ;
        RECT 2257.290 1172.700 2257.610 1172.960 ;
        RECT 2256.385 1124.960 2256.675 1125.005 ;
        RECT 2256.830 1124.960 2257.150 1125.020 ;
        RECT 2256.385 1124.820 2257.150 1124.960 ;
        RECT 2256.385 1124.775 2256.675 1124.820 ;
        RECT 2256.830 1124.760 2257.150 1124.820 ;
        RECT 2256.370 1111.020 2256.690 1111.080 ;
        RECT 2256.175 1110.880 2256.690 1111.020 ;
        RECT 2256.370 1110.820 2256.690 1110.880 ;
        RECT 2258.210 932.320 2258.530 932.580 ;
        RECT 2258.300 931.900 2258.440 932.320 ;
        RECT 2258.210 931.640 2258.530 931.900 ;
        RECT 2258.670 862.480 2258.990 862.540 ;
        RECT 2260.050 862.480 2260.370 862.540 ;
        RECT 2258.670 862.340 2260.370 862.480 ;
        RECT 2258.670 862.280 2258.990 862.340 ;
        RECT 2260.050 862.280 2260.370 862.340 ;
        RECT 2257.765 814.200 2258.055 814.245 ;
        RECT 2258.670 814.200 2258.990 814.260 ;
        RECT 2257.765 814.060 2258.990 814.200 ;
        RECT 2257.765 814.015 2258.055 814.060 ;
        RECT 2258.670 814.000 2258.990 814.060 ;
        RECT 2257.750 738.040 2258.070 738.100 ;
        RECT 2257.555 737.900 2258.070 738.040 ;
        RECT 2257.750 737.840 2258.070 737.900 ;
        RECT 2257.750 689.900 2258.070 690.160 ;
        RECT 2257.840 689.760 2257.980 689.900 ;
        RECT 2258.670 689.760 2258.990 689.820 ;
        RECT 2257.840 689.620 2258.990 689.760 ;
        RECT 2258.670 689.560 2258.990 689.620 ;
        RECT 2257.750 641.820 2258.070 641.880 ;
        RECT 2258.670 641.820 2258.990 641.880 ;
        RECT 2257.750 641.680 2258.990 641.820 ;
        RECT 2257.750 641.620 2258.070 641.680 ;
        RECT 2258.670 641.620 2258.990 641.680 ;
        RECT 2258.670 593.680 2258.990 593.940 ;
        RECT 2258.760 593.260 2258.900 593.680 ;
        RECT 2258.670 593.000 2258.990 593.260 ;
        RECT 2256.830 234.840 2257.150 234.900 ;
        RECT 2258.210 234.840 2258.530 234.900 ;
        RECT 2256.830 234.700 2258.530 234.840 ;
        RECT 2256.830 234.640 2257.150 234.700 ;
        RECT 2258.210 234.640 2258.530 234.700 ;
        RECT 2256.830 206.620 2257.150 206.680 ;
        RECT 2258.670 206.620 2258.990 206.680 ;
        RECT 2256.830 206.480 2258.990 206.620 ;
        RECT 2256.830 206.420 2257.150 206.480 ;
        RECT 2258.670 206.420 2258.990 206.480 ;
        RECT 2258.670 159.020 2258.990 159.080 ;
        RECT 2258.300 158.880 2258.990 159.020 ;
        RECT 2258.300 158.740 2258.440 158.880 ;
        RECT 2258.670 158.820 2258.990 158.880 ;
        RECT 2258.210 158.480 2258.530 158.740 ;
        RECT 2161.610 16.900 2161.930 16.960 ;
        RECT 2237.985 16.900 2238.275 16.945 ;
        RECT 2161.610 16.760 2238.275 16.900 ;
        RECT 2161.610 16.700 2161.930 16.760 ;
        RECT 2237.985 16.715 2238.275 16.760 ;
        RECT 2237.985 16.220 2238.275 16.265 ;
        RECT 2257.750 16.220 2258.070 16.280 ;
        RECT 2237.985 16.080 2258.070 16.220 ;
        RECT 2237.985 16.035 2238.275 16.080 ;
        RECT 2257.750 16.020 2258.070 16.080 ;
      LAYER via ;
        RECT 2256.860 1628.300 2257.120 1628.560 ;
        RECT 2257.780 1628.300 2258.040 1628.560 ;
        RECT 2257.780 1580.360 2258.040 1580.620 ;
        RECT 2258.700 1580.360 2258.960 1580.620 ;
        RECT 2257.780 1579.680 2258.040 1579.940 ;
        RECT 2257.780 1510.320 2258.040 1510.580 ;
        RECT 2257.780 1463.060 2258.040 1463.320 ;
        RECT 2257.320 1462.380 2257.580 1462.640 ;
        RECT 2256.400 1393.700 2256.660 1393.960 ;
        RECT 2257.780 1393.700 2258.040 1393.960 ;
        RECT 2257.780 1368.540 2258.040 1368.800 ;
        RECT 2257.780 1317.200 2258.040 1317.460 ;
        RECT 2257.780 1296.800 2258.040 1297.060 ;
        RECT 2257.780 1220.640 2258.040 1220.900 ;
        RECT 2257.780 1173.380 2258.040 1173.640 ;
        RECT 2257.320 1172.700 2257.580 1172.960 ;
        RECT 2256.860 1124.760 2257.120 1125.020 ;
        RECT 2256.400 1110.820 2256.660 1111.080 ;
        RECT 2258.240 932.320 2258.500 932.580 ;
        RECT 2258.240 931.640 2258.500 931.900 ;
        RECT 2258.700 862.280 2258.960 862.540 ;
        RECT 2260.080 862.280 2260.340 862.540 ;
        RECT 2258.700 814.000 2258.960 814.260 ;
        RECT 2257.780 737.840 2258.040 738.100 ;
        RECT 2257.780 689.900 2258.040 690.160 ;
        RECT 2258.700 689.560 2258.960 689.820 ;
        RECT 2257.780 641.620 2258.040 641.880 ;
        RECT 2258.700 641.620 2258.960 641.880 ;
        RECT 2258.700 593.680 2258.960 593.940 ;
        RECT 2258.700 593.000 2258.960 593.260 ;
        RECT 2256.860 234.640 2257.120 234.900 ;
        RECT 2258.240 234.640 2258.500 234.900 ;
        RECT 2256.860 206.420 2257.120 206.680 ;
        RECT 2258.700 206.420 2258.960 206.680 ;
        RECT 2258.700 158.820 2258.960 159.080 ;
        RECT 2258.240 158.480 2258.500 158.740 ;
        RECT 2161.640 16.700 2161.900 16.960 ;
        RECT 2257.780 16.020 2258.040 16.280 ;
      LAYER met2 ;
        RECT 2260.920 1700.410 2261.200 1704.000 ;
        RECT 2259.220 1700.270 2261.200 1700.410 ;
        RECT 2259.220 1676.725 2259.360 1700.270 ;
        RECT 2260.920 1700.000 2261.200 1700.270 ;
        RECT 2256.850 1676.355 2257.130 1676.725 ;
        RECT 2259.150 1676.355 2259.430 1676.725 ;
        RECT 2256.920 1628.590 2257.060 1676.355 ;
        RECT 2256.860 1628.270 2257.120 1628.590 ;
        RECT 2257.780 1628.445 2258.040 1628.590 ;
        RECT 2257.770 1628.075 2258.050 1628.445 ;
        RECT 2258.690 1628.075 2258.970 1628.445 ;
        RECT 2258.760 1580.650 2258.900 1628.075 ;
        RECT 2257.780 1580.330 2258.040 1580.650 ;
        RECT 2258.700 1580.330 2258.960 1580.650 ;
        RECT 2257.840 1579.970 2257.980 1580.330 ;
        RECT 2257.780 1579.650 2258.040 1579.970 ;
        RECT 2257.780 1510.290 2258.040 1510.610 ;
        RECT 2257.840 1463.350 2257.980 1510.290 ;
        RECT 2257.780 1463.030 2258.040 1463.350 ;
        RECT 2257.320 1462.350 2257.580 1462.670 ;
        RECT 2257.380 1442.125 2257.520 1462.350 ;
        RECT 2256.390 1441.755 2256.670 1442.125 ;
        RECT 2257.310 1441.755 2257.590 1442.125 ;
        RECT 2256.460 1393.990 2256.600 1441.755 ;
        RECT 2256.400 1393.670 2256.660 1393.990 ;
        RECT 2257.780 1393.670 2258.040 1393.990 ;
        RECT 2257.840 1368.830 2257.980 1393.670 ;
        RECT 2257.780 1368.510 2258.040 1368.830 ;
        RECT 2257.780 1317.170 2258.040 1317.490 ;
        RECT 2257.840 1297.090 2257.980 1317.170 ;
        RECT 2257.780 1296.770 2258.040 1297.090 ;
        RECT 2257.780 1220.610 2258.040 1220.930 ;
        RECT 2257.840 1173.670 2257.980 1220.610 ;
        RECT 2257.780 1173.350 2258.040 1173.670 ;
        RECT 2257.320 1172.670 2257.580 1172.990 ;
        RECT 2257.380 1159.130 2257.520 1172.670 ;
        RECT 2256.920 1158.990 2257.520 1159.130 ;
        RECT 2256.920 1125.050 2257.060 1158.990 ;
        RECT 2256.860 1124.730 2257.120 1125.050 ;
        RECT 2256.400 1110.965 2256.660 1111.110 ;
        RECT 2256.390 1110.595 2256.670 1110.965 ;
        RECT 2258.690 1109.915 2258.970 1110.285 ;
        RECT 2258.760 1027.890 2258.900 1109.915 ;
        RECT 2258.300 1027.750 2258.900 1027.890 ;
        RECT 2258.300 980.290 2258.440 1027.750 ;
        RECT 2257.840 980.150 2258.440 980.290 ;
        RECT 2257.840 979.610 2257.980 980.150 ;
        RECT 2257.840 979.470 2258.440 979.610 ;
        RECT 2258.300 932.610 2258.440 979.470 ;
        RECT 2258.240 932.290 2258.500 932.610 ;
        RECT 2258.240 931.610 2258.500 931.930 ;
        RECT 2258.300 910.930 2258.440 931.610 ;
        RECT 2258.300 910.790 2258.900 910.930 ;
        RECT 2258.760 862.570 2258.900 910.790 ;
        RECT 2258.700 862.250 2258.960 862.570 ;
        RECT 2260.080 862.250 2260.340 862.570 ;
        RECT 2260.140 814.485 2260.280 862.250 ;
        RECT 2259.150 814.370 2259.430 814.485 ;
        RECT 2258.760 814.290 2259.430 814.370 ;
        RECT 2258.700 814.230 2259.430 814.290 ;
        RECT 2258.700 813.970 2258.960 814.230 ;
        RECT 2259.150 814.115 2259.430 814.230 ;
        RECT 2260.070 814.115 2260.350 814.485 ;
        RECT 2257.780 737.810 2258.040 738.130 ;
        RECT 2257.840 690.190 2257.980 737.810 ;
        RECT 2257.780 689.870 2258.040 690.190 ;
        RECT 2258.700 689.530 2258.960 689.850 ;
        RECT 2258.760 641.910 2258.900 689.530 ;
        RECT 2257.780 641.650 2258.040 641.910 ;
        RECT 2258.700 641.650 2258.960 641.910 ;
        RECT 2257.780 641.590 2258.960 641.650 ;
        RECT 2257.840 641.510 2258.900 641.590 ;
        RECT 2258.760 593.970 2258.900 641.510 ;
        RECT 2258.700 593.650 2258.960 593.970 ;
        RECT 2258.700 592.970 2258.960 593.290 ;
        RECT 2258.760 579.770 2258.900 592.970 ;
        RECT 2258.760 579.630 2259.360 579.770 ;
        RECT 2259.220 545.090 2259.360 579.630 ;
        RECT 2258.300 544.950 2259.360 545.090 ;
        RECT 2258.300 497.605 2258.440 544.950 ;
        RECT 2258.230 497.235 2258.510 497.605 ;
        RECT 2258.230 482.955 2258.510 483.325 ;
        RECT 2258.300 234.930 2258.440 482.955 ;
        RECT 2256.860 234.610 2257.120 234.930 ;
        RECT 2258.240 234.610 2258.500 234.930 ;
        RECT 2256.920 206.710 2257.060 234.610 ;
        RECT 2256.860 206.390 2257.120 206.710 ;
        RECT 2258.700 206.390 2258.960 206.710 ;
        RECT 2258.760 159.110 2258.900 206.390 ;
        RECT 2258.700 158.790 2258.960 159.110 ;
        RECT 2258.240 158.450 2258.500 158.770 ;
        RECT 2258.300 110.570 2258.440 158.450 ;
        RECT 2258.300 110.430 2258.900 110.570 ;
        RECT 2258.760 62.290 2258.900 110.430 ;
        RECT 2257.840 62.150 2258.900 62.290 ;
        RECT 2161.640 16.670 2161.900 16.990 ;
        RECT 2161.700 2.400 2161.840 16.670 ;
        RECT 2257.840 16.310 2257.980 62.150 ;
        RECT 2257.780 15.990 2258.040 16.310 ;
        RECT 2161.490 -4.800 2162.050 2.400 ;
      LAYER via2 ;
        RECT 2256.850 1676.400 2257.130 1676.680 ;
        RECT 2259.150 1676.400 2259.430 1676.680 ;
        RECT 2257.770 1628.120 2258.050 1628.400 ;
        RECT 2258.690 1628.120 2258.970 1628.400 ;
        RECT 2256.390 1441.800 2256.670 1442.080 ;
        RECT 2257.310 1441.800 2257.590 1442.080 ;
        RECT 2256.390 1110.640 2256.670 1110.920 ;
        RECT 2258.690 1109.960 2258.970 1110.240 ;
        RECT 2259.150 814.160 2259.430 814.440 ;
        RECT 2260.070 814.160 2260.350 814.440 ;
        RECT 2258.230 497.280 2258.510 497.560 ;
        RECT 2258.230 483.000 2258.510 483.280 ;
      LAYER met3 ;
        RECT 2256.825 1676.690 2257.155 1676.705 ;
        RECT 2259.125 1676.690 2259.455 1676.705 ;
        RECT 2256.825 1676.390 2259.455 1676.690 ;
        RECT 2256.825 1676.375 2257.155 1676.390 ;
        RECT 2259.125 1676.375 2259.455 1676.390 ;
        RECT 2257.745 1628.410 2258.075 1628.425 ;
        RECT 2258.665 1628.410 2258.995 1628.425 ;
        RECT 2257.745 1628.110 2258.995 1628.410 ;
        RECT 2257.745 1628.095 2258.075 1628.110 ;
        RECT 2258.665 1628.095 2258.995 1628.110 ;
        RECT 2256.365 1442.090 2256.695 1442.105 ;
        RECT 2257.285 1442.090 2257.615 1442.105 ;
        RECT 2256.365 1441.790 2257.615 1442.090 ;
        RECT 2256.365 1441.775 2256.695 1441.790 ;
        RECT 2257.285 1441.775 2257.615 1441.790 ;
        RECT 2256.365 1110.930 2256.695 1110.945 ;
        RECT 2256.150 1110.615 2256.695 1110.930 ;
        RECT 2256.150 1110.250 2256.450 1110.615 ;
        RECT 2258.665 1110.250 2258.995 1110.265 ;
        RECT 2256.150 1109.950 2258.995 1110.250 ;
        RECT 2258.665 1109.935 2258.995 1109.950 ;
        RECT 2259.125 814.450 2259.455 814.465 ;
        RECT 2260.045 814.450 2260.375 814.465 ;
        RECT 2259.125 814.150 2260.375 814.450 ;
        RECT 2259.125 814.135 2259.455 814.150 ;
        RECT 2260.045 814.135 2260.375 814.150 ;
        RECT 2258.205 497.580 2258.535 497.585 ;
        RECT 2257.950 497.570 2258.535 497.580 ;
        RECT 2257.750 497.270 2258.535 497.570 ;
        RECT 2257.950 497.260 2258.535 497.270 ;
        RECT 2258.205 497.255 2258.535 497.260 ;
        RECT 2258.205 483.300 2258.535 483.305 ;
        RECT 2257.950 483.290 2258.535 483.300 ;
        RECT 2257.950 482.990 2258.760 483.290 ;
        RECT 2257.950 482.980 2258.535 482.990 ;
        RECT 2258.205 482.975 2258.535 482.980 ;
      LAYER via3 ;
        RECT 2257.980 497.260 2258.300 497.580 ;
        RECT 2257.980 482.980 2258.300 483.300 ;
      LAYER met4 ;
        RECT 2257.975 497.255 2258.305 497.585 ;
        RECT 2257.990 483.305 2258.290 497.255 ;
        RECT 2257.975 482.975 2258.305 483.305 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2180.010 1685.280 2180.330 1685.340 ;
        RECT 2270.170 1685.280 2270.490 1685.340 ;
        RECT 2180.010 1685.140 2270.490 1685.280 ;
        RECT 2180.010 1685.080 2180.330 1685.140 ;
        RECT 2270.170 1685.080 2270.490 1685.140 ;
        RECT 2179.090 2.960 2179.410 3.020 ;
        RECT 2180.010 2.960 2180.330 3.020 ;
        RECT 2179.090 2.820 2180.330 2.960 ;
        RECT 2179.090 2.760 2179.410 2.820 ;
        RECT 2180.010 2.760 2180.330 2.820 ;
      LAYER via ;
        RECT 2180.040 1685.080 2180.300 1685.340 ;
        RECT 2270.200 1685.080 2270.460 1685.340 ;
        RECT 2179.120 2.760 2179.380 3.020 ;
        RECT 2180.040 2.760 2180.300 3.020 ;
      LAYER met2 ;
        RECT 2270.120 1700.000 2270.400 1704.000 ;
        RECT 2270.260 1685.370 2270.400 1700.000 ;
        RECT 2180.040 1685.050 2180.300 1685.370 ;
        RECT 2270.200 1685.050 2270.460 1685.370 ;
        RECT 2180.100 3.050 2180.240 1685.050 ;
        RECT 2179.120 2.730 2179.380 3.050 ;
        RECT 2180.040 2.730 2180.300 3.050 ;
        RECT 2179.180 2.400 2179.320 2.730 ;
        RECT 2178.970 -4.800 2179.530 2.400 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2197.030 17.920 2197.350 17.980 ;
        RECT 2277.990 17.920 2278.310 17.980 ;
        RECT 2197.030 17.780 2278.310 17.920 ;
        RECT 2197.030 17.720 2197.350 17.780 ;
        RECT 2277.990 17.720 2278.310 17.780 ;
      LAYER via ;
        RECT 2197.060 17.720 2197.320 17.980 ;
        RECT 2278.020 17.720 2278.280 17.980 ;
      LAYER met2 ;
        RECT 2279.320 1700.410 2279.600 1704.000 ;
        RECT 2278.080 1700.270 2279.600 1700.410 ;
        RECT 2278.080 18.010 2278.220 1700.270 ;
        RECT 2279.320 1700.000 2279.600 1700.270 ;
        RECT 2197.060 17.690 2197.320 18.010 ;
        RECT 2278.020 17.690 2278.280 18.010 ;
        RECT 2197.120 2.400 2197.260 17.690 ;
        RECT 2196.910 -4.800 2197.470 2.400 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2214.970 18.260 2215.290 18.320 ;
        RECT 2284.890 18.260 2285.210 18.320 ;
        RECT 2214.970 18.120 2285.210 18.260 ;
        RECT 2214.970 18.060 2215.290 18.120 ;
        RECT 2284.890 18.060 2285.210 18.120 ;
      LAYER via ;
        RECT 2215.000 18.060 2215.260 18.320 ;
        RECT 2284.920 18.060 2285.180 18.320 ;
      LAYER met2 ;
        RECT 2288.520 1701.090 2288.800 1704.000 ;
        RECT 2286.360 1700.950 2288.800 1701.090 ;
        RECT 2286.360 1656.210 2286.500 1700.950 ;
        RECT 2288.520 1700.000 2288.800 1700.950 ;
        RECT 2284.980 1656.070 2286.500 1656.210 ;
        RECT 2284.980 18.350 2285.120 1656.070 ;
        RECT 2215.000 18.030 2215.260 18.350 ;
        RECT 2284.920 18.030 2285.180 18.350 ;
        RECT 2215.060 2.400 2215.200 18.030 ;
        RECT 2214.850 -4.800 2215.410 2.400 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2232.910 17.240 2233.230 17.300 ;
        RECT 2298.690 17.240 2299.010 17.300 ;
        RECT 2232.910 17.100 2299.010 17.240 ;
        RECT 2232.910 17.040 2233.230 17.100 ;
        RECT 2298.690 17.040 2299.010 17.100 ;
      LAYER via ;
        RECT 2232.940 17.040 2233.200 17.300 ;
        RECT 2298.720 17.040 2298.980 17.300 ;
      LAYER met2 ;
        RECT 2297.720 1700.410 2298.000 1704.000 ;
        RECT 2297.720 1700.270 2298.920 1700.410 ;
        RECT 2297.720 1700.000 2298.000 1700.270 ;
        RECT 2298.780 17.330 2298.920 1700.270 ;
        RECT 2232.940 17.010 2233.200 17.330 ;
        RECT 2298.720 17.010 2298.980 17.330 ;
        RECT 2233.000 2.400 2233.140 17.010 ;
        RECT 2232.790 -4.800 2233.350 2.400 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 793.110 50.220 793.430 50.280 ;
        RECT 1552.570 50.220 1552.890 50.280 ;
        RECT 793.110 50.080 1552.890 50.220 ;
        RECT 793.110 50.020 793.430 50.080 ;
        RECT 1552.570 50.020 1552.890 50.080 ;
      LAYER via ;
        RECT 793.140 50.020 793.400 50.280 ;
        RECT 1552.600 50.020 1552.860 50.280 ;
      LAYER met2 ;
        RECT 1553.900 1700.410 1554.180 1704.000 ;
        RECT 1552.660 1700.270 1554.180 1700.410 ;
        RECT 1552.660 50.310 1552.800 1700.270 ;
        RECT 1553.900 1700.000 1554.180 1700.270 ;
        RECT 793.140 49.990 793.400 50.310 ;
        RECT 1552.600 49.990 1552.860 50.310 ;
        RECT 793.200 16.730 793.340 49.990 ;
        RECT 787.680 16.590 793.340 16.730 ;
        RECT 787.680 2.400 787.820 16.590 ;
        RECT 787.470 -4.800 788.030 2.400 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2255.910 1687.660 2256.230 1687.720 ;
        RECT 2306.970 1687.660 2307.290 1687.720 ;
        RECT 2255.910 1687.520 2307.290 1687.660 ;
        RECT 2255.910 1687.460 2256.230 1687.520 ;
        RECT 2306.970 1687.460 2307.290 1687.520 ;
        RECT 2250.850 18.600 2251.170 18.660 ;
        RECT 2255.910 18.600 2256.230 18.660 ;
        RECT 2250.850 18.460 2256.230 18.600 ;
        RECT 2250.850 18.400 2251.170 18.460 ;
        RECT 2255.910 18.400 2256.230 18.460 ;
      LAYER via ;
        RECT 2255.940 1687.460 2256.200 1687.720 ;
        RECT 2307.000 1687.460 2307.260 1687.720 ;
        RECT 2250.880 18.400 2251.140 18.660 ;
        RECT 2255.940 18.400 2256.200 18.660 ;
      LAYER met2 ;
        RECT 2306.920 1700.000 2307.200 1704.000 ;
        RECT 2307.060 1687.750 2307.200 1700.000 ;
        RECT 2255.940 1687.430 2256.200 1687.750 ;
        RECT 2307.000 1687.430 2307.260 1687.750 ;
        RECT 2256.000 18.690 2256.140 1687.430 ;
        RECT 2250.880 18.370 2251.140 18.690 ;
        RECT 2255.940 18.370 2256.200 18.690 ;
        RECT 2250.940 2.400 2251.080 18.370 ;
        RECT 2250.730 -4.800 2251.290 2.400 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2269.710 1688.000 2270.030 1688.060 ;
        RECT 2316.170 1688.000 2316.490 1688.060 ;
        RECT 2269.710 1687.860 2316.490 1688.000 ;
        RECT 2269.710 1687.800 2270.030 1687.860 ;
        RECT 2316.170 1687.800 2316.490 1687.860 ;
        RECT 2268.330 2.960 2268.650 3.020 ;
        RECT 2269.710 2.960 2270.030 3.020 ;
        RECT 2268.330 2.820 2270.030 2.960 ;
        RECT 2268.330 2.760 2268.650 2.820 ;
        RECT 2269.710 2.760 2270.030 2.820 ;
      LAYER via ;
        RECT 2269.740 1687.800 2270.000 1688.060 ;
        RECT 2316.200 1687.800 2316.460 1688.060 ;
        RECT 2268.360 2.760 2268.620 3.020 ;
        RECT 2269.740 2.760 2270.000 3.020 ;
      LAYER met2 ;
        RECT 2316.120 1700.000 2316.400 1704.000 ;
        RECT 2316.260 1688.090 2316.400 1700.000 ;
        RECT 2269.740 1687.770 2270.000 1688.090 ;
        RECT 2316.200 1687.770 2316.460 1688.090 ;
        RECT 2269.800 3.050 2269.940 1687.770 ;
        RECT 2268.360 2.730 2268.620 3.050 ;
        RECT 2269.740 2.730 2270.000 3.050 ;
        RECT 2268.420 2.400 2268.560 2.730 ;
        RECT 2268.210 -4.800 2268.770 2.400 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2286.270 17.920 2286.590 17.980 ;
        RECT 2325.370 17.920 2325.690 17.980 ;
        RECT 2286.270 17.780 2325.690 17.920 ;
        RECT 2286.270 17.720 2286.590 17.780 ;
        RECT 2325.370 17.720 2325.690 17.780 ;
      LAYER via ;
        RECT 2286.300 17.720 2286.560 17.980 ;
        RECT 2325.400 17.720 2325.660 17.980 ;
      LAYER met2 ;
        RECT 2325.320 1700.000 2325.600 1704.000 ;
        RECT 2325.460 18.010 2325.600 1700.000 ;
        RECT 2286.300 17.690 2286.560 18.010 ;
        RECT 2325.400 17.690 2325.660 18.010 ;
        RECT 2286.360 2.400 2286.500 17.690 ;
        RECT 2286.150 -4.800 2286.710 2.400 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2304.210 1686.980 2304.530 1687.040 ;
        RECT 2334.570 1686.980 2334.890 1687.040 ;
        RECT 2304.210 1686.840 2334.890 1686.980 ;
        RECT 2304.210 1686.780 2304.530 1686.840 ;
        RECT 2334.570 1686.780 2334.890 1686.840 ;
      LAYER via ;
        RECT 2304.240 1686.780 2304.500 1687.040 ;
        RECT 2334.600 1686.780 2334.860 1687.040 ;
      LAYER met2 ;
        RECT 2334.520 1700.000 2334.800 1704.000 ;
        RECT 2334.660 1687.070 2334.800 1700.000 ;
        RECT 2304.240 1686.750 2304.500 1687.070 ;
        RECT 2334.600 1686.750 2334.860 1687.070 ;
        RECT 2304.300 2.400 2304.440 1686.750 ;
        RECT 2304.090 -4.800 2304.650 2.400 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2343.770 1684.600 2344.090 1684.660 ;
        RECT 2337.880 1684.460 2344.090 1684.600 ;
        RECT 2324.910 1684.260 2325.230 1684.320 ;
        RECT 2337.880 1684.260 2338.020 1684.460 ;
        RECT 2343.770 1684.400 2344.090 1684.460 ;
        RECT 2324.910 1684.120 2338.020 1684.260 ;
        RECT 2324.910 1684.060 2325.230 1684.120 ;
        RECT 2322.150 16.560 2322.470 16.620 ;
        RECT 2324.910 16.560 2325.230 16.620 ;
        RECT 2322.150 16.420 2325.230 16.560 ;
        RECT 2322.150 16.360 2322.470 16.420 ;
        RECT 2324.910 16.360 2325.230 16.420 ;
      LAYER via ;
        RECT 2324.940 1684.060 2325.200 1684.320 ;
        RECT 2343.800 1684.400 2344.060 1684.660 ;
        RECT 2322.180 16.360 2322.440 16.620 ;
        RECT 2324.940 16.360 2325.200 16.620 ;
      LAYER met2 ;
        RECT 2343.720 1700.000 2344.000 1704.000 ;
        RECT 2343.860 1684.690 2344.000 1700.000 ;
        RECT 2343.800 1684.370 2344.060 1684.690 ;
        RECT 2324.940 1684.030 2325.200 1684.350 ;
        RECT 2325.000 16.650 2325.140 1684.030 ;
        RECT 2322.180 16.330 2322.440 16.650 ;
        RECT 2324.940 16.330 2325.200 16.650 ;
        RECT 2322.240 2.400 2322.380 16.330 ;
        RECT 2322.030 -4.800 2322.590 2.400 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2339.630 19.280 2339.950 19.340 ;
        RECT 2353.430 19.280 2353.750 19.340 ;
        RECT 2339.630 19.140 2353.750 19.280 ;
        RECT 2339.630 19.080 2339.950 19.140 ;
        RECT 2353.430 19.080 2353.750 19.140 ;
      LAYER via ;
        RECT 2339.660 19.080 2339.920 19.340 ;
        RECT 2353.460 19.080 2353.720 19.340 ;
      LAYER met2 ;
        RECT 2352.920 1700.410 2353.200 1704.000 ;
        RECT 2352.920 1700.270 2353.660 1700.410 ;
        RECT 2352.920 1700.000 2353.200 1700.270 ;
        RECT 2353.520 19.370 2353.660 1700.270 ;
        RECT 2339.660 19.050 2339.920 19.370 ;
        RECT 2353.460 19.050 2353.720 19.370 ;
        RECT 2339.720 2.400 2339.860 19.050 ;
        RECT 2339.510 -4.800 2340.070 2.400 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2357.570 14.180 2357.890 14.240 ;
        RECT 2359.410 14.180 2359.730 14.240 ;
        RECT 2357.570 14.040 2359.730 14.180 ;
        RECT 2357.570 13.980 2357.890 14.040 ;
        RECT 2359.410 13.980 2359.730 14.040 ;
      LAYER via ;
        RECT 2357.600 13.980 2357.860 14.240 ;
        RECT 2359.440 13.980 2359.700 14.240 ;
      LAYER met2 ;
        RECT 2362.120 1700.410 2362.400 1704.000 ;
        RECT 2359.960 1700.270 2362.400 1700.410 ;
        RECT 2359.960 1683.920 2360.100 1700.270 ;
        RECT 2362.120 1700.000 2362.400 1700.270 ;
        RECT 2359.500 1683.780 2360.100 1683.920 ;
        RECT 2359.500 14.270 2359.640 1683.780 ;
        RECT 2357.600 13.950 2357.860 14.270 ;
        RECT 2359.440 13.950 2359.700 14.270 ;
        RECT 2357.660 2.400 2357.800 13.950 ;
        RECT 2357.450 -4.800 2358.010 2.400 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2373.210 20.640 2373.530 20.700 ;
        RECT 2375.510 20.640 2375.830 20.700 ;
        RECT 2373.210 20.500 2375.830 20.640 ;
        RECT 2373.210 20.440 2373.530 20.500 ;
        RECT 2375.510 20.440 2375.830 20.500 ;
      LAYER via ;
        RECT 2373.240 20.440 2373.500 20.700 ;
        RECT 2375.540 20.440 2375.800 20.700 ;
      LAYER met2 ;
        RECT 2371.320 1700.410 2371.600 1704.000 ;
        RECT 2371.320 1700.270 2373.440 1700.410 ;
        RECT 2371.320 1700.000 2371.600 1700.270 ;
        RECT 2373.300 20.730 2373.440 1700.270 ;
        RECT 2373.240 20.410 2373.500 20.730 ;
        RECT 2375.540 20.410 2375.800 20.730 ;
        RECT 2375.600 2.400 2375.740 20.410 ;
        RECT 2375.390 -4.800 2375.950 2.400 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2380.570 1683.920 2380.890 1683.980 ;
        RECT 2387.930 1683.920 2388.250 1683.980 ;
        RECT 2380.570 1683.780 2388.250 1683.920 ;
        RECT 2380.570 1683.720 2380.890 1683.780 ;
        RECT 2387.930 1683.720 2388.250 1683.780 ;
        RECT 2387.930 37.980 2388.250 38.040 ;
        RECT 2393.450 37.980 2393.770 38.040 ;
        RECT 2387.930 37.840 2393.770 37.980 ;
        RECT 2387.930 37.780 2388.250 37.840 ;
        RECT 2393.450 37.780 2393.770 37.840 ;
      LAYER via ;
        RECT 2380.600 1683.720 2380.860 1683.980 ;
        RECT 2387.960 1683.720 2388.220 1683.980 ;
        RECT 2387.960 37.780 2388.220 38.040 ;
        RECT 2393.480 37.780 2393.740 38.040 ;
      LAYER met2 ;
        RECT 2380.520 1700.000 2380.800 1704.000 ;
        RECT 2380.660 1684.010 2380.800 1700.000 ;
        RECT 2380.600 1683.690 2380.860 1684.010 ;
        RECT 2387.960 1683.690 2388.220 1684.010 ;
        RECT 2388.020 38.070 2388.160 1683.690 ;
        RECT 2387.960 37.750 2388.220 38.070 ;
        RECT 2393.480 37.750 2393.740 38.070 ;
        RECT 2393.540 2.400 2393.680 37.750 ;
        RECT 2393.330 -4.800 2393.890 2.400 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2389.770 1683.920 2390.090 1683.980 ;
        RECT 2393.910 1683.920 2394.230 1683.980 ;
        RECT 2389.770 1683.780 2394.230 1683.920 ;
        RECT 2389.770 1683.720 2390.090 1683.780 ;
        RECT 2393.910 1683.720 2394.230 1683.780 ;
        RECT 2393.910 20.640 2394.230 20.700 ;
        RECT 2411.390 20.640 2411.710 20.700 ;
        RECT 2393.910 20.500 2411.710 20.640 ;
        RECT 2393.910 20.440 2394.230 20.500 ;
        RECT 2411.390 20.440 2411.710 20.500 ;
      LAYER via ;
        RECT 2389.800 1683.720 2390.060 1683.980 ;
        RECT 2393.940 1683.720 2394.200 1683.980 ;
        RECT 2393.940 20.440 2394.200 20.700 ;
        RECT 2411.420 20.440 2411.680 20.700 ;
      LAYER met2 ;
        RECT 2389.720 1700.000 2390.000 1704.000 ;
        RECT 2389.860 1684.010 2390.000 1700.000 ;
        RECT 2389.800 1683.690 2390.060 1684.010 ;
        RECT 2393.940 1683.690 2394.200 1684.010 ;
        RECT 2394.000 20.730 2394.140 1683.690 ;
        RECT 2393.940 20.410 2394.200 20.730 ;
        RECT 2411.420 20.410 2411.680 20.730 ;
        RECT 2411.480 2.400 2411.620 20.410 ;
        RECT 2411.270 -4.800 2411.830 2.400 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1559.470 1689.360 1559.790 1689.420 ;
        RECT 1561.310 1689.360 1561.630 1689.420 ;
        RECT 1559.470 1689.220 1561.630 1689.360 ;
        RECT 1559.470 1689.160 1559.790 1689.220 ;
        RECT 1561.310 1689.160 1561.630 1689.220 ;
        RECT 806.910 49.880 807.230 49.940 ;
        RECT 1559.470 49.880 1559.790 49.940 ;
        RECT 806.910 49.740 1559.790 49.880 ;
        RECT 806.910 49.680 807.230 49.740 ;
        RECT 1559.470 49.680 1559.790 49.740 ;
      LAYER via ;
        RECT 1559.500 1689.160 1559.760 1689.420 ;
        RECT 1561.340 1689.160 1561.600 1689.420 ;
        RECT 806.940 49.680 807.200 49.940 ;
        RECT 1559.500 49.680 1559.760 49.940 ;
      LAYER met2 ;
        RECT 1563.100 1700.410 1563.380 1704.000 ;
        RECT 1561.400 1700.270 1563.380 1700.410 ;
        RECT 1561.400 1689.450 1561.540 1700.270 ;
        RECT 1563.100 1700.000 1563.380 1700.270 ;
        RECT 1559.500 1689.130 1559.760 1689.450 ;
        RECT 1561.340 1689.130 1561.600 1689.450 ;
        RECT 1559.560 49.970 1559.700 1689.130 ;
        RECT 806.940 49.650 807.200 49.970 ;
        RECT 1559.500 49.650 1559.760 49.970 ;
        RECT 807.000 16.730 807.140 49.650 ;
        RECT 805.620 16.590 807.140 16.730 ;
        RECT 805.620 2.400 805.760 16.590 ;
        RECT 805.410 -4.800 805.970 2.400 ;
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2.830 24.040 3.150 24.100 ;
        RECT 1145.470 24.040 1145.790 24.100 ;
        RECT 2.830 23.900 1145.790 24.040 ;
        RECT 2.830 23.840 3.150 23.900 ;
        RECT 1145.470 23.840 1145.790 23.900 ;
      LAYER via ;
        RECT 2.860 23.840 3.120 24.100 ;
        RECT 1145.500 23.840 1145.760 24.100 ;
      LAYER met2 ;
        RECT 1150.020 1700.410 1150.300 1704.000 ;
        RECT 1145.560 1700.270 1150.300 1700.410 ;
        RECT 1145.560 24.130 1145.700 1700.270 ;
        RECT 1150.020 1700.000 1150.300 1700.270 ;
        RECT 2.860 23.810 3.120 24.130 ;
        RECT 1145.500 23.810 1145.760 24.130 ;
        RECT 2.920 2.400 3.060 23.810 ;
        RECT 2.710 -4.800 3.270 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 8.350 24.380 8.670 24.440 ;
        RECT 1152.370 24.380 1152.690 24.440 ;
        RECT 8.350 24.240 1152.690 24.380 ;
        RECT 8.350 24.180 8.670 24.240 ;
        RECT 1152.370 24.180 1152.690 24.240 ;
      LAYER via ;
        RECT 8.380 24.180 8.640 24.440 ;
        RECT 1152.400 24.180 1152.660 24.440 ;
      LAYER met2 ;
        RECT 1152.780 1700.410 1153.060 1704.000 ;
        RECT 1152.460 1700.270 1153.060 1700.410 ;
        RECT 1152.460 24.470 1152.600 1700.270 ;
        RECT 1152.780 1700.000 1153.060 1700.270 ;
        RECT 8.380 24.150 8.640 24.470 ;
        RECT 1152.400 24.150 1152.660 24.470 ;
        RECT 8.440 2.400 8.580 24.150 ;
        RECT 8.230 -4.800 8.790 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 14.330 24.720 14.650 24.780 ;
        RECT 1153.750 24.720 1154.070 24.780 ;
        RECT 14.330 24.580 1154.070 24.720 ;
        RECT 14.330 24.520 14.650 24.580 ;
        RECT 1153.750 24.520 1154.070 24.580 ;
      LAYER via ;
        RECT 14.360 24.520 14.620 24.780 ;
        RECT 1153.780 24.520 1154.040 24.780 ;
      LAYER met2 ;
        RECT 1156.000 1700.410 1156.280 1704.000 ;
        RECT 1153.840 1700.270 1156.280 1700.410 ;
        RECT 1153.840 24.810 1153.980 1700.270 ;
        RECT 1156.000 1700.000 1156.280 1700.270 ;
        RECT 14.360 24.490 14.620 24.810 ;
        RECT 1153.780 24.490 1154.040 24.810 ;
        RECT 14.420 2.400 14.560 24.490 ;
        RECT 14.210 -4.800 14.770 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 38.250 25.060 38.570 25.120 ;
        RECT 1166.170 25.060 1166.490 25.120 ;
        RECT 38.250 24.920 1166.490 25.060 ;
        RECT 38.250 24.860 38.570 24.920 ;
        RECT 1166.170 24.860 1166.490 24.920 ;
      LAYER via ;
        RECT 38.280 24.860 38.540 25.120 ;
        RECT 1166.200 24.860 1166.460 25.120 ;
      LAYER met2 ;
        RECT 1167.960 1700.410 1168.240 1704.000 ;
        RECT 1166.260 1700.270 1168.240 1700.410 ;
        RECT 1166.260 25.150 1166.400 1700.270 ;
        RECT 1167.960 1700.000 1168.240 1700.270 ;
        RECT 38.280 24.830 38.540 25.150 ;
        RECT 1166.200 24.830 1166.460 25.150 ;
        RECT 38.340 2.400 38.480 24.830 ;
        RECT 38.130 -4.800 38.690 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1272.380 1700.410 1272.660 1704.000 ;
        RECT 1269.760 1700.270 1272.660 1700.410 ;
        RECT 1269.760 31.125 1269.900 1700.270 ;
        RECT 1272.380 1700.000 1272.660 1700.270 ;
        RECT 240.670 30.755 240.950 31.125 ;
        RECT 1269.690 30.755 1269.970 31.125 ;
        RECT 240.740 2.400 240.880 30.755 ;
        RECT 240.530 -4.800 241.090 2.400 ;
      LAYER via2 ;
        RECT 240.670 30.800 240.950 31.080 ;
        RECT 1269.690 30.800 1269.970 31.080 ;
      LAYER met3 ;
        RECT 240.645 31.090 240.975 31.105 ;
        RECT 1269.665 31.090 1269.995 31.105 ;
        RECT 240.645 30.790 1269.995 31.090 ;
        RECT 240.645 30.775 240.975 30.790 ;
        RECT 1269.665 30.775 1269.995 30.790 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1277.565 1490.645 1277.735 1579.895 ;
        RECT 1277.565 952.425 1277.735 1000.535 ;
        RECT 1277.565 834.785 1277.735 903.975 ;
        RECT 1277.565 372.725 1277.735 400.095 ;
        RECT 1277.565 276.165 1277.735 324.275 ;
      LAYER mcon ;
        RECT 1277.565 1579.725 1277.735 1579.895 ;
        RECT 1277.565 1000.365 1277.735 1000.535 ;
        RECT 1277.565 903.805 1277.735 903.975 ;
        RECT 1277.565 399.925 1277.735 400.095 ;
        RECT 1277.565 324.105 1277.735 324.275 ;
      LAYER met1 ;
        RECT 1277.030 1586.820 1277.350 1587.080 ;
        RECT 1277.120 1586.680 1277.260 1586.820 ;
        RECT 1278.410 1586.680 1278.730 1586.740 ;
        RECT 1277.120 1586.540 1278.730 1586.680 ;
        RECT 1278.410 1586.480 1278.730 1586.540 ;
        RECT 1277.505 1579.880 1277.795 1579.925 ;
        RECT 1278.410 1579.880 1278.730 1579.940 ;
        RECT 1277.505 1579.740 1278.730 1579.880 ;
        RECT 1277.505 1579.695 1277.795 1579.740 ;
        RECT 1278.410 1579.680 1278.730 1579.740 ;
        RECT 1277.490 1490.800 1277.810 1490.860 ;
        RECT 1277.295 1490.660 1277.810 1490.800 ;
        RECT 1277.490 1490.600 1277.810 1490.660 ;
        RECT 1277.490 1463.060 1277.810 1463.320 ;
        RECT 1277.580 1462.640 1277.720 1463.060 ;
        RECT 1277.490 1462.380 1277.810 1462.640 ;
        RECT 1277.950 1173.240 1278.270 1173.300 ;
        RECT 1277.580 1173.100 1278.270 1173.240 ;
        RECT 1277.580 1172.960 1277.720 1173.100 ;
        RECT 1277.950 1173.040 1278.270 1173.100 ;
        RECT 1277.490 1172.700 1277.810 1172.960 ;
        RECT 1277.950 1076.680 1278.270 1076.740 ;
        RECT 1277.580 1076.540 1278.270 1076.680 ;
        RECT 1277.580 1076.400 1277.720 1076.540 ;
        RECT 1277.950 1076.480 1278.270 1076.540 ;
        RECT 1277.490 1076.140 1277.810 1076.400 ;
        RECT 1276.570 1055.600 1276.890 1055.660 ;
        RECT 1277.490 1055.600 1277.810 1055.660 ;
        RECT 1276.570 1055.460 1277.810 1055.600 ;
        RECT 1276.570 1055.400 1276.890 1055.460 ;
        RECT 1277.490 1055.400 1277.810 1055.460 ;
        RECT 1277.490 1007.320 1277.810 1007.380 ;
        RECT 1277.950 1007.320 1278.270 1007.380 ;
        RECT 1277.490 1007.180 1278.270 1007.320 ;
        RECT 1277.490 1007.120 1277.810 1007.180 ;
        RECT 1277.950 1007.120 1278.270 1007.180 ;
        RECT 1277.490 1000.520 1277.810 1000.580 ;
        RECT 1277.295 1000.380 1277.810 1000.520 ;
        RECT 1277.490 1000.320 1277.810 1000.380 ;
        RECT 1277.490 952.580 1277.810 952.640 ;
        RECT 1277.295 952.440 1277.810 952.580 ;
        RECT 1277.490 952.380 1277.810 952.440 ;
        RECT 1277.490 903.960 1277.810 904.020 ;
        RECT 1277.295 903.820 1277.810 903.960 ;
        RECT 1277.490 903.760 1277.810 903.820 ;
        RECT 1277.490 834.940 1277.810 835.000 ;
        RECT 1277.295 834.800 1277.810 834.940 ;
        RECT 1277.490 834.740 1277.810 834.800 ;
        RECT 1277.490 400.080 1277.810 400.140 ;
        RECT 1277.295 399.940 1277.810 400.080 ;
        RECT 1277.490 399.880 1277.810 399.940 ;
        RECT 1277.490 372.880 1277.810 372.940 ;
        RECT 1277.295 372.740 1277.810 372.880 ;
        RECT 1277.490 372.680 1277.810 372.740 ;
        RECT 1277.490 324.260 1277.810 324.320 ;
        RECT 1277.295 324.120 1277.810 324.260 ;
        RECT 1277.490 324.060 1277.810 324.120 ;
        RECT 1277.490 276.320 1277.810 276.380 ;
        RECT 1277.295 276.180 1277.810 276.320 ;
        RECT 1277.490 276.120 1277.810 276.180 ;
        RECT 1277.950 228.040 1278.270 228.100 ;
        RECT 1278.870 228.040 1279.190 228.100 ;
        RECT 1277.950 227.900 1279.190 228.040 ;
        RECT 1277.950 227.840 1278.270 227.900 ;
        RECT 1278.870 227.840 1279.190 227.900 ;
        RECT 1277.950 96.260 1278.270 96.520 ;
        RECT 1278.040 95.840 1278.180 96.260 ;
        RECT 1277.950 95.580 1278.270 95.840 ;
        RECT 1276.570 48.520 1276.890 48.580 ;
        RECT 1277.950 48.520 1278.270 48.580 ;
        RECT 1276.570 48.380 1278.270 48.520 ;
        RECT 1276.570 48.320 1276.890 48.380 ;
        RECT 1277.950 48.320 1278.270 48.380 ;
        RECT 258.130 30.840 258.450 30.900 ;
        RECT 1276.570 30.840 1276.890 30.900 ;
        RECT 258.130 30.700 1276.890 30.840 ;
        RECT 258.130 30.640 258.450 30.700 ;
        RECT 1276.570 30.640 1276.890 30.700 ;
      LAYER via ;
        RECT 1277.060 1586.820 1277.320 1587.080 ;
        RECT 1278.440 1586.480 1278.700 1586.740 ;
        RECT 1278.440 1579.680 1278.700 1579.940 ;
        RECT 1277.520 1490.600 1277.780 1490.860 ;
        RECT 1277.520 1463.060 1277.780 1463.320 ;
        RECT 1277.520 1462.380 1277.780 1462.640 ;
        RECT 1277.980 1173.040 1278.240 1173.300 ;
        RECT 1277.520 1172.700 1277.780 1172.960 ;
        RECT 1277.980 1076.480 1278.240 1076.740 ;
        RECT 1277.520 1076.140 1277.780 1076.400 ;
        RECT 1276.600 1055.400 1276.860 1055.660 ;
        RECT 1277.520 1055.400 1277.780 1055.660 ;
        RECT 1277.520 1007.120 1277.780 1007.380 ;
        RECT 1277.980 1007.120 1278.240 1007.380 ;
        RECT 1277.520 1000.320 1277.780 1000.580 ;
        RECT 1277.520 952.380 1277.780 952.640 ;
        RECT 1277.520 903.760 1277.780 904.020 ;
        RECT 1277.520 834.740 1277.780 835.000 ;
        RECT 1277.520 399.880 1277.780 400.140 ;
        RECT 1277.520 372.680 1277.780 372.940 ;
        RECT 1277.520 324.060 1277.780 324.320 ;
        RECT 1277.520 276.120 1277.780 276.380 ;
        RECT 1277.980 227.840 1278.240 228.100 ;
        RECT 1278.900 227.840 1279.160 228.100 ;
        RECT 1277.980 96.260 1278.240 96.520 ;
        RECT 1277.980 95.580 1278.240 95.840 ;
        RECT 1276.600 48.320 1276.860 48.580 ;
        RECT 1277.980 48.320 1278.240 48.580 ;
        RECT 258.160 30.640 258.420 30.900 ;
        RECT 1276.600 30.640 1276.860 30.900 ;
      LAYER met2 ;
        RECT 1281.580 1700.410 1281.860 1704.000 ;
        RECT 1279.420 1700.270 1281.860 1700.410 ;
        RECT 1279.420 1656.210 1279.560 1700.270 ;
        RECT 1281.580 1700.000 1281.860 1700.270 ;
        RECT 1277.580 1656.070 1279.560 1656.210 ;
        RECT 1277.580 1587.530 1277.720 1656.070 ;
        RECT 1277.120 1587.390 1277.720 1587.530 ;
        RECT 1277.120 1587.110 1277.260 1587.390 ;
        RECT 1277.060 1586.790 1277.320 1587.110 ;
        RECT 1278.440 1586.450 1278.700 1586.770 ;
        RECT 1278.500 1579.970 1278.640 1586.450 ;
        RECT 1278.440 1579.650 1278.700 1579.970 ;
        RECT 1277.520 1490.570 1277.780 1490.890 ;
        RECT 1277.580 1463.350 1277.720 1490.570 ;
        RECT 1277.520 1463.030 1277.780 1463.350 ;
        RECT 1277.520 1462.350 1277.780 1462.670 ;
        RECT 1277.580 1366.530 1277.720 1462.350 ;
        RECT 1277.120 1366.390 1277.720 1366.530 ;
        RECT 1277.120 1365.850 1277.260 1366.390 ;
        RECT 1277.120 1365.710 1277.720 1365.850 ;
        RECT 1277.580 1269.970 1277.720 1365.710 ;
        RECT 1277.120 1269.830 1277.720 1269.970 ;
        RECT 1277.120 1269.290 1277.260 1269.830 ;
        RECT 1277.120 1269.150 1277.720 1269.290 ;
        RECT 1277.580 1207.410 1277.720 1269.150 ;
        RECT 1277.580 1207.270 1278.180 1207.410 ;
        RECT 1278.040 1173.330 1278.180 1207.270 ;
        RECT 1277.980 1173.010 1278.240 1173.330 ;
        RECT 1277.520 1172.670 1277.780 1172.990 ;
        RECT 1277.580 1110.850 1277.720 1172.670 ;
        RECT 1277.580 1110.710 1278.180 1110.850 ;
        RECT 1278.040 1076.770 1278.180 1110.710 ;
        RECT 1277.980 1076.450 1278.240 1076.770 ;
        RECT 1277.520 1076.110 1277.780 1076.430 ;
        RECT 1277.580 1055.690 1277.720 1076.110 ;
        RECT 1276.600 1055.370 1276.860 1055.690 ;
        RECT 1277.520 1055.370 1277.780 1055.690 ;
        RECT 1276.660 1007.605 1276.800 1055.370 ;
        RECT 1276.590 1007.235 1276.870 1007.605 ;
        RECT 1277.520 1007.090 1277.780 1007.410 ;
        RECT 1277.970 1007.235 1278.250 1007.605 ;
        RECT 1277.980 1007.090 1278.240 1007.235 ;
        RECT 1277.580 1000.610 1277.720 1007.090 ;
        RECT 1277.520 1000.290 1277.780 1000.610 ;
        RECT 1277.520 952.350 1277.780 952.670 ;
        RECT 1277.580 904.050 1277.720 952.350 ;
        RECT 1277.520 903.730 1277.780 904.050 ;
        RECT 1277.520 834.710 1277.780 835.030 ;
        RECT 1277.580 690.610 1277.720 834.710 ;
        RECT 1277.120 690.470 1277.720 690.610 ;
        RECT 1277.120 689.930 1277.260 690.470 ;
        RECT 1277.120 689.790 1277.720 689.930 ;
        RECT 1277.580 497.490 1277.720 689.790 ;
        RECT 1277.120 497.350 1277.720 497.490 ;
        RECT 1277.120 496.810 1277.260 497.350 ;
        RECT 1277.120 496.670 1277.720 496.810 ;
        RECT 1277.580 400.170 1277.720 496.670 ;
        RECT 1277.520 399.850 1277.780 400.170 ;
        RECT 1277.520 372.650 1277.780 372.970 ;
        RECT 1277.580 324.350 1277.720 372.650 ;
        RECT 1277.520 324.030 1277.780 324.350 ;
        RECT 1277.520 276.090 1277.780 276.410 ;
        RECT 1277.580 275.925 1277.720 276.090 ;
        RECT 1277.510 275.555 1277.790 275.925 ;
        RECT 1278.890 275.555 1279.170 275.925 ;
        RECT 1278.960 228.130 1279.100 275.555 ;
        RECT 1277.980 227.810 1278.240 228.130 ;
        RECT 1278.900 227.810 1279.160 228.130 ;
        RECT 1278.040 96.550 1278.180 227.810 ;
        RECT 1277.980 96.230 1278.240 96.550 ;
        RECT 1277.980 95.550 1278.240 95.870 ;
        RECT 1278.040 48.610 1278.180 95.550 ;
        RECT 1276.600 48.290 1276.860 48.610 ;
        RECT 1277.980 48.290 1278.240 48.610 ;
        RECT 1276.660 30.930 1276.800 48.290 ;
        RECT 258.160 30.610 258.420 30.930 ;
        RECT 1276.600 30.610 1276.860 30.930 ;
        RECT 258.220 2.400 258.360 30.610 ;
        RECT 258.010 -4.800 258.570 2.400 ;
      LAYER via2 ;
        RECT 1276.590 1007.280 1276.870 1007.560 ;
        RECT 1277.970 1007.280 1278.250 1007.560 ;
        RECT 1277.510 275.600 1277.790 275.880 ;
        RECT 1278.890 275.600 1279.170 275.880 ;
      LAYER met3 ;
        RECT 1276.565 1007.570 1276.895 1007.585 ;
        RECT 1277.945 1007.570 1278.275 1007.585 ;
        RECT 1276.565 1007.270 1278.275 1007.570 ;
        RECT 1276.565 1007.255 1276.895 1007.270 ;
        RECT 1277.945 1007.255 1278.275 1007.270 ;
        RECT 1277.485 275.890 1277.815 275.905 ;
        RECT 1278.865 275.890 1279.195 275.905 ;
        RECT 1277.485 275.590 1279.195 275.890 ;
        RECT 1277.485 275.575 1277.815 275.590 ;
        RECT 1278.865 275.575 1279.195 275.590 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 276.070 31.180 276.390 31.240 ;
        RECT 1291.290 31.180 1291.610 31.240 ;
        RECT 276.070 31.040 1291.610 31.180 ;
        RECT 276.070 30.980 276.390 31.040 ;
        RECT 1291.290 30.980 1291.610 31.040 ;
      LAYER via ;
        RECT 276.100 30.980 276.360 31.240 ;
        RECT 1291.320 30.980 1291.580 31.240 ;
      LAYER met2 ;
        RECT 1290.780 1700.410 1291.060 1704.000 ;
        RECT 1290.780 1700.270 1291.520 1700.410 ;
        RECT 1290.780 1700.000 1291.060 1700.270 ;
        RECT 1291.380 31.270 1291.520 1700.270 ;
        RECT 276.100 30.950 276.360 31.270 ;
        RECT 1291.320 30.950 1291.580 31.270 ;
        RECT 276.160 2.400 276.300 30.950 ;
        RECT 275.950 -4.800 276.510 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 294.010 31.520 294.330 31.580 ;
        RECT 1297.270 31.520 1297.590 31.580 ;
        RECT 294.010 31.380 1297.590 31.520 ;
        RECT 294.010 31.320 294.330 31.380 ;
        RECT 1297.270 31.320 1297.590 31.380 ;
      LAYER via ;
        RECT 294.040 31.320 294.300 31.580 ;
        RECT 1297.300 31.320 1297.560 31.580 ;
      LAYER met2 ;
        RECT 1299.980 1700.410 1300.260 1704.000 ;
        RECT 1297.360 1700.270 1300.260 1700.410 ;
        RECT 1297.360 31.610 1297.500 1700.270 ;
        RECT 1299.980 1700.000 1300.260 1700.270 ;
        RECT 294.040 31.290 294.300 31.610 ;
        RECT 1297.300 31.290 1297.560 31.610 ;
        RECT 294.100 2.400 294.240 31.290 ;
        RECT 293.890 -4.800 294.450 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1305.090 1608.240 1305.410 1608.500 ;
        RECT 1305.180 1607.820 1305.320 1608.240 ;
        RECT 1305.090 1607.560 1305.410 1607.820 ;
        RECT 1305.090 1539.080 1305.410 1539.140 ;
        RECT 1305.550 1539.080 1305.870 1539.140 ;
        RECT 1305.090 1538.940 1305.870 1539.080 ;
        RECT 1305.090 1538.880 1305.410 1538.940 ;
        RECT 1305.550 1538.880 1305.870 1538.940 ;
        RECT 1305.090 1490.800 1305.410 1490.860 ;
        RECT 1306.010 1490.800 1306.330 1490.860 ;
        RECT 1305.090 1490.660 1306.330 1490.800 ;
        RECT 1305.090 1490.600 1305.410 1490.660 ;
        RECT 1306.010 1490.600 1306.330 1490.660 ;
        RECT 1305.090 1269.940 1305.410 1270.200 ;
        RECT 1305.180 1269.520 1305.320 1269.940 ;
        RECT 1305.090 1269.260 1305.410 1269.520 ;
        RECT 1305.550 1173.240 1305.870 1173.300 ;
        RECT 1305.180 1173.100 1305.870 1173.240 ;
        RECT 1305.180 1172.960 1305.320 1173.100 ;
        RECT 1305.550 1173.040 1305.870 1173.100 ;
        RECT 1305.090 1172.700 1305.410 1172.960 ;
        RECT 1305.550 1076.680 1305.870 1076.740 ;
        RECT 1305.180 1076.540 1305.870 1076.680 ;
        RECT 1305.180 1076.400 1305.320 1076.540 ;
        RECT 1305.550 1076.480 1305.870 1076.540 ;
        RECT 1305.090 1076.140 1305.410 1076.400 ;
        RECT 1305.090 255.380 1305.410 255.640 ;
        RECT 1305.180 254.960 1305.320 255.380 ;
        RECT 1305.090 254.700 1305.410 254.960 ;
        RECT 1305.090 145.420 1305.410 145.480 ;
        RECT 1304.720 145.280 1305.410 145.420 ;
        RECT 1304.720 145.140 1304.860 145.280 ;
        RECT 1305.090 145.220 1305.410 145.280 ;
        RECT 1304.630 144.880 1304.950 145.140 ;
        RECT 1304.630 96.800 1304.950 96.860 ;
        RECT 1305.090 96.800 1305.410 96.860 ;
        RECT 1304.630 96.660 1305.410 96.800 ;
        RECT 1304.630 96.600 1304.950 96.660 ;
        RECT 1305.090 96.600 1305.410 96.660 ;
        RECT 311.950 32.200 312.270 32.260 ;
        RECT 1304.630 32.200 1304.950 32.260 ;
        RECT 311.950 32.060 1304.950 32.200 ;
        RECT 311.950 32.000 312.270 32.060 ;
        RECT 1304.630 32.000 1304.950 32.060 ;
      LAYER via ;
        RECT 1305.120 1608.240 1305.380 1608.500 ;
        RECT 1305.120 1607.560 1305.380 1607.820 ;
        RECT 1305.120 1538.880 1305.380 1539.140 ;
        RECT 1305.580 1538.880 1305.840 1539.140 ;
        RECT 1305.120 1490.600 1305.380 1490.860 ;
        RECT 1306.040 1490.600 1306.300 1490.860 ;
        RECT 1305.120 1269.940 1305.380 1270.200 ;
        RECT 1305.120 1269.260 1305.380 1269.520 ;
        RECT 1305.580 1173.040 1305.840 1173.300 ;
        RECT 1305.120 1172.700 1305.380 1172.960 ;
        RECT 1305.580 1076.480 1305.840 1076.740 ;
        RECT 1305.120 1076.140 1305.380 1076.400 ;
        RECT 1305.120 255.380 1305.380 255.640 ;
        RECT 1305.120 254.700 1305.380 254.960 ;
        RECT 1305.120 145.220 1305.380 145.480 ;
        RECT 1304.660 144.880 1304.920 145.140 ;
        RECT 1304.660 96.600 1304.920 96.860 ;
        RECT 1305.120 96.600 1305.380 96.860 ;
        RECT 311.980 32.000 312.240 32.260 ;
        RECT 1304.660 32.000 1304.920 32.260 ;
      LAYER met2 ;
        RECT 1309.180 1701.090 1309.460 1704.000 ;
        RECT 1306.560 1700.950 1309.460 1701.090 ;
        RECT 1306.560 1677.970 1306.700 1700.950 ;
        RECT 1309.180 1700.000 1309.460 1700.950 ;
        RECT 1305.180 1677.830 1306.700 1677.970 ;
        RECT 1305.180 1608.530 1305.320 1677.830 ;
        RECT 1305.120 1608.210 1305.380 1608.530 ;
        RECT 1305.120 1607.530 1305.380 1607.850 ;
        RECT 1305.180 1595.125 1305.320 1607.530 ;
        RECT 1305.110 1594.755 1305.390 1595.125 ;
        RECT 1305.110 1594.075 1305.390 1594.445 ;
        RECT 1305.180 1559.650 1305.320 1594.075 ;
        RECT 1305.180 1559.510 1305.780 1559.650 ;
        RECT 1305.640 1539.170 1305.780 1559.510 ;
        RECT 1305.120 1538.850 1305.380 1539.170 ;
        RECT 1305.580 1538.850 1305.840 1539.170 ;
        RECT 1305.180 1538.685 1305.320 1538.850 ;
        RECT 1305.110 1538.315 1305.390 1538.685 ;
        RECT 1306.030 1538.315 1306.310 1538.685 ;
        RECT 1306.100 1490.890 1306.240 1538.315 ;
        RECT 1305.120 1490.570 1305.380 1490.890 ;
        RECT 1306.040 1490.570 1306.300 1490.890 ;
        RECT 1305.180 1490.290 1305.320 1490.570 ;
        RECT 1305.180 1490.150 1305.780 1490.290 ;
        RECT 1305.640 1461.730 1305.780 1490.150 ;
        RECT 1305.180 1461.590 1305.780 1461.730 ;
        RECT 1305.180 1400.700 1305.320 1461.590 ;
        RECT 1304.260 1400.560 1305.320 1400.700 ;
        RECT 1304.260 1364.490 1304.400 1400.560 ;
        RECT 1304.260 1364.350 1305.320 1364.490 ;
        RECT 1305.180 1270.230 1305.320 1364.350 ;
        RECT 1305.120 1269.910 1305.380 1270.230 ;
        RECT 1305.120 1269.230 1305.380 1269.550 ;
        RECT 1305.180 1207.410 1305.320 1269.230 ;
        RECT 1305.180 1207.270 1305.780 1207.410 ;
        RECT 1305.640 1173.330 1305.780 1207.270 ;
        RECT 1305.580 1173.010 1305.840 1173.330 ;
        RECT 1305.120 1172.670 1305.380 1172.990 ;
        RECT 1305.180 1110.850 1305.320 1172.670 ;
        RECT 1305.180 1110.710 1305.780 1110.850 ;
        RECT 1305.640 1076.770 1305.780 1110.710 ;
        RECT 1305.580 1076.450 1305.840 1076.770 ;
        RECT 1305.120 1076.110 1305.380 1076.430 ;
        RECT 1305.180 893.930 1305.320 1076.110 ;
        RECT 1304.720 893.790 1305.320 893.930 ;
        RECT 1304.720 834.770 1304.860 893.790 ;
        RECT 1304.720 834.630 1305.320 834.770 ;
        RECT 1305.180 497.490 1305.320 834.630 ;
        RECT 1304.720 497.350 1305.320 497.490 ;
        RECT 1304.720 496.810 1304.860 497.350 ;
        RECT 1304.720 496.670 1305.320 496.810 ;
        RECT 1305.180 400.930 1305.320 496.670 ;
        RECT 1305.180 400.790 1305.780 400.930 ;
        RECT 1305.640 399.570 1305.780 400.790 ;
        RECT 1305.180 399.430 1305.780 399.570 ;
        RECT 1305.180 303.690 1305.320 399.430 ;
        RECT 1304.720 303.550 1305.320 303.690 ;
        RECT 1304.720 303.010 1304.860 303.550 ;
        RECT 1304.720 302.870 1305.320 303.010 ;
        RECT 1305.180 255.670 1305.320 302.870 ;
        RECT 1305.120 255.350 1305.380 255.670 ;
        RECT 1305.120 254.670 1305.380 254.990 ;
        RECT 1305.180 145.510 1305.320 254.670 ;
        RECT 1305.120 145.190 1305.380 145.510 ;
        RECT 1304.660 144.850 1304.920 145.170 ;
        RECT 1304.720 96.890 1304.860 144.850 ;
        RECT 1304.660 96.570 1304.920 96.890 ;
        RECT 1305.120 96.570 1305.380 96.890 ;
        RECT 1305.180 60.930 1305.320 96.570 ;
        RECT 1304.720 60.790 1305.320 60.930 ;
        RECT 1304.720 32.290 1304.860 60.790 ;
        RECT 311.980 31.970 312.240 32.290 ;
        RECT 1304.660 31.970 1304.920 32.290 ;
        RECT 312.040 2.400 312.180 31.970 ;
        RECT 311.830 -4.800 312.390 2.400 ;
      LAYER via2 ;
        RECT 1305.110 1594.800 1305.390 1595.080 ;
        RECT 1305.110 1594.120 1305.390 1594.400 ;
        RECT 1305.110 1538.360 1305.390 1538.640 ;
        RECT 1306.030 1538.360 1306.310 1538.640 ;
      LAYER met3 ;
        RECT 1305.085 1595.090 1305.415 1595.105 ;
        RECT 1304.870 1594.775 1305.415 1595.090 ;
        RECT 1304.870 1594.425 1305.170 1594.775 ;
        RECT 1304.870 1594.110 1305.415 1594.425 ;
        RECT 1305.085 1594.095 1305.415 1594.110 ;
        RECT 1305.085 1538.650 1305.415 1538.665 ;
        RECT 1306.005 1538.650 1306.335 1538.665 ;
        RECT 1305.085 1538.350 1306.335 1538.650 ;
        RECT 1305.085 1538.335 1305.415 1538.350 ;
        RECT 1306.005 1538.335 1306.335 1538.350 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 329.890 31.860 330.210 31.920 ;
        RECT 1318.430 31.860 1318.750 31.920 ;
        RECT 329.890 31.720 1318.750 31.860 ;
        RECT 329.890 31.660 330.210 31.720 ;
        RECT 1318.430 31.660 1318.750 31.720 ;
      LAYER via ;
        RECT 329.920 31.660 330.180 31.920 ;
        RECT 1318.460 31.660 1318.720 31.920 ;
      LAYER met2 ;
        RECT 1318.380 1700.000 1318.660 1704.000 ;
        RECT 1318.520 31.950 1318.660 1700.000 ;
        RECT 329.920 31.630 330.180 31.950 ;
        RECT 1318.460 31.630 1318.720 31.950 ;
        RECT 329.980 2.400 330.120 31.630 ;
        RECT 329.770 -4.800 330.330 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 347.370 32.540 347.690 32.600 ;
        RECT 1324.870 32.540 1325.190 32.600 ;
        RECT 347.370 32.400 1325.190 32.540 ;
        RECT 347.370 32.340 347.690 32.400 ;
        RECT 1324.870 32.340 1325.190 32.400 ;
      LAYER via ;
        RECT 347.400 32.340 347.660 32.600 ;
        RECT 1324.900 32.340 1325.160 32.600 ;
      LAYER met2 ;
        RECT 1327.120 1700.410 1327.400 1704.000 ;
        RECT 1324.960 1700.270 1327.400 1700.410 ;
        RECT 1324.960 32.630 1325.100 1700.270 ;
        RECT 1327.120 1700.000 1327.400 1700.270 ;
        RECT 347.400 32.310 347.660 32.630 ;
        RECT 1324.900 32.310 1325.160 32.630 ;
        RECT 347.460 2.400 347.600 32.310 ;
        RECT 347.250 -4.800 347.810 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1332.305 462.485 1332.475 510.595 ;
        RECT 1332.305 324.445 1332.475 389.895 ;
        RECT 1333.225 95.965 1333.395 137.955 ;
      LAYER mcon ;
        RECT 1332.305 510.425 1332.475 510.595 ;
        RECT 1332.305 389.725 1332.475 389.895 ;
        RECT 1333.225 137.785 1333.395 137.955 ;
      LAYER met1 ;
        RECT 1332.230 869.620 1332.550 869.680 ;
        RECT 1332.690 869.620 1333.010 869.680 ;
        RECT 1332.230 869.480 1333.010 869.620 ;
        RECT 1332.230 869.420 1332.550 869.480 ;
        RECT 1332.690 869.420 1333.010 869.480 ;
        RECT 1332.690 773.060 1333.010 773.120 ;
        RECT 1333.150 773.060 1333.470 773.120 ;
        RECT 1332.690 772.920 1333.470 773.060 ;
        RECT 1332.690 772.860 1333.010 772.920 ;
        RECT 1333.150 772.860 1333.470 772.920 ;
        RECT 1332.230 717.640 1332.550 717.700 ;
        RECT 1333.610 717.640 1333.930 717.700 ;
        RECT 1332.230 717.500 1333.930 717.640 ;
        RECT 1332.230 717.440 1332.550 717.500 ;
        RECT 1333.610 717.440 1333.930 717.500 ;
        RECT 1333.150 614.280 1333.470 614.340 ;
        RECT 1333.610 614.280 1333.930 614.340 ;
        RECT 1333.150 614.140 1333.930 614.280 ;
        RECT 1333.150 614.080 1333.470 614.140 ;
        RECT 1333.610 614.080 1333.930 614.140 ;
        RECT 1332.245 510.580 1332.535 510.625 ;
        RECT 1332.690 510.580 1333.010 510.640 ;
        RECT 1332.245 510.440 1333.010 510.580 ;
        RECT 1332.245 510.395 1332.535 510.440 ;
        RECT 1332.690 510.380 1333.010 510.440 ;
        RECT 1332.230 462.640 1332.550 462.700 ;
        RECT 1332.035 462.500 1332.550 462.640 ;
        RECT 1332.230 462.440 1332.550 462.500 ;
        RECT 1332.245 389.880 1332.535 389.925 ;
        RECT 1333.150 389.880 1333.470 389.940 ;
        RECT 1332.245 389.740 1333.470 389.880 ;
        RECT 1332.245 389.695 1332.535 389.740 ;
        RECT 1333.150 389.680 1333.470 389.740 ;
        RECT 1332.230 324.600 1332.550 324.660 ;
        RECT 1332.035 324.460 1332.550 324.600 ;
        RECT 1332.230 324.400 1332.550 324.460 ;
        RECT 1332.690 144.740 1333.010 144.800 ;
        RECT 1333.150 144.740 1333.470 144.800 ;
        RECT 1332.690 144.600 1333.470 144.740 ;
        RECT 1332.690 144.540 1333.010 144.600 ;
        RECT 1333.150 144.540 1333.470 144.600 ;
        RECT 1333.150 137.940 1333.470 138.000 ;
        RECT 1332.955 137.800 1333.470 137.940 ;
        RECT 1333.150 137.740 1333.470 137.800 ;
        RECT 1333.150 96.120 1333.470 96.180 ;
        RECT 1332.955 95.980 1333.470 96.120 ;
        RECT 1333.150 95.920 1333.470 95.980 ;
        RECT 365.310 32.880 365.630 32.940 ;
        RECT 1331.770 32.880 1332.090 32.940 ;
        RECT 365.310 32.740 1332.090 32.880 ;
        RECT 365.310 32.680 365.630 32.740 ;
        RECT 1331.770 32.680 1332.090 32.740 ;
      LAYER via ;
        RECT 1332.260 869.420 1332.520 869.680 ;
        RECT 1332.720 869.420 1332.980 869.680 ;
        RECT 1332.720 772.860 1332.980 773.120 ;
        RECT 1333.180 772.860 1333.440 773.120 ;
        RECT 1332.260 717.440 1332.520 717.700 ;
        RECT 1333.640 717.440 1333.900 717.700 ;
        RECT 1333.180 614.080 1333.440 614.340 ;
        RECT 1333.640 614.080 1333.900 614.340 ;
        RECT 1332.720 510.380 1332.980 510.640 ;
        RECT 1332.260 462.440 1332.520 462.700 ;
        RECT 1333.180 389.680 1333.440 389.940 ;
        RECT 1332.260 324.400 1332.520 324.660 ;
        RECT 1332.720 144.540 1332.980 144.800 ;
        RECT 1333.180 144.540 1333.440 144.800 ;
        RECT 1333.180 137.740 1333.440 138.000 ;
        RECT 1333.180 95.920 1333.440 96.180 ;
        RECT 365.340 32.680 365.600 32.940 ;
        RECT 1331.800 32.680 1332.060 32.940 ;
      LAYER met2 ;
        RECT 1336.320 1701.090 1336.600 1704.000 ;
        RECT 1334.160 1700.950 1336.600 1701.090 ;
        RECT 1334.160 1677.970 1334.300 1700.950 ;
        RECT 1336.320 1700.000 1336.600 1700.950 ;
        RECT 1332.780 1677.830 1334.300 1677.970 ;
        RECT 1332.780 1607.930 1332.920 1677.830 ;
        RECT 1332.320 1607.790 1332.920 1607.930 ;
        RECT 1332.320 1607.250 1332.460 1607.790 ;
        RECT 1332.320 1607.110 1332.920 1607.250 ;
        RECT 1332.780 1463.090 1332.920 1607.110 ;
        RECT 1332.320 1462.950 1332.920 1463.090 ;
        RECT 1332.320 1462.410 1332.460 1462.950 ;
        RECT 1332.320 1462.270 1332.920 1462.410 ;
        RECT 1332.780 869.710 1332.920 1462.270 ;
        RECT 1332.260 869.565 1332.520 869.710 ;
        RECT 1332.250 869.195 1332.530 869.565 ;
        RECT 1332.720 869.390 1332.980 869.710 ;
        RECT 1333.170 869.195 1333.450 869.565 ;
        RECT 1333.240 773.150 1333.380 869.195 ;
        RECT 1332.720 772.830 1332.980 773.150 ;
        RECT 1333.180 772.830 1333.440 773.150 ;
        RECT 1332.780 725.405 1332.920 772.830 ;
        RECT 1332.710 725.035 1332.990 725.405 ;
        RECT 1332.250 724.355 1332.530 724.725 ;
        RECT 1332.320 717.730 1332.460 724.355 ;
        RECT 1332.260 717.410 1332.520 717.730 ;
        RECT 1333.640 717.410 1333.900 717.730 ;
        RECT 1333.700 614.370 1333.840 717.410 ;
        RECT 1333.180 614.050 1333.440 614.370 ;
        RECT 1333.640 614.050 1333.900 614.370 ;
        RECT 1333.240 566.170 1333.380 614.050 ;
        RECT 1332.320 566.030 1333.380 566.170 ;
        RECT 1332.320 545.770 1332.460 566.030 ;
        RECT 1332.320 545.630 1333.380 545.770 ;
        RECT 1333.240 517.890 1333.380 545.630 ;
        RECT 1332.780 517.750 1333.380 517.890 ;
        RECT 1332.780 510.670 1332.920 517.750 ;
        RECT 1332.720 510.350 1332.980 510.670 ;
        RECT 1332.260 462.410 1332.520 462.730 ;
        RECT 1332.320 413.965 1332.460 462.410 ;
        RECT 1332.250 413.595 1332.530 413.965 ;
        RECT 1333.170 412.915 1333.450 413.285 ;
        RECT 1333.240 389.970 1333.380 412.915 ;
        RECT 1333.180 389.650 1333.440 389.970 ;
        RECT 1332.260 324.370 1332.520 324.690 ;
        RECT 1332.320 258.810 1332.460 324.370 ;
        RECT 1332.320 258.670 1332.920 258.810 ;
        RECT 1332.780 144.830 1332.920 258.670 ;
        RECT 1332.720 144.510 1332.980 144.830 ;
        RECT 1333.180 144.510 1333.440 144.830 ;
        RECT 1333.240 138.030 1333.380 144.510 ;
        RECT 1333.180 137.710 1333.440 138.030 ;
        RECT 1333.180 95.890 1333.440 96.210 ;
        RECT 1333.240 72.490 1333.380 95.890 ;
        RECT 1331.860 72.350 1333.380 72.490 ;
        RECT 1331.860 32.970 1332.000 72.350 ;
        RECT 365.340 32.650 365.600 32.970 ;
        RECT 1331.800 32.650 1332.060 32.970 ;
        RECT 365.400 2.400 365.540 32.650 ;
        RECT 365.190 -4.800 365.750 2.400 ;
      LAYER via2 ;
        RECT 1332.250 869.240 1332.530 869.520 ;
        RECT 1333.170 869.240 1333.450 869.520 ;
        RECT 1332.710 725.080 1332.990 725.360 ;
        RECT 1332.250 724.400 1332.530 724.680 ;
        RECT 1332.250 413.640 1332.530 413.920 ;
        RECT 1333.170 412.960 1333.450 413.240 ;
      LAYER met3 ;
        RECT 1332.225 869.530 1332.555 869.545 ;
        RECT 1333.145 869.530 1333.475 869.545 ;
        RECT 1332.225 869.230 1333.475 869.530 ;
        RECT 1332.225 869.215 1332.555 869.230 ;
        RECT 1333.145 869.215 1333.475 869.230 ;
        RECT 1332.685 725.370 1333.015 725.385 ;
        RECT 1331.550 725.070 1333.015 725.370 ;
        RECT 1331.550 724.690 1331.850 725.070 ;
        RECT 1332.685 725.055 1333.015 725.070 ;
        RECT 1332.225 724.690 1332.555 724.705 ;
        RECT 1331.550 724.390 1332.555 724.690 ;
        RECT 1332.225 724.375 1332.555 724.390 ;
        RECT 1332.225 413.930 1332.555 413.945 ;
        RECT 1331.550 413.630 1332.555 413.930 ;
        RECT 1331.550 413.250 1331.850 413.630 ;
        RECT 1332.225 413.615 1332.555 413.630 ;
        RECT 1333.145 413.250 1333.475 413.265 ;
        RECT 1331.550 412.950 1333.475 413.250 ;
        RECT 1333.145 412.935 1333.475 412.950 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 383.250 33.220 383.570 33.280 ;
        RECT 1345.570 33.220 1345.890 33.280 ;
        RECT 383.250 33.080 1345.890 33.220 ;
        RECT 383.250 33.020 383.570 33.080 ;
        RECT 1345.570 33.020 1345.890 33.080 ;
      LAYER via ;
        RECT 383.280 33.020 383.540 33.280 ;
        RECT 1345.600 33.020 1345.860 33.280 ;
      LAYER met2 ;
        RECT 1345.520 1700.000 1345.800 1704.000 ;
        RECT 1345.660 33.310 1345.800 1700.000 ;
        RECT 383.280 32.990 383.540 33.310 ;
        RECT 1345.600 32.990 1345.860 33.310 ;
        RECT 383.340 2.400 383.480 32.990 ;
        RECT 383.130 -4.800 383.690 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 401.190 33.560 401.510 33.620 ;
        RECT 1352.930 33.560 1353.250 33.620 ;
        RECT 401.190 33.420 1353.250 33.560 ;
        RECT 401.190 33.360 401.510 33.420 ;
        RECT 1352.930 33.360 1353.250 33.420 ;
      LAYER via ;
        RECT 401.220 33.360 401.480 33.620 ;
        RECT 1352.960 33.360 1353.220 33.620 ;
      LAYER met2 ;
        RECT 1354.720 1700.410 1355.000 1704.000 ;
        RECT 1352.560 1700.270 1355.000 1700.410 ;
        RECT 1352.560 48.010 1352.700 1700.270 ;
        RECT 1354.720 1700.000 1355.000 1700.270 ;
        RECT 1352.560 47.870 1353.160 48.010 ;
        RECT 1353.020 33.650 1353.160 47.870 ;
        RECT 401.220 33.330 401.480 33.650 ;
        RECT 1352.960 33.330 1353.220 33.650 ;
        RECT 401.280 2.400 401.420 33.330 ;
        RECT 401.070 -4.800 401.630 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 62.170 25.400 62.490 25.460 ;
        RECT 1180.430 25.400 1180.750 25.460 ;
        RECT 62.170 25.260 1180.750 25.400 ;
        RECT 62.170 25.200 62.490 25.260 ;
        RECT 1180.430 25.200 1180.750 25.260 ;
      LAYER via ;
        RECT 62.200 25.200 62.460 25.460 ;
        RECT 1180.460 25.200 1180.720 25.460 ;
      LAYER met2 ;
        RECT 1180.380 1700.000 1180.660 1704.000 ;
        RECT 1180.520 25.490 1180.660 1700.000 ;
        RECT 62.200 25.170 62.460 25.490 ;
        RECT 1180.460 25.170 1180.720 25.490 ;
        RECT 62.260 2.400 62.400 25.170 ;
        RECT 62.050 -4.800 62.610 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1360.365 1256.045 1360.535 1304.155 ;
        RECT 1359.905 917.745 1360.075 932.195 ;
        RECT 1359.905 814.385 1360.075 862.495 ;
        RECT 1359.905 742.985 1360.075 790.075 ;
        RECT 1359.905 576.725 1360.075 620.755 ;
        RECT 1359.905 365.925 1360.075 414.035 ;
        RECT 1359.905 234.685 1360.075 258.995 ;
        RECT 1360.365 144.925 1360.535 214.795 ;
      LAYER mcon ;
        RECT 1360.365 1303.985 1360.535 1304.155 ;
        RECT 1359.905 932.025 1360.075 932.195 ;
        RECT 1359.905 862.325 1360.075 862.495 ;
        RECT 1359.905 789.905 1360.075 790.075 ;
        RECT 1359.905 620.585 1360.075 620.755 ;
        RECT 1359.905 413.865 1360.075 414.035 ;
        RECT 1359.905 258.825 1360.075 258.995 ;
        RECT 1360.365 214.625 1360.535 214.795 ;
      LAYER met1 ;
        RECT 1360.290 1365.820 1360.610 1366.080 ;
        RECT 1360.380 1365.400 1360.520 1365.820 ;
        RECT 1360.290 1365.140 1360.610 1365.400 ;
        RECT 1360.290 1304.140 1360.610 1304.200 ;
        RECT 1360.095 1304.000 1360.610 1304.140 ;
        RECT 1360.290 1303.940 1360.610 1304.000 ;
        RECT 1360.290 1256.200 1360.610 1256.260 ;
        RECT 1360.095 1256.060 1360.610 1256.200 ;
        RECT 1360.290 1256.000 1360.610 1256.060 ;
        RECT 1359.370 1159.300 1359.690 1159.360 ;
        RECT 1360.290 1159.300 1360.610 1159.360 ;
        RECT 1359.370 1159.160 1360.610 1159.300 ;
        RECT 1359.370 1159.100 1359.690 1159.160 ;
        RECT 1360.290 1159.100 1360.610 1159.160 ;
        RECT 1359.370 1062.740 1359.690 1062.800 ;
        RECT 1360.290 1062.740 1360.610 1062.800 ;
        RECT 1359.370 1062.600 1360.610 1062.740 ;
        RECT 1359.370 1062.540 1359.690 1062.600 ;
        RECT 1360.290 1062.540 1360.610 1062.600 ;
        RECT 1359.845 932.180 1360.135 932.225 ;
        RECT 1360.290 932.180 1360.610 932.240 ;
        RECT 1359.845 932.040 1360.610 932.180 ;
        RECT 1359.845 931.995 1360.135 932.040 ;
        RECT 1360.290 931.980 1360.610 932.040 ;
        RECT 1359.830 917.900 1360.150 917.960 ;
        RECT 1359.635 917.760 1360.150 917.900 ;
        RECT 1359.830 917.700 1360.150 917.760 ;
        RECT 1359.830 869.620 1360.150 869.680 ;
        RECT 1360.290 869.620 1360.610 869.680 ;
        RECT 1359.830 869.480 1360.610 869.620 ;
        RECT 1359.830 869.420 1360.150 869.480 ;
        RECT 1360.290 869.420 1360.610 869.480 ;
        RECT 1359.845 862.480 1360.135 862.525 ;
        RECT 1360.290 862.480 1360.610 862.540 ;
        RECT 1359.845 862.340 1360.610 862.480 ;
        RECT 1359.845 862.295 1360.135 862.340 ;
        RECT 1360.290 862.280 1360.610 862.340 ;
        RECT 1359.830 814.540 1360.150 814.600 ;
        RECT 1359.635 814.400 1360.150 814.540 ;
        RECT 1359.830 814.340 1360.150 814.400 ;
        RECT 1359.830 790.060 1360.150 790.120 ;
        RECT 1359.635 789.920 1360.150 790.060 ;
        RECT 1359.830 789.860 1360.150 789.920 ;
        RECT 1359.830 743.140 1360.150 743.200 ;
        RECT 1359.635 743.000 1360.150 743.140 ;
        RECT 1359.830 742.940 1360.150 743.000 ;
        RECT 1359.830 724.440 1360.150 724.500 ;
        RECT 1360.290 724.440 1360.610 724.500 ;
        RECT 1359.830 724.300 1360.610 724.440 ;
        RECT 1359.830 724.240 1360.150 724.300 ;
        RECT 1360.290 724.240 1360.610 724.300 ;
        RECT 1359.370 676.160 1359.690 676.220 ;
        RECT 1359.830 676.160 1360.150 676.220 ;
        RECT 1359.370 676.020 1360.150 676.160 ;
        RECT 1359.370 675.960 1359.690 676.020 ;
        RECT 1359.830 675.960 1360.150 676.020 ;
        RECT 1359.830 627.880 1360.150 627.940 ;
        RECT 1360.290 627.880 1360.610 627.940 ;
        RECT 1359.830 627.740 1360.610 627.880 ;
        RECT 1359.830 627.680 1360.150 627.740 ;
        RECT 1360.290 627.680 1360.610 627.740 ;
        RECT 1359.830 620.740 1360.150 620.800 ;
        RECT 1359.635 620.600 1360.150 620.740 ;
        RECT 1359.830 620.540 1360.150 620.600 ;
        RECT 1359.830 576.880 1360.150 576.940 ;
        RECT 1359.635 576.740 1360.150 576.880 ;
        RECT 1359.830 576.680 1360.150 576.740 ;
        RECT 1359.370 524.520 1359.690 524.580 ;
        RECT 1359.830 524.520 1360.150 524.580 ;
        RECT 1359.370 524.380 1360.150 524.520 ;
        RECT 1359.370 524.320 1359.690 524.380 ;
        RECT 1359.830 524.320 1360.150 524.380 ;
        RECT 1359.370 496.640 1359.690 496.700 ;
        RECT 1360.290 496.640 1360.610 496.700 ;
        RECT 1359.370 496.500 1360.610 496.640 ;
        RECT 1359.370 496.440 1359.690 496.500 ;
        RECT 1360.290 496.440 1360.610 496.500 ;
        RECT 1360.290 421.500 1360.610 421.560 ;
        RECT 1359.920 421.360 1360.610 421.500 ;
        RECT 1359.920 421.220 1360.060 421.360 ;
        RECT 1360.290 421.300 1360.610 421.360 ;
        RECT 1359.830 420.960 1360.150 421.220 ;
        RECT 1359.830 414.020 1360.150 414.080 ;
        RECT 1359.635 413.880 1360.150 414.020 ;
        RECT 1359.830 413.820 1360.150 413.880 ;
        RECT 1359.830 366.080 1360.150 366.140 ;
        RECT 1359.635 365.940 1360.150 366.080 ;
        RECT 1359.830 365.880 1360.150 365.940 ;
        RECT 1359.830 324.260 1360.150 324.320 ;
        RECT 1360.290 324.260 1360.610 324.320 ;
        RECT 1359.830 324.120 1360.610 324.260 ;
        RECT 1359.830 324.060 1360.150 324.120 ;
        RECT 1360.290 324.060 1360.610 324.120 ;
        RECT 1359.845 258.980 1360.135 259.025 ;
        RECT 1360.290 258.980 1360.610 259.040 ;
        RECT 1359.845 258.840 1360.610 258.980 ;
        RECT 1359.845 258.795 1360.135 258.840 ;
        RECT 1360.290 258.780 1360.610 258.840 ;
        RECT 1359.830 234.840 1360.150 234.900 ;
        RECT 1359.635 234.700 1360.150 234.840 ;
        RECT 1359.830 234.640 1360.150 234.700 ;
        RECT 1359.830 214.780 1360.150 214.840 ;
        RECT 1360.305 214.780 1360.595 214.825 ;
        RECT 1359.830 214.640 1360.595 214.780 ;
        RECT 1359.830 214.580 1360.150 214.640 ;
        RECT 1360.305 214.595 1360.595 214.640 ;
        RECT 1360.290 145.080 1360.610 145.140 ;
        RECT 1360.095 144.940 1360.610 145.080 ;
        RECT 1360.290 144.880 1360.610 144.940 ;
        RECT 1360.290 90.340 1360.610 90.400 ;
        RECT 1359.920 90.200 1360.610 90.340 ;
        RECT 1359.920 90.060 1360.060 90.200 ;
        RECT 1360.290 90.140 1360.610 90.200 ;
        RECT 1359.830 89.800 1360.150 90.060 ;
        RECT 419.130 33.900 419.450 33.960 ;
        RECT 1359.370 33.900 1359.690 33.960 ;
        RECT 419.130 33.760 1359.690 33.900 ;
        RECT 419.130 33.700 419.450 33.760 ;
        RECT 1359.370 33.700 1359.690 33.760 ;
      LAYER via ;
        RECT 1360.320 1365.820 1360.580 1366.080 ;
        RECT 1360.320 1365.140 1360.580 1365.400 ;
        RECT 1360.320 1303.940 1360.580 1304.200 ;
        RECT 1360.320 1256.000 1360.580 1256.260 ;
        RECT 1359.400 1159.100 1359.660 1159.360 ;
        RECT 1360.320 1159.100 1360.580 1159.360 ;
        RECT 1359.400 1062.540 1359.660 1062.800 ;
        RECT 1360.320 1062.540 1360.580 1062.800 ;
        RECT 1360.320 931.980 1360.580 932.240 ;
        RECT 1359.860 917.700 1360.120 917.960 ;
        RECT 1359.860 869.420 1360.120 869.680 ;
        RECT 1360.320 869.420 1360.580 869.680 ;
        RECT 1360.320 862.280 1360.580 862.540 ;
        RECT 1359.860 814.340 1360.120 814.600 ;
        RECT 1359.860 789.860 1360.120 790.120 ;
        RECT 1359.860 742.940 1360.120 743.200 ;
        RECT 1359.860 724.240 1360.120 724.500 ;
        RECT 1360.320 724.240 1360.580 724.500 ;
        RECT 1359.400 675.960 1359.660 676.220 ;
        RECT 1359.860 675.960 1360.120 676.220 ;
        RECT 1359.860 627.680 1360.120 627.940 ;
        RECT 1360.320 627.680 1360.580 627.940 ;
        RECT 1359.860 620.540 1360.120 620.800 ;
        RECT 1359.860 576.680 1360.120 576.940 ;
        RECT 1359.400 524.320 1359.660 524.580 ;
        RECT 1359.860 524.320 1360.120 524.580 ;
        RECT 1359.400 496.440 1359.660 496.700 ;
        RECT 1360.320 496.440 1360.580 496.700 ;
        RECT 1360.320 421.300 1360.580 421.560 ;
        RECT 1359.860 420.960 1360.120 421.220 ;
        RECT 1359.860 413.820 1360.120 414.080 ;
        RECT 1359.860 365.880 1360.120 366.140 ;
        RECT 1359.860 324.060 1360.120 324.320 ;
        RECT 1360.320 324.060 1360.580 324.320 ;
        RECT 1360.320 258.780 1360.580 259.040 ;
        RECT 1359.860 234.640 1360.120 234.900 ;
        RECT 1359.860 214.580 1360.120 214.840 ;
        RECT 1360.320 144.880 1360.580 145.140 ;
        RECT 1360.320 90.140 1360.580 90.400 ;
        RECT 1359.860 89.800 1360.120 90.060 ;
        RECT 419.160 33.700 419.420 33.960 ;
        RECT 1359.400 33.700 1359.660 33.960 ;
      LAYER met2 ;
        RECT 1363.920 1700.410 1364.200 1704.000 ;
        RECT 1362.220 1700.270 1364.200 1700.410 ;
        RECT 1362.220 1678.650 1362.360 1700.270 ;
        RECT 1363.920 1700.000 1364.200 1700.270 ;
        RECT 1360.380 1678.510 1362.360 1678.650 ;
        RECT 1360.380 1607.930 1360.520 1678.510 ;
        RECT 1359.920 1607.790 1360.520 1607.930 ;
        RECT 1359.920 1607.250 1360.060 1607.790 ;
        RECT 1359.920 1607.110 1360.520 1607.250 ;
        RECT 1360.380 1463.090 1360.520 1607.110 ;
        RECT 1359.920 1462.950 1360.520 1463.090 ;
        RECT 1359.920 1462.410 1360.060 1462.950 ;
        RECT 1359.920 1462.270 1360.520 1462.410 ;
        RECT 1360.380 1366.110 1360.520 1462.270 ;
        RECT 1360.320 1365.790 1360.580 1366.110 ;
        RECT 1360.320 1365.110 1360.580 1365.430 ;
        RECT 1360.380 1304.230 1360.520 1365.110 ;
        RECT 1360.320 1303.910 1360.580 1304.230 ;
        RECT 1360.320 1255.970 1360.580 1256.290 ;
        RECT 1360.380 1207.525 1360.520 1255.970 ;
        RECT 1359.390 1207.155 1359.670 1207.525 ;
        RECT 1360.310 1207.155 1360.590 1207.525 ;
        RECT 1359.460 1159.390 1359.600 1207.155 ;
        RECT 1359.400 1159.070 1359.660 1159.390 ;
        RECT 1360.320 1159.070 1360.580 1159.390 ;
        RECT 1360.380 1110.965 1360.520 1159.070 ;
        RECT 1359.390 1110.595 1359.670 1110.965 ;
        RECT 1360.310 1110.595 1360.590 1110.965 ;
        RECT 1359.460 1062.830 1359.600 1110.595 ;
        RECT 1359.400 1062.510 1359.660 1062.830 ;
        RECT 1360.320 1062.510 1360.580 1062.830 ;
        RECT 1360.380 980.290 1360.520 1062.510 ;
        RECT 1359.920 980.150 1360.520 980.290 ;
        RECT 1359.920 979.610 1360.060 980.150 ;
        RECT 1359.920 979.470 1360.520 979.610 ;
        RECT 1360.380 932.270 1360.520 979.470 ;
        RECT 1360.320 931.950 1360.580 932.270 ;
        RECT 1359.860 917.670 1360.120 917.990 ;
        RECT 1359.920 869.710 1360.060 917.670 ;
        RECT 1359.860 869.390 1360.120 869.710 ;
        RECT 1360.320 869.390 1360.580 869.710 ;
        RECT 1360.380 862.570 1360.520 869.390 ;
        RECT 1360.320 862.250 1360.580 862.570 ;
        RECT 1359.860 814.310 1360.120 814.630 ;
        RECT 1359.920 790.150 1360.060 814.310 ;
        RECT 1359.860 789.830 1360.120 790.150 ;
        RECT 1359.860 742.910 1360.120 743.230 ;
        RECT 1359.920 724.530 1360.060 742.910 ;
        RECT 1359.860 724.210 1360.120 724.530 ;
        RECT 1360.320 724.210 1360.580 724.530 ;
        RECT 1360.380 699.450 1360.520 724.210 ;
        RECT 1359.920 699.310 1360.520 699.450 ;
        RECT 1359.920 676.250 1360.060 699.310 ;
        RECT 1359.400 675.930 1359.660 676.250 ;
        RECT 1359.860 675.930 1360.120 676.250 ;
        RECT 1359.460 628.165 1359.600 675.930 ;
        RECT 1359.390 627.795 1359.670 628.165 ;
        RECT 1359.860 627.650 1360.120 627.970 ;
        RECT 1360.310 627.795 1360.590 628.165 ;
        RECT 1360.320 627.650 1360.580 627.795 ;
        RECT 1359.920 620.830 1360.060 627.650 ;
        RECT 1359.860 620.510 1360.120 620.830 ;
        RECT 1359.860 576.650 1360.120 576.970 ;
        RECT 1359.920 524.610 1360.060 576.650 ;
        RECT 1359.400 524.290 1359.660 524.610 ;
        RECT 1359.860 524.290 1360.120 524.610 ;
        RECT 1359.460 496.730 1359.600 524.290 ;
        RECT 1359.400 496.410 1359.660 496.730 ;
        RECT 1360.320 496.410 1360.580 496.730 ;
        RECT 1360.380 421.590 1360.520 496.410 ;
        RECT 1360.320 421.270 1360.580 421.590 ;
        RECT 1359.860 420.930 1360.120 421.250 ;
        RECT 1359.920 414.110 1360.060 420.930 ;
        RECT 1359.860 413.790 1360.120 414.110 ;
        RECT 1359.860 365.850 1360.120 366.170 ;
        RECT 1359.920 324.350 1360.060 365.850 ;
        RECT 1359.860 324.030 1360.120 324.350 ;
        RECT 1360.320 324.030 1360.580 324.350 ;
        RECT 1360.380 259.070 1360.520 324.030 ;
        RECT 1360.320 258.750 1360.580 259.070 ;
        RECT 1359.860 234.610 1360.120 234.930 ;
        RECT 1359.920 214.870 1360.060 234.610 ;
        RECT 1359.860 214.550 1360.120 214.870 ;
        RECT 1360.320 144.850 1360.580 145.170 ;
        RECT 1360.380 90.430 1360.520 144.850 ;
        RECT 1360.320 90.110 1360.580 90.430 ;
        RECT 1359.860 89.770 1360.120 90.090 ;
        RECT 1359.920 65.690 1360.060 89.770 ;
        RECT 1359.000 65.550 1360.060 65.690 ;
        RECT 1359.000 61.610 1359.140 65.550 ;
        RECT 1359.000 61.470 1359.600 61.610 ;
        RECT 1359.460 33.990 1359.600 61.470 ;
        RECT 419.160 33.670 419.420 33.990 ;
        RECT 1359.400 33.670 1359.660 33.990 ;
        RECT 419.220 2.400 419.360 33.670 ;
        RECT 419.010 -4.800 419.570 2.400 ;
      LAYER via2 ;
        RECT 1359.390 1207.200 1359.670 1207.480 ;
        RECT 1360.310 1207.200 1360.590 1207.480 ;
        RECT 1359.390 1110.640 1359.670 1110.920 ;
        RECT 1360.310 1110.640 1360.590 1110.920 ;
        RECT 1359.390 627.840 1359.670 628.120 ;
        RECT 1360.310 627.840 1360.590 628.120 ;
      LAYER met3 ;
        RECT 1359.365 1207.490 1359.695 1207.505 ;
        RECT 1360.285 1207.490 1360.615 1207.505 ;
        RECT 1359.365 1207.190 1360.615 1207.490 ;
        RECT 1359.365 1207.175 1359.695 1207.190 ;
        RECT 1360.285 1207.175 1360.615 1207.190 ;
        RECT 1359.365 1110.930 1359.695 1110.945 ;
        RECT 1360.285 1110.930 1360.615 1110.945 ;
        RECT 1359.365 1110.630 1360.615 1110.930 ;
        RECT 1359.365 1110.615 1359.695 1110.630 ;
        RECT 1360.285 1110.615 1360.615 1110.630 ;
        RECT 1359.365 628.130 1359.695 628.145 ;
        RECT 1360.285 628.130 1360.615 628.145 ;
        RECT 1359.365 627.830 1360.615 628.130 ;
        RECT 1359.365 627.815 1359.695 627.830 ;
        RECT 1360.285 627.815 1360.615 627.830 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 436.610 37.640 436.930 37.700 ;
        RECT 1373.170 37.640 1373.490 37.700 ;
        RECT 436.610 37.500 1373.490 37.640 ;
        RECT 436.610 37.440 436.930 37.500 ;
        RECT 1373.170 37.440 1373.490 37.500 ;
      LAYER via ;
        RECT 436.640 37.440 436.900 37.700 ;
        RECT 1373.200 37.440 1373.460 37.700 ;
      LAYER met2 ;
        RECT 1373.120 1700.000 1373.400 1704.000 ;
        RECT 1373.260 37.730 1373.400 1700.000 ;
        RECT 436.640 37.410 436.900 37.730 ;
        RECT 1373.200 37.410 1373.460 37.730 ;
        RECT 436.700 2.400 436.840 37.410 ;
        RECT 436.490 -4.800 437.050 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 454.550 37.300 454.870 37.360 ;
        RECT 1380.070 37.300 1380.390 37.360 ;
        RECT 454.550 37.160 1380.390 37.300 ;
        RECT 454.550 37.100 454.870 37.160 ;
        RECT 1380.070 37.100 1380.390 37.160 ;
      LAYER via ;
        RECT 454.580 37.100 454.840 37.360 ;
        RECT 1380.100 37.100 1380.360 37.360 ;
      LAYER met2 ;
        RECT 1382.320 1700.410 1382.600 1704.000 ;
        RECT 1380.160 1700.270 1382.600 1700.410 ;
        RECT 1380.160 37.390 1380.300 1700.270 ;
        RECT 1382.320 1700.000 1382.600 1700.270 ;
        RECT 454.580 37.070 454.840 37.390 ;
        RECT 1380.100 37.070 1380.360 37.390 ;
        RECT 454.640 2.400 454.780 37.070 ;
        RECT 454.430 -4.800 454.990 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1387.965 1545.045 1388.135 1559.835 ;
        RECT 1387.965 1490.985 1388.135 1538.755 ;
        RECT 1387.965 1400.885 1388.135 1490.475 ;
      LAYER mcon ;
        RECT 1387.965 1559.665 1388.135 1559.835 ;
        RECT 1387.965 1538.585 1388.135 1538.755 ;
        RECT 1387.965 1490.305 1388.135 1490.475 ;
      LAYER met1 ;
        RECT 1386.510 1617.960 1386.830 1618.020 ;
        RECT 1387.890 1617.960 1388.210 1618.020 ;
        RECT 1386.510 1617.820 1388.210 1617.960 ;
        RECT 1386.510 1617.760 1386.830 1617.820 ;
        RECT 1387.890 1617.760 1388.210 1617.820 ;
        RECT 1387.890 1559.820 1388.210 1559.880 ;
        RECT 1387.695 1559.680 1388.210 1559.820 ;
        RECT 1387.890 1559.620 1388.210 1559.680 ;
        RECT 1387.430 1545.200 1387.750 1545.260 ;
        RECT 1387.905 1545.200 1388.195 1545.245 ;
        RECT 1387.430 1545.060 1388.195 1545.200 ;
        RECT 1387.430 1545.000 1387.750 1545.060 ;
        RECT 1387.905 1545.015 1388.195 1545.060 ;
        RECT 1387.890 1538.740 1388.210 1538.800 ;
        RECT 1387.695 1538.600 1388.210 1538.740 ;
        RECT 1387.890 1538.540 1388.210 1538.600 ;
        RECT 1387.890 1491.140 1388.210 1491.200 ;
        RECT 1387.695 1491.000 1388.210 1491.140 ;
        RECT 1387.890 1490.940 1388.210 1491.000 ;
        RECT 1387.890 1490.460 1388.210 1490.520 ;
        RECT 1387.695 1490.320 1388.210 1490.460 ;
        RECT 1387.890 1490.260 1388.210 1490.320 ;
        RECT 1387.905 1401.040 1388.195 1401.085 ;
        RECT 1388.350 1401.040 1388.670 1401.100 ;
        RECT 1387.905 1400.900 1388.670 1401.040 ;
        RECT 1387.905 1400.855 1388.195 1400.900 ;
        RECT 1388.350 1400.840 1388.670 1400.900 ;
        RECT 1387.890 1304.140 1388.210 1304.200 ;
        RECT 1388.350 1304.140 1388.670 1304.200 ;
        RECT 1387.890 1304.000 1388.670 1304.140 ;
        RECT 1387.890 1303.940 1388.210 1304.000 ;
        RECT 1388.350 1303.940 1388.670 1304.000 ;
        RECT 1387.890 1159.300 1388.210 1159.360 ;
        RECT 1388.350 1159.300 1388.670 1159.360 ;
        RECT 1387.890 1159.160 1388.670 1159.300 ;
        RECT 1387.890 1159.100 1388.210 1159.160 ;
        RECT 1388.350 1159.100 1388.670 1159.160 ;
        RECT 1387.890 1062.740 1388.210 1062.800 ;
        RECT 1388.350 1062.740 1388.670 1062.800 ;
        RECT 1387.890 1062.600 1388.670 1062.740 ;
        RECT 1387.890 1062.540 1388.210 1062.600 ;
        RECT 1388.350 1062.540 1388.670 1062.600 ;
        RECT 1387.430 979.780 1387.750 979.840 ;
        RECT 1388.350 979.780 1388.670 979.840 ;
        RECT 1387.430 979.640 1388.670 979.780 ;
        RECT 1387.430 979.580 1387.750 979.640 ;
        RECT 1388.350 979.580 1388.670 979.640 ;
        RECT 1388.350 931.980 1388.670 932.240 ;
        RECT 1388.440 931.220 1388.580 931.980 ;
        RECT 1388.350 930.960 1388.670 931.220 ;
        RECT 1388.350 690.440 1388.670 690.500 ;
        RECT 1387.980 690.300 1388.670 690.440 ;
        RECT 1387.980 689.820 1388.120 690.300 ;
        RECT 1388.350 690.240 1388.670 690.300 ;
        RECT 1387.890 689.560 1388.210 689.820 ;
        RECT 1387.430 579.600 1387.750 579.660 ;
        RECT 1388.350 579.600 1388.670 579.660 ;
        RECT 1387.430 579.460 1388.670 579.600 ;
        RECT 1387.430 579.400 1387.750 579.460 ;
        RECT 1388.350 579.400 1388.670 579.460 ;
        RECT 1387.890 497.120 1388.210 497.380 ;
        RECT 1387.980 496.700 1388.120 497.120 ;
        RECT 1387.890 496.440 1388.210 496.700 ;
        RECT 1387.890 352.280 1388.210 352.540 ;
        RECT 1387.980 351.860 1388.120 352.280 ;
        RECT 1387.890 351.600 1388.210 351.860 ;
        RECT 1387.890 110.740 1388.210 110.800 ;
        RECT 1387.520 110.600 1388.210 110.740 ;
        RECT 1387.520 110.460 1387.660 110.600 ;
        RECT 1387.890 110.540 1388.210 110.600 ;
        RECT 1387.430 110.200 1387.750 110.460 ;
        RECT 472.490 36.960 472.810 37.020 ;
        RECT 1387.430 36.960 1387.750 37.020 ;
        RECT 472.490 36.820 1387.750 36.960 ;
        RECT 472.490 36.760 472.810 36.820 ;
        RECT 1387.430 36.760 1387.750 36.820 ;
      LAYER via ;
        RECT 1386.540 1617.760 1386.800 1618.020 ;
        RECT 1387.920 1617.760 1388.180 1618.020 ;
        RECT 1387.920 1559.620 1388.180 1559.880 ;
        RECT 1387.460 1545.000 1387.720 1545.260 ;
        RECT 1387.920 1538.540 1388.180 1538.800 ;
        RECT 1387.920 1490.940 1388.180 1491.200 ;
        RECT 1387.920 1490.260 1388.180 1490.520 ;
        RECT 1388.380 1400.840 1388.640 1401.100 ;
        RECT 1387.920 1303.940 1388.180 1304.200 ;
        RECT 1388.380 1303.940 1388.640 1304.200 ;
        RECT 1387.920 1159.100 1388.180 1159.360 ;
        RECT 1388.380 1159.100 1388.640 1159.360 ;
        RECT 1387.920 1062.540 1388.180 1062.800 ;
        RECT 1388.380 1062.540 1388.640 1062.800 ;
        RECT 1387.460 979.580 1387.720 979.840 ;
        RECT 1388.380 979.580 1388.640 979.840 ;
        RECT 1388.380 931.980 1388.640 932.240 ;
        RECT 1388.380 930.960 1388.640 931.220 ;
        RECT 1388.380 690.240 1388.640 690.500 ;
        RECT 1387.920 689.560 1388.180 689.820 ;
        RECT 1387.460 579.400 1387.720 579.660 ;
        RECT 1388.380 579.400 1388.640 579.660 ;
        RECT 1387.920 497.120 1388.180 497.380 ;
        RECT 1387.920 496.440 1388.180 496.700 ;
        RECT 1387.920 352.280 1388.180 352.540 ;
        RECT 1387.920 351.600 1388.180 351.860 ;
        RECT 1387.920 110.540 1388.180 110.800 ;
        RECT 1387.460 110.200 1387.720 110.460 ;
        RECT 472.520 36.760 472.780 37.020 ;
        RECT 1387.460 36.760 1387.720 37.020 ;
      LAYER met2 ;
        RECT 1391.520 1700.410 1391.800 1704.000 ;
        RECT 1389.820 1700.270 1391.800 1700.410 ;
        RECT 1389.820 1678.650 1389.960 1700.270 ;
        RECT 1391.520 1700.000 1391.800 1700.270 ;
        RECT 1387.980 1678.510 1389.960 1678.650 ;
        RECT 1387.980 1618.050 1388.120 1678.510 ;
        RECT 1386.540 1617.730 1386.800 1618.050 ;
        RECT 1387.920 1617.730 1388.180 1618.050 ;
        RECT 1386.600 1594.445 1386.740 1617.730 ;
        RECT 1386.530 1594.075 1386.810 1594.445 ;
        RECT 1387.910 1594.075 1388.190 1594.445 ;
        RECT 1387.980 1559.910 1388.120 1594.075 ;
        RECT 1387.920 1559.590 1388.180 1559.910 ;
        RECT 1387.460 1544.970 1387.720 1545.290 ;
        RECT 1387.520 1539.250 1387.660 1544.970 ;
        RECT 1387.520 1539.110 1388.120 1539.250 ;
        RECT 1387.980 1538.830 1388.120 1539.110 ;
        RECT 1387.920 1538.510 1388.180 1538.830 ;
        RECT 1387.920 1490.910 1388.180 1491.230 ;
        RECT 1387.980 1490.550 1388.120 1490.910 ;
        RECT 1387.920 1490.230 1388.180 1490.550 ;
        RECT 1388.380 1400.810 1388.640 1401.130 ;
        RECT 1388.440 1352.365 1388.580 1400.810 ;
        RECT 1388.370 1351.995 1388.650 1352.365 ;
        RECT 1388.830 1351.315 1389.110 1351.685 ;
        RECT 1388.900 1304.650 1389.040 1351.315 ;
        RECT 1387.980 1304.510 1389.040 1304.650 ;
        RECT 1387.980 1304.230 1388.120 1304.510 ;
        RECT 1387.920 1303.910 1388.180 1304.230 ;
        RECT 1388.380 1303.910 1388.640 1304.230 ;
        RECT 1388.440 1221.010 1388.580 1303.910 ;
        RECT 1387.980 1220.870 1388.580 1221.010 ;
        RECT 1387.980 1159.390 1388.120 1220.870 ;
        RECT 1387.920 1159.070 1388.180 1159.390 ;
        RECT 1388.380 1159.070 1388.640 1159.390 ;
        RECT 1388.440 1124.450 1388.580 1159.070 ;
        RECT 1387.980 1124.310 1388.580 1124.450 ;
        RECT 1387.980 1062.830 1388.120 1124.310 ;
        RECT 1387.920 1062.510 1388.180 1062.830 ;
        RECT 1388.380 1062.510 1388.640 1062.830 ;
        RECT 1388.440 1027.890 1388.580 1062.510 ;
        RECT 1387.980 1027.750 1388.580 1027.890 ;
        RECT 1387.980 980.290 1388.120 1027.750 ;
        RECT 1387.520 980.150 1388.120 980.290 ;
        RECT 1387.520 979.870 1387.660 980.150 ;
        RECT 1387.460 979.550 1387.720 979.870 ;
        RECT 1388.380 979.550 1388.640 979.870 ;
        RECT 1388.440 932.270 1388.580 979.550 ;
        RECT 1388.380 931.950 1388.640 932.270 ;
        RECT 1388.380 930.930 1388.640 931.250 ;
        RECT 1388.440 917.730 1388.580 930.930 ;
        RECT 1387.980 917.590 1388.580 917.730 ;
        RECT 1387.980 835.450 1388.120 917.590 ;
        RECT 1387.520 835.310 1388.120 835.450 ;
        RECT 1387.520 834.770 1387.660 835.310 ;
        RECT 1387.520 834.630 1388.120 834.770 ;
        RECT 1387.980 738.890 1388.120 834.630 ;
        RECT 1387.520 738.750 1388.120 738.890 ;
        RECT 1387.520 738.210 1387.660 738.750 ;
        RECT 1387.520 738.070 1388.580 738.210 ;
        RECT 1388.440 690.530 1388.580 738.070 ;
        RECT 1388.380 690.210 1388.640 690.530 ;
        RECT 1387.920 689.530 1388.180 689.850 ;
        RECT 1387.980 580.565 1388.120 689.530 ;
        RECT 1387.910 580.195 1388.190 580.565 ;
        RECT 1387.450 579.515 1387.730 579.885 ;
        RECT 1387.460 579.370 1387.720 579.515 ;
        RECT 1388.380 579.370 1388.640 579.690 ;
        RECT 1388.440 554.610 1388.580 579.370 ;
        RECT 1387.980 554.470 1388.580 554.610 ;
        RECT 1387.980 497.410 1388.120 554.470 ;
        RECT 1387.920 497.090 1388.180 497.410 ;
        RECT 1387.920 496.410 1388.180 496.730 ;
        RECT 1387.980 352.570 1388.120 496.410 ;
        RECT 1387.920 352.250 1388.180 352.570 ;
        RECT 1387.920 351.570 1388.180 351.890 ;
        RECT 1387.980 258.810 1388.120 351.570 ;
        RECT 1387.980 258.670 1388.580 258.810 ;
        RECT 1388.440 145.250 1388.580 258.670 ;
        RECT 1387.980 145.110 1388.580 145.250 ;
        RECT 1387.980 110.830 1388.120 145.110 ;
        RECT 1387.920 110.510 1388.180 110.830 ;
        RECT 1387.460 110.170 1387.720 110.490 ;
        RECT 1387.520 37.050 1387.660 110.170 ;
        RECT 472.520 36.730 472.780 37.050 ;
        RECT 1387.460 36.730 1387.720 37.050 ;
        RECT 472.580 2.400 472.720 36.730 ;
        RECT 472.370 -4.800 472.930 2.400 ;
      LAYER via2 ;
        RECT 1386.530 1594.120 1386.810 1594.400 ;
        RECT 1387.910 1594.120 1388.190 1594.400 ;
        RECT 1388.370 1352.040 1388.650 1352.320 ;
        RECT 1388.830 1351.360 1389.110 1351.640 ;
        RECT 1387.910 580.240 1388.190 580.520 ;
        RECT 1387.450 579.560 1387.730 579.840 ;
      LAYER met3 ;
        RECT 1386.505 1594.410 1386.835 1594.425 ;
        RECT 1387.885 1594.410 1388.215 1594.425 ;
        RECT 1386.505 1594.110 1388.215 1594.410 ;
        RECT 1386.505 1594.095 1386.835 1594.110 ;
        RECT 1387.885 1594.095 1388.215 1594.110 ;
        RECT 1388.345 1352.330 1388.675 1352.345 ;
        RECT 1387.670 1352.030 1388.675 1352.330 ;
        RECT 1387.670 1351.650 1387.970 1352.030 ;
        RECT 1388.345 1352.015 1388.675 1352.030 ;
        RECT 1388.805 1351.650 1389.135 1351.665 ;
        RECT 1387.670 1351.350 1389.135 1351.650 ;
        RECT 1388.805 1351.335 1389.135 1351.350 ;
        RECT 1387.885 580.530 1388.215 580.545 ;
        RECT 1387.670 580.215 1388.215 580.530 ;
        RECT 1387.670 579.865 1387.970 580.215 ;
        RECT 1387.425 579.550 1387.970 579.865 ;
        RECT 1387.425 579.535 1387.755 579.550 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 495.950 51.920 496.270 51.980 ;
        RECT 1400.770 51.920 1401.090 51.980 ;
        RECT 495.950 51.780 1401.090 51.920 ;
        RECT 495.950 51.720 496.270 51.780 ;
        RECT 1400.770 51.720 1401.090 51.780 ;
        RECT 490.430 15.540 490.750 15.600 ;
        RECT 495.950 15.540 496.270 15.600 ;
        RECT 490.430 15.400 496.270 15.540 ;
        RECT 490.430 15.340 490.750 15.400 ;
        RECT 495.950 15.340 496.270 15.400 ;
      LAYER via ;
        RECT 495.980 51.720 496.240 51.980 ;
        RECT 1400.800 51.720 1401.060 51.980 ;
        RECT 490.460 15.340 490.720 15.600 ;
        RECT 495.980 15.340 496.240 15.600 ;
      LAYER met2 ;
        RECT 1400.720 1700.000 1401.000 1704.000 ;
        RECT 1400.860 52.010 1401.000 1700.000 ;
        RECT 495.980 51.690 496.240 52.010 ;
        RECT 1400.800 51.690 1401.060 52.010 ;
        RECT 496.040 15.630 496.180 51.690 ;
        RECT 490.460 15.310 490.720 15.630 ;
        RECT 495.980 15.310 496.240 15.630 ;
        RECT 490.520 2.400 490.660 15.310 ;
        RECT 490.310 -4.800 490.870 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 507.910 52.260 508.230 52.320 ;
        RECT 1407.670 52.260 1407.990 52.320 ;
        RECT 507.910 52.120 1407.990 52.260 ;
        RECT 507.910 52.060 508.230 52.120 ;
        RECT 1407.670 52.060 1407.990 52.120 ;
      LAYER via ;
        RECT 507.940 52.060 508.200 52.320 ;
        RECT 1407.700 52.060 1407.960 52.320 ;
      LAYER met2 ;
        RECT 1409.920 1700.410 1410.200 1704.000 ;
        RECT 1407.760 1700.270 1410.200 1700.410 ;
        RECT 1407.760 52.350 1407.900 1700.270 ;
        RECT 1409.920 1700.000 1410.200 1700.270 ;
        RECT 507.940 52.030 508.200 52.350 ;
        RECT 1407.700 52.030 1407.960 52.350 ;
        RECT 508.000 2.400 508.140 52.030 ;
        RECT 507.790 -4.800 508.350 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1415.105 1538.925 1415.275 1587.035 ;
        RECT 1415.565 1449.165 1415.735 1497.275 ;
        RECT 1415.105 662.405 1415.275 710.515 ;
        RECT 1414.645 476.085 1414.815 524.195 ;
        RECT 1415.565 282.965 1415.735 331.075 ;
        RECT 1414.645 179.605 1414.815 227.715 ;
      LAYER mcon ;
        RECT 1415.105 1586.865 1415.275 1587.035 ;
        RECT 1415.565 1497.105 1415.735 1497.275 ;
        RECT 1415.105 710.345 1415.275 710.515 ;
        RECT 1414.645 524.025 1414.815 524.195 ;
        RECT 1415.565 330.905 1415.735 331.075 ;
        RECT 1414.645 227.545 1414.815 227.715 ;
      LAYER met1 ;
        RECT 1415.030 1593.820 1415.350 1593.880 ;
        RECT 1415.490 1593.820 1415.810 1593.880 ;
        RECT 1415.030 1593.680 1415.810 1593.820 ;
        RECT 1415.030 1593.620 1415.350 1593.680 ;
        RECT 1415.490 1593.620 1415.810 1593.680 ;
        RECT 1415.030 1587.020 1415.350 1587.080 ;
        RECT 1414.835 1586.880 1415.350 1587.020 ;
        RECT 1415.030 1586.820 1415.350 1586.880 ;
        RECT 1415.030 1539.080 1415.350 1539.140 ;
        RECT 1414.835 1538.940 1415.350 1539.080 ;
        RECT 1415.030 1538.880 1415.350 1538.940 ;
        RECT 1415.030 1511.340 1415.350 1511.600 ;
        RECT 1415.120 1510.520 1415.260 1511.340 ;
        RECT 1415.490 1510.520 1415.810 1510.580 ;
        RECT 1415.120 1510.380 1415.810 1510.520 ;
        RECT 1415.490 1510.320 1415.810 1510.380 ;
        RECT 1415.490 1497.260 1415.810 1497.320 ;
        RECT 1415.295 1497.120 1415.810 1497.260 ;
        RECT 1415.490 1497.060 1415.810 1497.120 ;
        RECT 1415.490 1449.320 1415.810 1449.380 ;
        RECT 1415.295 1449.180 1415.810 1449.320 ;
        RECT 1415.490 1449.120 1415.810 1449.180 ;
        RECT 1415.490 1365.820 1415.810 1366.080 ;
        RECT 1415.580 1365.400 1415.720 1365.820 ;
        RECT 1415.490 1365.140 1415.810 1365.400 ;
        RECT 1415.490 1269.260 1415.810 1269.520 ;
        RECT 1415.580 1268.840 1415.720 1269.260 ;
        RECT 1415.490 1268.580 1415.810 1268.840 ;
        RECT 1415.490 1076.140 1415.810 1076.400 ;
        RECT 1415.580 1075.720 1415.720 1076.140 ;
        RECT 1415.490 1075.460 1415.810 1075.720 ;
        RECT 1415.490 724.780 1415.810 724.840 ;
        RECT 1415.120 724.640 1415.810 724.780 ;
        RECT 1415.120 724.500 1415.260 724.640 ;
        RECT 1415.490 724.580 1415.810 724.640 ;
        RECT 1415.030 724.240 1415.350 724.500 ;
        RECT 1415.030 710.500 1415.350 710.560 ;
        RECT 1414.835 710.360 1415.350 710.500 ;
        RECT 1415.030 710.300 1415.350 710.360 ;
        RECT 1415.045 662.560 1415.335 662.605 ;
        RECT 1415.490 662.560 1415.810 662.620 ;
        RECT 1415.045 662.420 1415.810 662.560 ;
        RECT 1415.045 662.375 1415.335 662.420 ;
        RECT 1415.490 662.360 1415.810 662.420 ;
        RECT 1415.490 572.800 1415.810 572.860 ;
        RECT 1415.950 572.800 1416.270 572.860 ;
        RECT 1415.490 572.660 1416.270 572.800 ;
        RECT 1415.490 572.600 1415.810 572.660 ;
        RECT 1415.950 572.600 1416.270 572.660 ;
        RECT 1414.570 548.660 1414.890 548.720 ;
        RECT 1415.490 548.660 1415.810 548.720 ;
        RECT 1414.570 548.520 1415.810 548.660 ;
        RECT 1414.570 548.460 1414.890 548.520 ;
        RECT 1415.490 548.460 1415.810 548.520 ;
        RECT 1414.570 524.180 1414.890 524.240 ;
        RECT 1414.375 524.040 1414.890 524.180 ;
        RECT 1414.570 523.980 1414.890 524.040 ;
        RECT 1414.570 476.240 1414.890 476.300 ;
        RECT 1414.375 476.100 1414.890 476.240 ;
        RECT 1414.570 476.040 1414.890 476.100 ;
        RECT 1415.950 331.740 1416.270 331.800 ;
        RECT 1415.580 331.600 1416.270 331.740 ;
        RECT 1415.580 331.105 1415.720 331.600 ;
        RECT 1415.950 331.540 1416.270 331.600 ;
        RECT 1415.505 330.875 1415.795 331.105 ;
        RECT 1415.490 283.120 1415.810 283.180 ;
        RECT 1415.295 282.980 1415.810 283.120 ;
        RECT 1415.490 282.920 1415.810 282.980 ;
        RECT 1414.585 227.700 1414.875 227.745 ;
        RECT 1415.950 227.700 1416.270 227.760 ;
        RECT 1414.585 227.560 1416.270 227.700 ;
        RECT 1414.585 227.515 1414.875 227.560 ;
        RECT 1415.950 227.500 1416.270 227.560 ;
        RECT 1414.570 179.760 1414.890 179.820 ;
        RECT 1414.375 179.620 1414.890 179.760 ;
        RECT 1414.570 179.560 1414.890 179.620 ;
        RECT 525.850 52.940 526.170 53.000 ;
        RECT 1415.030 52.940 1415.350 53.000 ;
        RECT 525.850 52.800 1415.350 52.940 ;
        RECT 525.850 52.740 526.170 52.800 ;
        RECT 1415.030 52.740 1415.350 52.800 ;
      LAYER via ;
        RECT 1415.060 1593.620 1415.320 1593.880 ;
        RECT 1415.520 1593.620 1415.780 1593.880 ;
        RECT 1415.060 1586.820 1415.320 1587.080 ;
        RECT 1415.060 1538.880 1415.320 1539.140 ;
        RECT 1415.060 1511.340 1415.320 1511.600 ;
        RECT 1415.520 1510.320 1415.780 1510.580 ;
        RECT 1415.520 1497.060 1415.780 1497.320 ;
        RECT 1415.520 1449.120 1415.780 1449.380 ;
        RECT 1415.520 1365.820 1415.780 1366.080 ;
        RECT 1415.520 1365.140 1415.780 1365.400 ;
        RECT 1415.520 1269.260 1415.780 1269.520 ;
        RECT 1415.520 1268.580 1415.780 1268.840 ;
        RECT 1415.520 1076.140 1415.780 1076.400 ;
        RECT 1415.520 1075.460 1415.780 1075.720 ;
        RECT 1415.520 724.580 1415.780 724.840 ;
        RECT 1415.060 724.240 1415.320 724.500 ;
        RECT 1415.060 710.300 1415.320 710.560 ;
        RECT 1415.520 662.360 1415.780 662.620 ;
        RECT 1415.520 572.600 1415.780 572.860 ;
        RECT 1415.980 572.600 1416.240 572.860 ;
        RECT 1414.600 548.460 1414.860 548.720 ;
        RECT 1415.520 548.460 1415.780 548.720 ;
        RECT 1414.600 523.980 1414.860 524.240 ;
        RECT 1414.600 476.040 1414.860 476.300 ;
        RECT 1415.980 331.540 1416.240 331.800 ;
        RECT 1415.520 282.920 1415.780 283.180 ;
        RECT 1415.980 227.500 1416.240 227.760 ;
        RECT 1414.600 179.560 1414.860 179.820 ;
        RECT 525.880 52.740 526.140 53.000 ;
        RECT 1415.060 52.740 1415.320 53.000 ;
      LAYER met2 ;
        RECT 1419.120 1701.090 1419.400 1704.000 ;
        RECT 1416.500 1700.950 1419.400 1701.090 ;
        RECT 1416.500 1677.970 1416.640 1700.950 ;
        RECT 1419.120 1700.000 1419.400 1700.950 ;
        RECT 1415.580 1677.830 1416.640 1677.970 ;
        RECT 1415.580 1593.910 1415.720 1677.830 ;
        RECT 1415.060 1593.590 1415.320 1593.910 ;
        RECT 1415.520 1593.590 1415.780 1593.910 ;
        RECT 1415.120 1587.110 1415.260 1593.590 ;
        RECT 1415.060 1586.790 1415.320 1587.110 ;
        RECT 1415.060 1538.850 1415.320 1539.170 ;
        RECT 1415.120 1511.630 1415.260 1538.850 ;
        RECT 1415.060 1511.310 1415.320 1511.630 ;
        RECT 1415.520 1510.290 1415.780 1510.610 ;
        RECT 1415.580 1497.350 1415.720 1510.290 ;
        RECT 1415.520 1497.030 1415.780 1497.350 ;
        RECT 1415.520 1449.090 1415.780 1449.410 ;
        RECT 1415.580 1366.110 1415.720 1449.090 ;
        RECT 1415.520 1365.790 1415.780 1366.110 ;
        RECT 1415.520 1365.110 1415.780 1365.430 ;
        RECT 1415.580 1269.550 1415.720 1365.110 ;
        RECT 1415.520 1269.230 1415.780 1269.550 ;
        RECT 1415.520 1268.550 1415.780 1268.870 ;
        RECT 1415.580 1173.410 1415.720 1268.550 ;
        RECT 1415.120 1173.270 1415.720 1173.410 ;
        RECT 1415.120 1172.730 1415.260 1173.270 ;
        RECT 1415.120 1172.590 1415.720 1172.730 ;
        RECT 1415.580 1076.430 1415.720 1172.590 ;
        RECT 1415.520 1076.110 1415.780 1076.430 ;
        RECT 1415.520 1075.430 1415.780 1075.750 ;
        RECT 1415.580 835.450 1415.720 1075.430 ;
        RECT 1415.120 835.310 1415.720 835.450 ;
        RECT 1415.120 834.770 1415.260 835.310 ;
        RECT 1415.120 834.630 1415.720 834.770 ;
        RECT 1415.580 773.685 1415.720 834.630 ;
        RECT 1415.510 773.315 1415.790 773.685 ;
        RECT 1415.510 772.635 1415.790 773.005 ;
        RECT 1415.580 724.870 1415.720 772.635 ;
        RECT 1415.520 724.550 1415.780 724.870 ;
        RECT 1415.060 724.210 1415.320 724.530 ;
        RECT 1415.120 710.590 1415.260 724.210 ;
        RECT 1415.060 710.270 1415.320 710.590 ;
        RECT 1415.520 662.330 1415.780 662.650 ;
        RECT 1415.580 628.845 1415.720 662.330 ;
        RECT 1415.510 628.475 1415.790 628.845 ;
        RECT 1415.510 627.795 1415.790 628.165 ;
        RECT 1415.580 594.050 1415.720 627.795 ;
        RECT 1415.580 593.910 1416.180 594.050 ;
        RECT 1416.040 572.890 1416.180 593.910 ;
        RECT 1415.520 572.570 1415.780 572.890 ;
        RECT 1415.980 572.570 1416.240 572.890 ;
        RECT 1415.580 548.750 1415.720 572.570 ;
        RECT 1414.600 548.430 1414.860 548.750 ;
        RECT 1415.520 548.430 1415.780 548.750 ;
        RECT 1414.660 524.270 1414.800 548.430 ;
        RECT 1414.600 523.950 1414.860 524.270 ;
        RECT 1414.600 476.010 1414.860 476.330 ;
        RECT 1414.660 458.730 1414.800 476.010 ;
        RECT 1414.660 458.590 1415.720 458.730 ;
        RECT 1415.580 353.330 1415.720 458.590 ;
        RECT 1415.580 353.190 1416.180 353.330 ;
        RECT 1416.040 331.830 1416.180 353.190 ;
        RECT 1415.980 331.510 1416.240 331.830 ;
        RECT 1415.520 282.890 1415.780 283.210 ;
        RECT 1415.580 234.500 1415.720 282.890 ;
        RECT 1415.580 234.360 1416.180 234.500 ;
        RECT 1416.040 227.790 1416.180 234.360 ;
        RECT 1415.980 227.470 1416.240 227.790 ;
        RECT 1414.600 179.530 1414.860 179.850 ;
        RECT 1414.660 158.170 1414.800 179.530 ;
        RECT 1414.660 158.030 1415.260 158.170 ;
        RECT 1415.120 53.030 1415.260 158.030 ;
        RECT 525.880 52.710 526.140 53.030 ;
        RECT 1415.060 52.710 1415.320 53.030 ;
        RECT 525.940 2.400 526.080 52.710 ;
        RECT 525.730 -4.800 526.290 2.400 ;
      LAYER via2 ;
        RECT 1415.510 773.360 1415.790 773.640 ;
        RECT 1415.510 772.680 1415.790 772.960 ;
        RECT 1415.510 628.520 1415.790 628.800 ;
        RECT 1415.510 627.840 1415.790 628.120 ;
      LAYER met3 ;
        RECT 1415.485 773.650 1415.815 773.665 ;
        RECT 1415.270 773.335 1415.815 773.650 ;
        RECT 1415.270 772.985 1415.570 773.335 ;
        RECT 1415.270 772.670 1415.815 772.985 ;
        RECT 1415.485 772.655 1415.815 772.670 ;
        RECT 1415.485 628.810 1415.815 628.825 ;
        RECT 1415.270 628.495 1415.815 628.810 ;
        RECT 1415.270 628.145 1415.570 628.495 ;
        RECT 1415.270 627.830 1415.815 628.145 ;
        RECT 1415.485 627.815 1415.815 627.830 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 543.790 52.600 544.110 52.660 ;
        RECT 1428.370 52.600 1428.690 52.660 ;
        RECT 543.790 52.460 1428.690 52.600 ;
        RECT 543.790 52.400 544.110 52.460 ;
        RECT 1428.370 52.400 1428.690 52.460 ;
      LAYER via ;
        RECT 543.820 52.400 544.080 52.660 ;
        RECT 1428.400 52.400 1428.660 52.660 ;
      LAYER met2 ;
        RECT 1428.320 1700.000 1428.600 1704.000 ;
        RECT 1428.460 52.690 1428.600 1700.000 ;
        RECT 543.820 52.370 544.080 52.690 ;
        RECT 1428.400 52.370 1428.660 52.690 ;
        RECT 543.880 2.400 544.020 52.370 ;
        RECT 543.670 -4.800 544.230 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 565.410 53.280 565.730 53.340 ;
        RECT 1435.270 53.280 1435.590 53.340 ;
        RECT 565.410 53.140 1435.590 53.280 ;
        RECT 565.410 53.080 565.730 53.140 ;
        RECT 1435.270 53.080 1435.590 53.140 ;
        RECT 561.730 14.860 562.050 14.920 ;
        RECT 565.410 14.860 565.730 14.920 ;
        RECT 561.730 14.720 565.730 14.860 ;
        RECT 561.730 14.660 562.050 14.720 ;
        RECT 565.410 14.660 565.730 14.720 ;
      LAYER via ;
        RECT 565.440 53.080 565.700 53.340 ;
        RECT 1435.300 53.080 1435.560 53.340 ;
        RECT 561.760 14.660 562.020 14.920 ;
        RECT 565.440 14.660 565.700 14.920 ;
      LAYER met2 ;
        RECT 1437.520 1700.410 1437.800 1704.000 ;
        RECT 1435.360 1700.270 1437.800 1700.410 ;
        RECT 1435.360 53.370 1435.500 1700.270 ;
        RECT 1437.520 1700.000 1437.800 1700.270 ;
        RECT 565.440 53.050 565.700 53.370 ;
        RECT 1435.300 53.050 1435.560 53.370 ;
        RECT 565.500 14.950 565.640 53.050 ;
        RECT 561.760 14.630 562.020 14.950 ;
        RECT 565.440 14.630 565.700 14.950 ;
        RECT 561.820 2.400 561.960 14.630 ;
        RECT 561.610 -4.800 562.170 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1443.165 1545.725 1443.335 1593.835 ;
        RECT 1443.165 1449.165 1443.335 1497.275 ;
        RECT 1443.165 1352.605 1443.335 1400.715 ;
        RECT 1443.165 1256.045 1443.335 1304.155 ;
        RECT 1443.165 483.225 1443.335 496.995 ;
        RECT 1443.165 386.325 1443.335 434.775 ;
        RECT 1442.705 53.465 1442.875 96.475 ;
      LAYER mcon ;
        RECT 1443.165 1593.665 1443.335 1593.835 ;
        RECT 1443.165 1497.105 1443.335 1497.275 ;
        RECT 1443.165 1400.545 1443.335 1400.715 ;
        RECT 1443.165 1303.985 1443.335 1304.155 ;
        RECT 1443.165 496.825 1443.335 496.995 ;
        RECT 1443.165 434.605 1443.335 434.775 ;
        RECT 1442.705 96.305 1442.875 96.475 ;
      LAYER met1 ;
        RECT 1443.090 1593.820 1443.410 1593.880 ;
        RECT 1442.895 1593.680 1443.410 1593.820 ;
        RECT 1443.090 1593.620 1443.410 1593.680 ;
        RECT 1443.090 1545.880 1443.410 1545.940 ;
        RECT 1442.895 1545.740 1443.410 1545.880 ;
        RECT 1443.090 1545.680 1443.410 1545.740 ;
        RECT 1443.090 1497.260 1443.410 1497.320 ;
        RECT 1442.895 1497.120 1443.410 1497.260 ;
        RECT 1443.090 1497.060 1443.410 1497.120 ;
        RECT 1443.090 1449.320 1443.410 1449.380 ;
        RECT 1442.895 1449.180 1443.410 1449.320 ;
        RECT 1443.090 1449.120 1443.410 1449.180 ;
        RECT 1443.090 1400.700 1443.410 1400.760 ;
        RECT 1442.895 1400.560 1443.410 1400.700 ;
        RECT 1443.090 1400.500 1443.410 1400.560 ;
        RECT 1443.090 1352.760 1443.410 1352.820 ;
        RECT 1442.895 1352.620 1443.410 1352.760 ;
        RECT 1443.090 1352.560 1443.410 1352.620 ;
        RECT 1443.090 1304.140 1443.410 1304.200 ;
        RECT 1442.895 1304.000 1443.410 1304.140 ;
        RECT 1443.090 1303.940 1443.410 1304.000 ;
        RECT 1443.090 1256.200 1443.410 1256.260 ;
        RECT 1442.895 1256.060 1443.410 1256.200 ;
        RECT 1443.090 1256.000 1443.410 1256.060 ;
        RECT 1442.170 1062.740 1442.490 1062.800 ;
        RECT 1443.090 1062.740 1443.410 1062.800 ;
        RECT 1442.170 1062.600 1443.410 1062.740 ;
        RECT 1442.170 1062.540 1442.490 1062.600 ;
        RECT 1443.090 1062.540 1443.410 1062.600 ;
        RECT 1442.170 966.180 1442.490 966.240 ;
        RECT 1443.090 966.180 1443.410 966.240 ;
        RECT 1442.170 966.040 1443.410 966.180 ;
        RECT 1442.170 965.980 1442.490 966.040 ;
        RECT 1443.090 965.980 1443.410 966.040 ;
        RECT 1442.170 869.620 1442.490 869.680 ;
        RECT 1443.090 869.620 1443.410 869.680 ;
        RECT 1442.170 869.480 1443.410 869.620 ;
        RECT 1442.170 869.420 1442.490 869.480 ;
        RECT 1443.090 869.420 1443.410 869.480 ;
        RECT 1443.090 496.980 1443.410 497.040 ;
        RECT 1442.895 496.840 1443.410 496.980 ;
        RECT 1443.090 496.780 1443.410 496.840 ;
        RECT 1443.090 483.380 1443.410 483.440 ;
        RECT 1442.895 483.240 1443.410 483.380 ;
        RECT 1443.090 483.180 1443.410 483.240 ;
        RECT 1443.090 434.760 1443.410 434.820 ;
        RECT 1442.895 434.620 1443.410 434.760 ;
        RECT 1443.090 434.560 1443.410 434.620 ;
        RECT 1443.090 386.480 1443.410 386.540 ;
        RECT 1442.895 386.340 1443.410 386.480 ;
        RECT 1443.090 386.280 1443.410 386.340 ;
        RECT 1442.630 234.500 1442.950 234.560 ;
        RECT 1443.090 234.500 1443.410 234.560 ;
        RECT 1442.630 234.360 1443.410 234.500 ;
        RECT 1442.630 234.300 1442.950 234.360 ;
        RECT 1443.090 234.300 1443.410 234.360 ;
        RECT 1442.170 144.740 1442.490 144.800 ;
        RECT 1443.090 144.740 1443.410 144.800 ;
        RECT 1442.170 144.600 1443.410 144.740 ;
        RECT 1442.170 144.540 1442.490 144.600 ;
        RECT 1443.090 144.540 1443.410 144.600 ;
        RECT 1442.630 96.460 1442.950 96.520 ;
        RECT 1442.435 96.320 1442.950 96.460 ;
        RECT 1442.630 96.260 1442.950 96.320 ;
        RECT 585.650 53.620 585.970 53.680 ;
        RECT 1442.645 53.620 1442.935 53.665 ;
        RECT 585.650 53.480 1442.935 53.620 ;
        RECT 585.650 53.420 585.970 53.480 ;
        RECT 1442.645 53.435 1442.935 53.480 ;
        RECT 579.670 14.860 579.990 14.920 ;
        RECT 584.730 14.860 585.050 14.920 ;
        RECT 579.670 14.720 585.050 14.860 ;
        RECT 579.670 14.660 579.990 14.720 ;
        RECT 584.730 14.660 585.050 14.720 ;
      LAYER via ;
        RECT 1443.120 1593.620 1443.380 1593.880 ;
        RECT 1443.120 1545.680 1443.380 1545.940 ;
        RECT 1443.120 1497.060 1443.380 1497.320 ;
        RECT 1443.120 1449.120 1443.380 1449.380 ;
        RECT 1443.120 1400.500 1443.380 1400.760 ;
        RECT 1443.120 1352.560 1443.380 1352.820 ;
        RECT 1443.120 1303.940 1443.380 1304.200 ;
        RECT 1443.120 1256.000 1443.380 1256.260 ;
        RECT 1442.200 1062.540 1442.460 1062.800 ;
        RECT 1443.120 1062.540 1443.380 1062.800 ;
        RECT 1442.200 965.980 1442.460 966.240 ;
        RECT 1443.120 965.980 1443.380 966.240 ;
        RECT 1442.200 869.420 1442.460 869.680 ;
        RECT 1443.120 869.420 1443.380 869.680 ;
        RECT 1443.120 496.780 1443.380 497.040 ;
        RECT 1443.120 483.180 1443.380 483.440 ;
        RECT 1443.120 434.560 1443.380 434.820 ;
        RECT 1443.120 386.280 1443.380 386.540 ;
        RECT 1442.660 234.300 1442.920 234.560 ;
        RECT 1443.120 234.300 1443.380 234.560 ;
        RECT 1442.200 144.540 1442.460 144.800 ;
        RECT 1443.120 144.540 1443.380 144.800 ;
        RECT 1442.660 96.260 1442.920 96.520 ;
        RECT 585.680 53.420 585.940 53.680 ;
        RECT 579.700 14.660 579.960 14.920 ;
        RECT 584.760 14.660 585.020 14.920 ;
      LAYER met2 ;
        RECT 1446.720 1701.090 1447.000 1704.000 ;
        RECT 1444.100 1700.950 1447.000 1701.090 ;
        RECT 1444.100 1677.970 1444.240 1700.950 ;
        RECT 1446.720 1700.000 1447.000 1700.950 ;
        RECT 1442.720 1677.830 1444.240 1677.970 ;
        RECT 1442.720 1606.570 1442.860 1677.830 ;
        RECT 1442.720 1606.430 1443.320 1606.570 ;
        RECT 1443.180 1593.910 1443.320 1606.430 ;
        RECT 1443.120 1593.590 1443.380 1593.910 ;
        RECT 1443.120 1545.650 1443.380 1545.970 ;
        RECT 1443.180 1497.350 1443.320 1545.650 ;
        RECT 1443.120 1497.030 1443.380 1497.350 ;
        RECT 1443.120 1449.090 1443.380 1449.410 ;
        RECT 1443.180 1400.790 1443.320 1449.090 ;
        RECT 1443.120 1400.470 1443.380 1400.790 ;
        RECT 1443.120 1352.530 1443.380 1352.850 ;
        RECT 1443.180 1304.230 1443.320 1352.530 ;
        RECT 1443.120 1303.910 1443.380 1304.230 ;
        RECT 1443.120 1255.970 1443.380 1256.290 ;
        RECT 1443.180 1173.410 1443.320 1255.970 ;
        RECT 1442.720 1173.270 1443.320 1173.410 ;
        RECT 1442.720 1172.730 1442.860 1173.270 ;
        RECT 1442.720 1172.590 1443.320 1172.730 ;
        RECT 1443.180 1110.965 1443.320 1172.590 ;
        RECT 1442.190 1110.595 1442.470 1110.965 ;
        RECT 1443.110 1110.595 1443.390 1110.965 ;
        RECT 1442.260 1062.830 1442.400 1110.595 ;
        RECT 1442.200 1062.510 1442.460 1062.830 ;
        RECT 1443.120 1062.510 1443.380 1062.830 ;
        RECT 1443.180 1014.405 1443.320 1062.510 ;
        RECT 1442.190 1014.035 1442.470 1014.405 ;
        RECT 1443.110 1014.035 1443.390 1014.405 ;
        RECT 1442.260 966.270 1442.400 1014.035 ;
        RECT 1442.200 965.950 1442.460 966.270 ;
        RECT 1443.120 965.950 1443.380 966.270 ;
        RECT 1443.180 917.845 1443.320 965.950 ;
        RECT 1442.190 917.475 1442.470 917.845 ;
        RECT 1443.110 917.475 1443.390 917.845 ;
        RECT 1442.260 869.710 1442.400 917.475 ;
        RECT 1442.200 869.390 1442.460 869.710 ;
        RECT 1443.120 869.390 1443.380 869.710 ;
        RECT 1443.180 787.170 1443.320 869.390 ;
        RECT 1442.720 787.030 1443.320 787.170 ;
        RECT 1442.720 785.810 1442.860 787.030 ;
        RECT 1442.720 785.670 1443.320 785.810 ;
        RECT 1443.180 690.610 1443.320 785.670 ;
        RECT 1442.720 690.470 1443.320 690.610 ;
        RECT 1442.720 689.930 1442.860 690.470 ;
        RECT 1442.720 689.790 1443.320 689.930 ;
        RECT 1443.180 628.845 1443.320 689.790 ;
        RECT 1443.110 628.475 1443.390 628.845 ;
        RECT 1443.110 627.795 1443.390 628.165 ;
        RECT 1443.180 594.050 1443.320 627.795 ;
        RECT 1443.180 593.910 1443.780 594.050 ;
        RECT 1443.640 592.690 1443.780 593.910 ;
        RECT 1443.180 592.550 1443.780 592.690 ;
        RECT 1443.180 497.070 1443.320 592.550 ;
        RECT 1443.120 496.750 1443.380 497.070 ;
        RECT 1443.120 483.150 1443.380 483.470 ;
        RECT 1443.180 434.850 1443.320 483.150 ;
        RECT 1443.120 434.530 1443.380 434.850 ;
        RECT 1443.120 386.250 1443.380 386.570 ;
        RECT 1443.180 235.010 1443.320 386.250 ;
        RECT 1442.720 234.870 1443.320 235.010 ;
        RECT 1442.720 234.590 1442.860 234.870 ;
        RECT 1442.660 234.270 1442.920 234.590 ;
        RECT 1443.120 234.270 1443.380 234.590 ;
        RECT 1443.180 144.830 1443.320 234.270 ;
        RECT 1442.200 144.510 1442.460 144.830 ;
        RECT 1443.120 144.510 1443.380 144.830 ;
        RECT 1442.260 96.970 1442.400 144.510 ;
        RECT 1442.260 96.830 1442.860 96.970 ;
        RECT 1442.720 96.550 1442.860 96.830 ;
        RECT 1442.660 96.230 1442.920 96.550 ;
        RECT 585.680 53.390 585.940 53.710 ;
        RECT 585.740 18.090 585.880 53.390 ;
        RECT 584.820 17.950 585.880 18.090 ;
        RECT 584.820 14.950 584.960 17.950 ;
        RECT 579.700 14.630 579.960 14.950 ;
        RECT 584.760 14.630 585.020 14.950 ;
        RECT 579.760 2.400 579.900 14.630 ;
        RECT 579.550 -4.800 580.110 2.400 ;
      LAYER via2 ;
        RECT 1442.190 1110.640 1442.470 1110.920 ;
        RECT 1443.110 1110.640 1443.390 1110.920 ;
        RECT 1442.190 1014.080 1442.470 1014.360 ;
        RECT 1443.110 1014.080 1443.390 1014.360 ;
        RECT 1442.190 917.520 1442.470 917.800 ;
        RECT 1443.110 917.520 1443.390 917.800 ;
        RECT 1443.110 628.520 1443.390 628.800 ;
        RECT 1443.110 627.840 1443.390 628.120 ;
      LAYER met3 ;
        RECT 1442.165 1110.930 1442.495 1110.945 ;
        RECT 1443.085 1110.930 1443.415 1110.945 ;
        RECT 1442.165 1110.630 1443.415 1110.930 ;
        RECT 1442.165 1110.615 1442.495 1110.630 ;
        RECT 1443.085 1110.615 1443.415 1110.630 ;
        RECT 1442.165 1014.370 1442.495 1014.385 ;
        RECT 1443.085 1014.370 1443.415 1014.385 ;
        RECT 1442.165 1014.070 1443.415 1014.370 ;
        RECT 1442.165 1014.055 1442.495 1014.070 ;
        RECT 1443.085 1014.055 1443.415 1014.070 ;
        RECT 1442.165 917.810 1442.495 917.825 ;
        RECT 1443.085 917.810 1443.415 917.825 ;
        RECT 1442.165 917.510 1443.415 917.810 ;
        RECT 1442.165 917.495 1442.495 917.510 ;
        RECT 1443.085 917.495 1443.415 917.510 ;
        RECT 1443.085 628.810 1443.415 628.825 ;
        RECT 1442.870 628.495 1443.415 628.810 ;
        RECT 1442.870 628.145 1443.170 628.495 ;
        RECT 1442.870 627.830 1443.415 628.145 ;
        RECT 1443.085 627.815 1443.415 627.830 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1187.330 1678.140 1187.650 1678.200 ;
        RECT 1191.470 1678.140 1191.790 1678.200 ;
        RECT 1187.330 1678.000 1191.790 1678.140 ;
        RECT 1187.330 1677.940 1187.650 1678.000 ;
        RECT 1191.470 1677.940 1191.790 1678.000 ;
        RECT 86.550 25.740 86.870 25.800 ;
        RECT 1187.330 25.740 1187.650 25.800 ;
        RECT 86.550 25.600 1187.650 25.740 ;
        RECT 86.550 25.540 86.870 25.600 ;
        RECT 1187.330 25.540 1187.650 25.600 ;
      LAYER via ;
        RECT 1187.360 1677.940 1187.620 1678.200 ;
        RECT 1191.500 1677.940 1191.760 1678.200 ;
        RECT 86.580 25.540 86.840 25.800 ;
        RECT 1187.360 25.540 1187.620 25.800 ;
      LAYER met2 ;
        RECT 1192.800 1700.410 1193.080 1704.000 ;
        RECT 1191.560 1700.270 1193.080 1700.410 ;
        RECT 1191.560 1678.230 1191.700 1700.270 ;
        RECT 1192.800 1700.000 1193.080 1700.270 ;
        RECT 1187.360 1677.910 1187.620 1678.230 ;
        RECT 1191.500 1677.910 1191.760 1678.230 ;
        RECT 1187.420 25.830 1187.560 1677.910 ;
        RECT 86.580 25.510 86.840 25.830 ;
        RECT 1187.360 25.510 1187.620 25.830 ;
        RECT 86.640 5.170 86.780 25.510 ;
        RECT 86.180 5.030 86.780 5.170 ;
        RECT 86.180 2.400 86.320 5.030 ;
        RECT 85.970 -4.800 86.530 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 599.910 53.960 600.230 54.020 ;
        RECT 1455.970 53.960 1456.290 54.020 ;
        RECT 599.910 53.820 1456.290 53.960 ;
        RECT 599.910 53.760 600.230 53.820 ;
        RECT 1455.970 53.760 1456.290 53.820 ;
        RECT 597.150 14.860 597.470 14.920 ;
        RECT 599.910 14.860 600.230 14.920 ;
        RECT 597.150 14.720 600.230 14.860 ;
        RECT 597.150 14.660 597.470 14.720 ;
        RECT 599.910 14.660 600.230 14.720 ;
      LAYER via ;
        RECT 599.940 53.760 600.200 54.020 ;
        RECT 1456.000 53.760 1456.260 54.020 ;
        RECT 597.180 14.660 597.440 14.920 ;
        RECT 599.940 14.660 600.200 14.920 ;
      LAYER met2 ;
        RECT 1455.920 1700.000 1456.200 1704.000 ;
        RECT 1456.060 54.050 1456.200 1700.000 ;
        RECT 599.940 53.730 600.200 54.050 ;
        RECT 1456.000 53.730 1456.260 54.050 ;
        RECT 600.000 14.950 600.140 53.730 ;
        RECT 597.180 14.630 597.440 14.950 ;
        RECT 599.940 14.630 600.200 14.950 ;
        RECT 597.240 2.400 597.380 14.630 ;
        RECT 597.030 -4.800 597.590 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 620.610 54.300 620.930 54.360 ;
        RECT 1462.870 54.300 1463.190 54.360 ;
        RECT 620.610 54.160 1463.190 54.300 ;
        RECT 620.610 54.100 620.930 54.160 ;
        RECT 1462.870 54.100 1463.190 54.160 ;
      LAYER via ;
        RECT 620.640 54.100 620.900 54.360 ;
        RECT 1462.900 54.100 1463.160 54.360 ;
      LAYER met2 ;
        RECT 1465.120 1700.410 1465.400 1704.000 ;
        RECT 1462.960 1700.270 1465.400 1700.410 ;
        RECT 1462.960 54.390 1463.100 1700.270 ;
        RECT 1465.120 1700.000 1465.400 1700.270 ;
        RECT 620.640 54.070 620.900 54.390 ;
        RECT 1462.900 54.070 1463.160 54.390 ;
        RECT 620.700 17.410 620.840 54.070 ;
        RECT 615.180 17.270 620.840 17.410 ;
        RECT 615.180 2.400 615.320 17.270 ;
        RECT 614.970 -4.800 615.530 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1200.745 572.645 1200.915 620.755 ;
        RECT 1200.745 483.225 1200.915 531.335 ;
        RECT 1200.745 428.145 1200.915 475.915 ;
        RECT 1201.205 234.685 1201.375 282.795 ;
        RECT 1201.205 131.665 1201.375 159.375 ;
      LAYER mcon ;
        RECT 1200.745 620.585 1200.915 620.755 ;
        RECT 1200.745 531.165 1200.915 531.335 ;
        RECT 1200.745 475.745 1200.915 475.915 ;
        RECT 1201.205 282.625 1201.375 282.795 ;
        RECT 1201.205 159.205 1201.375 159.375 ;
      LAYER met1 ;
        RECT 1201.130 765.920 1201.450 765.980 ;
        RECT 1202.510 765.920 1202.830 765.980 ;
        RECT 1201.130 765.780 1202.830 765.920 ;
        RECT 1201.130 765.720 1201.450 765.780 ;
        RECT 1202.510 765.720 1202.830 765.780 ;
        RECT 1200.670 628.220 1200.990 628.280 ;
        RECT 1201.590 628.220 1201.910 628.280 ;
        RECT 1200.670 628.080 1201.910 628.220 ;
        RECT 1200.670 628.020 1200.990 628.080 ;
        RECT 1201.590 628.020 1201.910 628.080 ;
        RECT 1200.670 620.740 1200.990 620.800 ;
        RECT 1200.670 620.600 1201.185 620.740 ;
        RECT 1200.670 620.540 1200.990 620.600 ;
        RECT 1200.685 572.800 1200.975 572.845 ;
        RECT 1201.130 572.800 1201.450 572.860 ;
        RECT 1200.685 572.660 1201.450 572.800 ;
        RECT 1200.685 572.615 1200.975 572.660 ;
        RECT 1201.130 572.600 1201.450 572.660 ;
        RECT 1200.685 531.320 1200.975 531.365 ;
        RECT 1201.130 531.320 1201.450 531.380 ;
        RECT 1200.685 531.180 1201.450 531.320 ;
        RECT 1200.685 531.135 1200.975 531.180 ;
        RECT 1201.130 531.120 1201.450 531.180 ;
        RECT 1200.670 483.380 1200.990 483.440 ;
        RECT 1200.475 483.240 1200.990 483.380 ;
        RECT 1200.670 483.180 1200.990 483.240 ;
        RECT 1200.670 475.900 1200.990 475.960 ;
        RECT 1200.670 475.760 1201.185 475.900 ;
        RECT 1200.670 475.700 1200.990 475.760 ;
        RECT 1200.685 428.300 1200.975 428.345 ;
        RECT 1201.130 428.300 1201.450 428.360 ;
        RECT 1200.685 428.160 1201.450 428.300 ;
        RECT 1200.685 428.115 1200.975 428.160 ;
        RECT 1201.130 428.100 1201.450 428.160 ;
        RECT 1201.130 379.680 1201.450 379.740 ;
        RECT 1202.050 379.680 1202.370 379.740 ;
        RECT 1201.130 379.540 1202.370 379.680 ;
        RECT 1201.130 379.480 1201.450 379.540 ;
        RECT 1202.050 379.480 1202.370 379.540 ;
        RECT 1200.670 338.200 1200.990 338.260 ;
        RECT 1201.590 338.200 1201.910 338.260 ;
        RECT 1200.670 338.060 1201.910 338.200 ;
        RECT 1200.670 338.000 1200.990 338.060 ;
        RECT 1201.590 338.000 1201.910 338.060 ;
        RECT 1200.670 289.920 1200.990 289.980 ;
        RECT 1201.130 289.920 1201.450 289.980 ;
        RECT 1200.670 289.780 1201.450 289.920 ;
        RECT 1200.670 289.720 1200.990 289.780 ;
        RECT 1201.130 289.720 1201.450 289.780 ;
        RECT 1201.130 282.780 1201.450 282.840 ;
        RECT 1200.935 282.640 1201.450 282.780 ;
        RECT 1201.130 282.580 1201.450 282.640 ;
        RECT 1201.130 234.840 1201.450 234.900 ;
        RECT 1200.935 234.700 1201.450 234.840 ;
        RECT 1201.130 234.640 1201.450 234.700 ;
        RECT 1201.130 159.360 1201.450 159.420 ;
        RECT 1200.935 159.220 1201.450 159.360 ;
        RECT 1201.130 159.160 1201.450 159.220 ;
        RECT 1201.130 131.820 1201.450 131.880 ;
        RECT 1200.935 131.680 1201.450 131.820 ;
        RECT 1201.130 131.620 1201.450 131.680 ;
        RECT 1201.130 130.940 1201.450 131.200 ;
        RECT 1201.220 130.800 1201.360 130.940 ;
        RECT 1201.590 130.800 1201.910 130.860 ;
        RECT 1201.220 130.660 1201.910 130.800 ;
        RECT 1201.590 130.600 1201.910 130.660 ;
        RECT 109.550 26.080 109.870 26.140 ;
        RECT 1201.130 26.080 1201.450 26.140 ;
        RECT 109.550 25.940 1201.450 26.080 ;
        RECT 109.550 25.880 109.870 25.940 ;
        RECT 1201.130 25.880 1201.450 25.940 ;
      LAYER via ;
        RECT 1201.160 765.720 1201.420 765.980 ;
        RECT 1202.540 765.720 1202.800 765.980 ;
        RECT 1200.700 628.020 1200.960 628.280 ;
        RECT 1201.620 628.020 1201.880 628.280 ;
        RECT 1200.700 620.540 1200.960 620.800 ;
        RECT 1201.160 572.600 1201.420 572.860 ;
        RECT 1201.160 531.120 1201.420 531.380 ;
        RECT 1200.700 483.180 1200.960 483.440 ;
        RECT 1200.700 475.700 1200.960 475.960 ;
        RECT 1201.160 428.100 1201.420 428.360 ;
        RECT 1201.160 379.480 1201.420 379.740 ;
        RECT 1202.080 379.480 1202.340 379.740 ;
        RECT 1200.700 338.000 1200.960 338.260 ;
        RECT 1201.620 338.000 1201.880 338.260 ;
        RECT 1200.700 289.720 1200.960 289.980 ;
        RECT 1201.160 289.720 1201.420 289.980 ;
        RECT 1201.160 282.580 1201.420 282.840 ;
        RECT 1201.160 234.640 1201.420 234.900 ;
        RECT 1201.160 159.160 1201.420 159.420 ;
        RECT 1201.160 131.620 1201.420 131.880 ;
        RECT 1201.160 130.940 1201.420 131.200 ;
        RECT 1201.620 130.600 1201.880 130.860 ;
        RECT 109.580 25.880 109.840 26.140 ;
        RECT 1201.160 25.880 1201.420 26.140 ;
      LAYER met2 ;
        RECT 1204.760 1701.090 1205.040 1704.000 ;
        RECT 1202.600 1700.950 1205.040 1701.090 ;
        RECT 1202.600 1656.210 1202.740 1700.950 ;
        RECT 1204.760 1700.000 1205.040 1700.950 ;
        RECT 1200.760 1656.070 1202.740 1656.210 ;
        RECT 1200.760 1655.530 1200.900 1656.070 ;
        RECT 1200.760 1655.390 1201.360 1655.530 ;
        RECT 1201.220 1511.370 1201.360 1655.390 ;
        RECT 1200.760 1511.230 1201.360 1511.370 ;
        RECT 1200.760 1510.690 1200.900 1511.230 ;
        RECT 1200.760 1510.550 1201.360 1510.690 ;
        RECT 1201.220 1414.810 1201.360 1510.550 ;
        RECT 1200.760 1414.670 1201.360 1414.810 ;
        RECT 1200.760 1414.130 1200.900 1414.670 ;
        RECT 1200.760 1413.990 1201.360 1414.130 ;
        RECT 1201.220 1318.250 1201.360 1413.990 ;
        RECT 1200.760 1318.110 1201.360 1318.250 ;
        RECT 1200.760 1317.570 1200.900 1318.110 ;
        RECT 1200.760 1317.430 1201.360 1317.570 ;
        RECT 1201.220 1221.690 1201.360 1317.430 ;
        RECT 1200.760 1221.550 1201.360 1221.690 ;
        RECT 1200.760 1221.010 1200.900 1221.550 ;
        RECT 1200.760 1220.870 1201.360 1221.010 ;
        RECT 1201.220 1125.130 1201.360 1220.870 ;
        RECT 1200.760 1124.990 1201.360 1125.130 ;
        RECT 1200.760 1124.450 1200.900 1124.990 ;
        RECT 1200.760 1124.310 1201.360 1124.450 ;
        RECT 1201.220 1028.570 1201.360 1124.310 ;
        RECT 1200.760 1028.430 1201.360 1028.570 ;
        RECT 1200.760 1027.890 1200.900 1028.430 ;
        RECT 1200.760 1027.750 1201.360 1027.890 ;
        RECT 1201.220 932.010 1201.360 1027.750 ;
        RECT 1200.760 931.870 1201.360 932.010 ;
        RECT 1200.760 931.330 1200.900 931.870 ;
        RECT 1200.760 931.190 1201.360 931.330 ;
        RECT 1201.220 835.450 1201.360 931.190 ;
        RECT 1200.760 835.310 1201.360 835.450 ;
        RECT 1200.760 834.770 1200.900 835.310 ;
        RECT 1200.760 834.630 1201.360 834.770 ;
        RECT 1201.220 773.685 1201.360 834.630 ;
        RECT 1201.150 773.315 1201.430 773.685 ;
        RECT 1201.150 772.635 1201.430 773.005 ;
        RECT 1201.220 766.010 1201.360 772.635 ;
        RECT 1201.160 765.690 1201.420 766.010 ;
        RECT 1202.540 765.690 1202.800 766.010 ;
        RECT 1202.600 717.925 1202.740 765.690 ;
        RECT 1201.610 717.555 1201.890 717.925 ;
        RECT 1202.530 717.555 1202.810 717.925 ;
        RECT 1201.680 628.310 1201.820 717.555 ;
        RECT 1200.700 627.990 1200.960 628.310 ;
        RECT 1201.620 627.990 1201.880 628.310 ;
        RECT 1200.760 620.830 1200.900 627.990 ;
        RECT 1200.700 620.510 1200.960 620.830 ;
        RECT 1201.160 572.570 1201.420 572.890 ;
        RECT 1201.220 531.410 1201.360 572.570 ;
        RECT 1201.160 531.090 1201.420 531.410 ;
        RECT 1200.700 483.150 1200.960 483.470 ;
        RECT 1200.760 475.990 1200.900 483.150 ;
        RECT 1200.700 475.670 1200.960 475.990 ;
        RECT 1201.160 428.070 1201.420 428.390 ;
        RECT 1201.220 427.620 1201.360 428.070 ;
        RECT 1201.220 427.480 1202.280 427.620 ;
        RECT 1202.140 379.770 1202.280 427.480 ;
        RECT 1201.160 379.450 1201.420 379.770 ;
        RECT 1202.080 379.450 1202.340 379.770 ;
        RECT 1201.220 362.850 1201.360 379.450 ;
        RECT 1201.220 362.710 1201.820 362.850 ;
        RECT 1201.680 338.290 1201.820 362.710 ;
        RECT 1200.700 337.970 1200.960 338.290 ;
        RECT 1201.620 337.970 1201.880 338.290 ;
        RECT 1200.760 290.010 1200.900 337.970 ;
        RECT 1200.700 289.690 1200.960 290.010 ;
        RECT 1201.160 289.690 1201.420 290.010 ;
        RECT 1201.220 282.870 1201.360 289.690 ;
        RECT 1201.160 282.550 1201.420 282.870 ;
        RECT 1201.160 234.610 1201.420 234.930 ;
        RECT 1201.220 159.450 1201.360 234.610 ;
        RECT 1201.160 159.130 1201.420 159.450 ;
        RECT 1201.160 131.590 1201.420 131.910 ;
        RECT 1201.220 131.230 1201.360 131.590 ;
        RECT 1201.160 130.910 1201.420 131.230 ;
        RECT 1201.620 130.570 1201.880 130.890 ;
        RECT 1201.680 61.610 1201.820 130.570 ;
        RECT 1201.220 61.470 1201.820 61.610 ;
        RECT 1201.220 26.170 1201.360 61.470 ;
        RECT 109.580 25.850 109.840 26.170 ;
        RECT 1201.160 25.850 1201.420 26.170 ;
        RECT 109.640 2.400 109.780 25.850 ;
        RECT 109.430 -4.800 109.990 2.400 ;
      LAYER via2 ;
        RECT 1201.150 773.360 1201.430 773.640 ;
        RECT 1201.150 772.680 1201.430 772.960 ;
        RECT 1201.610 717.600 1201.890 717.880 ;
        RECT 1202.530 717.600 1202.810 717.880 ;
      LAYER met3 ;
        RECT 1201.125 773.650 1201.455 773.665 ;
        RECT 1200.910 773.335 1201.455 773.650 ;
        RECT 1200.910 772.985 1201.210 773.335 ;
        RECT 1200.910 772.670 1201.455 772.985 ;
        RECT 1201.125 772.655 1201.455 772.670 ;
        RECT 1201.585 717.890 1201.915 717.905 ;
        RECT 1202.505 717.890 1202.835 717.905 ;
        RECT 1201.585 717.590 1202.835 717.890 ;
        RECT 1201.585 717.575 1201.915 717.590 ;
        RECT 1202.505 717.575 1202.835 717.590 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 133.470 38.660 133.790 38.720 ;
        RECT 1214.470 38.660 1214.790 38.720 ;
        RECT 133.470 38.520 1214.790 38.660 ;
        RECT 133.470 38.460 133.790 38.520 ;
        RECT 1214.470 38.460 1214.790 38.520 ;
      LAYER via ;
        RECT 133.500 38.460 133.760 38.720 ;
        RECT 1214.500 38.460 1214.760 38.720 ;
      LAYER met2 ;
        RECT 1217.180 1700.410 1217.460 1704.000 ;
        RECT 1214.560 1700.270 1217.460 1700.410 ;
        RECT 1214.560 38.750 1214.700 1700.270 ;
        RECT 1217.180 1700.000 1217.460 1700.270 ;
        RECT 133.500 38.430 133.760 38.750 ;
        RECT 1214.500 38.430 1214.760 38.750 ;
        RECT 133.560 2.400 133.700 38.430 ;
        RECT 133.350 -4.800 133.910 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1222.365 338.045 1222.535 352.495 ;
        RECT 1222.365 186.405 1222.535 234.515 ;
        RECT 1221.445 83.045 1221.615 97.155 ;
      LAYER mcon ;
        RECT 1222.365 352.325 1222.535 352.495 ;
        RECT 1222.365 234.345 1222.535 234.515 ;
        RECT 1221.445 96.985 1221.615 97.155 ;
      LAYER met1 ;
        RECT 1222.290 1462.380 1222.610 1462.640 ;
        RECT 1222.380 1461.960 1222.520 1462.380 ;
        RECT 1222.290 1461.700 1222.610 1461.960 ;
        RECT 1222.290 1365.820 1222.610 1366.080 ;
        RECT 1222.380 1365.400 1222.520 1365.820 ;
        RECT 1222.290 1365.140 1222.610 1365.400 ;
        RECT 1222.290 1269.260 1222.610 1269.520 ;
        RECT 1222.380 1268.840 1222.520 1269.260 ;
        RECT 1222.290 1268.580 1222.610 1268.840 ;
        RECT 1222.290 883.020 1222.610 883.280 ;
        RECT 1222.380 882.600 1222.520 883.020 ;
        RECT 1222.290 882.340 1222.610 882.600 ;
        RECT 1221.830 593.540 1222.150 593.600 ;
        RECT 1221.830 593.400 1222.520 593.540 ;
        RECT 1221.830 593.340 1222.150 593.400 ;
        RECT 1222.380 593.260 1222.520 593.400 ;
        RECT 1222.290 593.000 1222.610 593.260 ;
        RECT 1222.290 497.120 1222.610 497.380 ;
        RECT 1222.380 496.700 1222.520 497.120 ;
        RECT 1222.290 496.440 1222.610 496.700 ;
        RECT 1222.290 352.480 1222.610 352.540 ;
        RECT 1222.095 352.340 1222.610 352.480 ;
        RECT 1222.290 352.280 1222.610 352.340 ;
        RECT 1222.290 338.200 1222.610 338.260 ;
        RECT 1222.095 338.060 1222.610 338.200 ;
        RECT 1222.290 338.000 1222.610 338.060 ;
        RECT 1221.830 289.920 1222.150 289.980 ;
        RECT 1222.750 289.920 1223.070 289.980 ;
        RECT 1221.830 289.780 1223.070 289.920 ;
        RECT 1221.830 289.720 1222.150 289.780 ;
        RECT 1222.750 289.720 1223.070 289.780 ;
        RECT 1222.290 234.500 1222.610 234.560 ;
        RECT 1222.095 234.360 1222.610 234.500 ;
        RECT 1222.290 234.300 1222.610 234.360 ;
        RECT 1222.305 186.560 1222.595 186.605 ;
        RECT 1222.750 186.560 1223.070 186.620 ;
        RECT 1222.305 186.420 1223.070 186.560 ;
        RECT 1222.305 186.375 1222.595 186.420 ;
        RECT 1222.750 186.360 1223.070 186.420 ;
        RECT 1221.830 145.080 1222.150 145.140 ;
        RECT 1222.750 145.080 1223.070 145.140 ;
        RECT 1221.830 144.940 1223.070 145.080 ;
        RECT 1221.830 144.880 1222.150 144.940 ;
        RECT 1222.750 144.880 1223.070 144.940 ;
        RECT 1221.385 97.140 1221.675 97.185 ;
        RECT 1221.830 97.140 1222.150 97.200 ;
        RECT 1221.385 97.000 1222.150 97.140 ;
        RECT 1221.385 96.955 1221.675 97.000 ;
        RECT 1221.830 96.940 1222.150 97.000 ;
        RECT 1221.370 83.200 1221.690 83.260 ;
        RECT 1221.175 83.060 1221.690 83.200 ;
        RECT 1221.370 83.000 1221.690 83.060 ;
        RECT 151.410 39.000 151.730 39.060 ;
        RECT 1221.370 39.000 1221.690 39.060 ;
        RECT 151.410 38.860 1221.690 39.000 ;
        RECT 151.410 38.800 151.730 38.860 ;
        RECT 1221.370 38.800 1221.690 38.860 ;
      LAYER via ;
        RECT 1222.320 1462.380 1222.580 1462.640 ;
        RECT 1222.320 1461.700 1222.580 1461.960 ;
        RECT 1222.320 1365.820 1222.580 1366.080 ;
        RECT 1222.320 1365.140 1222.580 1365.400 ;
        RECT 1222.320 1269.260 1222.580 1269.520 ;
        RECT 1222.320 1268.580 1222.580 1268.840 ;
        RECT 1222.320 883.020 1222.580 883.280 ;
        RECT 1222.320 882.340 1222.580 882.600 ;
        RECT 1221.860 593.340 1222.120 593.600 ;
        RECT 1222.320 593.000 1222.580 593.260 ;
        RECT 1222.320 497.120 1222.580 497.380 ;
        RECT 1222.320 496.440 1222.580 496.700 ;
        RECT 1222.320 352.280 1222.580 352.540 ;
        RECT 1222.320 338.000 1222.580 338.260 ;
        RECT 1221.860 289.720 1222.120 289.980 ;
        RECT 1222.780 289.720 1223.040 289.980 ;
        RECT 1222.320 234.300 1222.580 234.560 ;
        RECT 1222.780 186.360 1223.040 186.620 ;
        RECT 1221.860 144.880 1222.120 145.140 ;
        RECT 1222.780 144.880 1223.040 145.140 ;
        RECT 1221.860 96.940 1222.120 97.200 ;
        RECT 1221.400 83.000 1221.660 83.260 ;
        RECT 151.440 38.800 151.700 39.060 ;
        RECT 1221.400 38.800 1221.660 39.060 ;
      LAYER met2 ;
        RECT 1226.380 1700.410 1226.660 1704.000 ;
        RECT 1224.220 1700.270 1226.660 1700.410 ;
        RECT 1224.220 1678.650 1224.360 1700.270 ;
        RECT 1226.380 1700.000 1226.660 1700.270 ;
        RECT 1222.380 1678.510 1224.360 1678.650 ;
        RECT 1222.380 1559.650 1222.520 1678.510 ;
        RECT 1221.920 1559.510 1222.520 1559.650 ;
        RECT 1221.920 1558.970 1222.060 1559.510 ;
        RECT 1221.920 1558.830 1222.520 1558.970 ;
        RECT 1222.380 1462.670 1222.520 1558.830 ;
        RECT 1222.320 1462.350 1222.580 1462.670 ;
        RECT 1222.320 1461.670 1222.580 1461.990 ;
        RECT 1222.380 1366.110 1222.520 1461.670 ;
        RECT 1222.320 1365.790 1222.580 1366.110 ;
        RECT 1222.320 1365.110 1222.580 1365.430 ;
        RECT 1222.380 1269.550 1222.520 1365.110 ;
        RECT 1222.320 1269.230 1222.580 1269.550 ;
        RECT 1222.320 1268.550 1222.580 1268.870 ;
        RECT 1222.380 883.310 1222.520 1268.550 ;
        RECT 1222.320 882.990 1222.580 883.310 ;
        RECT 1222.320 882.310 1222.580 882.630 ;
        RECT 1222.380 677.125 1222.520 882.310 ;
        RECT 1222.310 676.755 1222.590 677.125 ;
        RECT 1222.310 675.395 1222.590 675.765 ;
        RECT 1222.380 620.740 1222.520 675.395 ;
        RECT 1221.920 620.600 1222.520 620.740 ;
        RECT 1221.920 593.630 1222.060 620.600 ;
        RECT 1221.860 593.310 1222.120 593.630 ;
        RECT 1222.320 592.970 1222.580 593.290 ;
        RECT 1222.380 497.410 1222.520 592.970 ;
        RECT 1222.320 497.090 1222.580 497.410 ;
        RECT 1222.320 496.410 1222.580 496.730 ;
        RECT 1222.380 352.570 1222.520 496.410 ;
        RECT 1222.320 352.250 1222.580 352.570 ;
        RECT 1222.320 337.970 1222.580 338.290 ;
        RECT 1222.380 314.570 1222.520 337.970 ;
        RECT 1222.380 314.430 1222.980 314.570 ;
        RECT 1222.840 290.010 1222.980 314.430 ;
        RECT 1221.860 289.690 1222.120 290.010 ;
        RECT 1222.780 289.690 1223.040 290.010 ;
        RECT 1221.920 254.730 1222.060 289.690 ;
        RECT 1221.920 254.590 1222.520 254.730 ;
        RECT 1222.380 234.590 1222.520 254.590 ;
        RECT 1222.320 234.270 1222.580 234.590 ;
        RECT 1222.780 186.330 1223.040 186.650 ;
        RECT 1222.840 145.170 1222.980 186.330 ;
        RECT 1221.860 144.850 1222.120 145.170 ;
        RECT 1222.780 144.850 1223.040 145.170 ;
        RECT 1221.920 97.230 1222.060 144.850 ;
        RECT 1221.860 96.910 1222.120 97.230 ;
        RECT 1221.400 82.970 1221.660 83.290 ;
        RECT 1221.460 39.090 1221.600 82.970 ;
        RECT 151.440 38.770 151.700 39.090 ;
        RECT 1221.400 38.770 1221.660 39.090 ;
        RECT 151.500 2.400 151.640 38.770 ;
        RECT 151.290 -4.800 151.850 2.400 ;
      LAYER via2 ;
        RECT 1222.310 676.800 1222.590 677.080 ;
        RECT 1222.310 675.440 1222.590 675.720 ;
      LAYER met3 ;
        RECT 1222.285 677.090 1222.615 677.105 ;
        RECT 1222.070 676.775 1222.615 677.090 ;
        RECT 1222.070 675.745 1222.370 676.775 ;
        RECT 1222.070 675.430 1222.615 675.745 ;
        RECT 1222.285 675.415 1222.615 675.430 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 169.350 39.340 169.670 39.400 ;
        RECT 1236.090 39.340 1236.410 39.400 ;
        RECT 169.350 39.200 1236.410 39.340 ;
        RECT 169.350 39.140 169.670 39.200 ;
        RECT 1236.090 39.140 1236.410 39.200 ;
      LAYER via ;
        RECT 169.380 39.140 169.640 39.400 ;
        RECT 1236.120 39.140 1236.380 39.400 ;
      LAYER met2 ;
        RECT 1235.580 1700.410 1235.860 1704.000 ;
        RECT 1235.580 1700.270 1236.320 1700.410 ;
        RECT 1235.580 1700.000 1235.860 1700.270 ;
        RECT 1236.180 39.430 1236.320 1700.270 ;
        RECT 169.380 39.110 169.640 39.430 ;
        RECT 1236.120 39.110 1236.380 39.430 ;
        RECT 169.440 2.400 169.580 39.110 ;
        RECT 169.230 -4.800 169.790 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 186.830 39.680 187.150 39.740 ;
        RECT 1242.530 39.680 1242.850 39.740 ;
        RECT 186.830 39.540 1242.850 39.680 ;
        RECT 186.830 39.480 187.150 39.540 ;
        RECT 1242.530 39.480 1242.850 39.540 ;
      LAYER via ;
        RECT 186.860 39.480 187.120 39.740 ;
        RECT 1242.560 39.480 1242.820 39.740 ;
      LAYER met2 ;
        RECT 1244.780 1700.410 1245.060 1704.000 ;
        RECT 1242.620 1700.270 1245.060 1700.410 ;
        RECT 1242.620 39.770 1242.760 1700.270 ;
        RECT 1244.780 1700.000 1245.060 1700.270 ;
        RECT 186.860 39.450 187.120 39.770 ;
        RECT 1242.560 39.450 1242.820 39.770 ;
        RECT 186.920 2.400 187.060 39.450 ;
        RECT 186.710 -4.800 187.270 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1249.965 1587.205 1250.135 1608.455 ;
        RECT 1249.965 1449.165 1250.135 1497.275 ;
        RECT 1249.965 572.645 1250.135 620.755 ;
        RECT 1249.965 396.525 1250.135 427.635 ;
        RECT 1249.505 282.625 1249.675 324.275 ;
        RECT 1249.505 235.025 1249.675 255.935 ;
        RECT 1249.505 186.405 1249.675 234.515 ;
      LAYER mcon ;
        RECT 1249.965 1608.285 1250.135 1608.455 ;
        RECT 1249.965 1497.105 1250.135 1497.275 ;
        RECT 1249.965 620.585 1250.135 620.755 ;
        RECT 1249.965 427.465 1250.135 427.635 ;
        RECT 1249.505 324.105 1249.675 324.275 ;
        RECT 1249.505 255.765 1249.675 255.935 ;
        RECT 1249.505 234.345 1249.675 234.515 ;
      LAYER met1 ;
        RECT 1249.890 1608.440 1250.210 1608.500 ;
        RECT 1249.695 1608.300 1250.210 1608.440 ;
        RECT 1249.890 1608.240 1250.210 1608.300 ;
        RECT 1249.890 1587.360 1250.210 1587.420 ;
        RECT 1249.695 1587.220 1250.210 1587.360 ;
        RECT 1249.890 1587.160 1250.210 1587.220 ;
        RECT 1249.430 1562.880 1249.750 1562.940 ;
        RECT 1250.350 1562.880 1250.670 1562.940 ;
        RECT 1249.430 1562.740 1250.670 1562.880 ;
        RECT 1249.430 1562.680 1249.750 1562.740 ;
        RECT 1250.350 1562.680 1250.670 1562.740 ;
        RECT 1249.890 1497.260 1250.210 1497.320 ;
        RECT 1249.695 1497.120 1250.210 1497.260 ;
        RECT 1249.890 1497.060 1250.210 1497.120 ;
        RECT 1249.890 1449.320 1250.210 1449.380 ;
        RECT 1249.695 1449.180 1250.210 1449.320 ;
        RECT 1249.890 1449.120 1250.210 1449.180 ;
        RECT 1249.890 1365.140 1250.210 1365.400 ;
        RECT 1249.980 1364.720 1250.120 1365.140 ;
        RECT 1249.890 1364.460 1250.210 1364.720 ;
        RECT 1249.890 1268.580 1250.210 1268.840 ;
        RECT 1249.980 1268.160 1250.120 1268.580 ;
        RECT 1249.890 1267.900 1250.210 1268.160 ;
        RECT 1249.890 882.340 1250.210 882.600 ;
        RECT 1249.980 881.920 1250.120 882.340 ;
        RECT 1249.890 881.660 1250.210 881.920 ;
        RECT 1249.890 620.740 1250.210 620.800 ;
        RECT 1249.695 620.600 1250.210 620.740 ;
        RECT 1249.890 620.540 1250.210 620.600 ;
        RECT 1249.890 572.800 1250.210 572.860 ;
        RECT 1249.695 572.660 1250.210 572.800 ;
        RECT 1249.890 572.600 1250.210 572.660 ;
        RECT 1249.890 427.620 1250.210 427.680 ;
        RECT 1249.695 427.480 1250.210 427.620 ;
        RECT 1249.890 427.420 1250.210 427.480 ;
        RECT 1249.890 396.680 1250.210 396.740 ;
        RECT 1249.695 396.540 1250.210 396.680 ;
        RECT 1249.890 396.480 1250.210 396.540 ;
        RECT 1249.430 331.060 1249.750 331.120 ;
        RECT 1249.890 331.060 1250.210 331.120 ;
        RECT 1249.430 330.920 1250.210 331.060 ;
        RECT 1249.430 330.860 1249.750 330.920 ;
        RECT 1249.890 330.860 1250.210 330.920 ;
        RECT 1249.430 324.260 1249.750 324.320 ;
        RECT 1249.235 324.120 1249.750 324.260 ;
        RECT 1249.430 324.060 1249.750 324.120 ;
        RECT 1249.430 282.780 1249.750 282.840 ;
        RECT 1249.235 282.640 1249.750 282.780 ;
        RECT 1249.430 282.580 1249.750 282.640 ;
        RECT 1249.430 255.920 1249.750 255.980 ;
        RECT 1249.235 255.780 1249.750 255.920 ;
        RECT 1249.430 255.720 1249.750 255.780 ;
        RECT 1249.430 235.180 1249.750 235.240 ;
        RECT 1249.235 235.040 1249.750 235.180 ;
        RECT 1249.430 234.980 1249.750 235.040 ;
        RECT 1249.430 234.500 1249.750 234.560 ;
        RECT 1249.235 234.360 1249.750 234.500 ;
        RECT 1249.430 234.300 1249.750 234.360 ;
        RECT 1249.430 186.560 1249.750 186.620 ;
        RECT 1249.235 186.420 1249.750 186.560 ;
        RECT 1249.430 186.360 1249.750 186.420 ;
        RECT 1249.430 145.080 1249.750 145.140 ;
        RECT 1249.890 145.080 1250.210 145.140 ;
        RECT 1249.430 144.940 1250.210 145.080 ;
        RECT 1249.430 144.880 1249.750 144.940 ;
        RECT 1249.890 144.880 1250.210 144.940 ;
        RECT 1249.890 48.520 1250.210 48.580 ;
        RECT 1250.350 48.520 1250.670 48.580 ;
        RECT 1249.890 48.380 1250.670 48.520 ;
        RECT 1249.890 48.320 1250.210 48.380 ;
        RECT 1250.350 48.320 1250.670 48.380 ;
        RECT 204.770 40.020 205.090 40.080 ;
        RECT 1249.890 40.020 1250.210 40.080 ;
        RECT 204.770 39.880 1250.210 40.020 ;
        RECT 204.770 39.820 205.090 39.880 ;
        RECT 1249.890 39.820 1250.210 39.880 ;
      LAYER via ;
        RECT 1249.920 1608.240 1250.180 1608.500 ;
        RECT 1249.920 1587.160 1250.180 1587.420 ;
        RECT 1249.460 1562.680 1249.720 1562.940 ;
        RECT 1250.380 1562.680 1250.640 1562.940 ;
        RECT 1249.920 1497.060 1250.180 1497.320 ;
        RECT 1249.920 1449.120 1250.180 1449.380 ;
        RECT 1249.920 1365.140 1250.180 1365.400 ;
        RECT 1249.920 1364.460 1250.180 1364.720 ;
        RECT 1249.920 1268.580 1250.180 1268.840 ;
        RECT 1249.920 1267.900 1250.180 1268.160 ;
        RECT 1249.920 882.340 1250.180 882.600 ;
        RECT 1249.920 881.660 1250.180 881.920 ;
        RECT 1249.920 620.540 1250.180 620.800 ;
        RECT 1249.920 572.600 1250.180 572.860 ;
        RECT 1249.920 427.420 1250.180 427.680 ;
        RECT 1249.920 396.480 1250.180 396.740 ;
        RECT 1249.460 330.860 1249.720 331.120 ;
        RECT 1249.920 330.860 1250.180 331.120 ;
        RECT 1249.460 324.060 1249.720 324.320 ;
        RECT 1249.460 282.580 1249.720 282.840 ;
        RECT 1249.460 255.720 1249.720 255.980 ;
        RECT 1249.460 234.980 1249.720 235.240 ;
        RECT 1249.460 234.300 1249.720 234.560 ;
        RECT 1249.460 186.360 1249.720 186.620 ;
        RECT 1249.460 144.880 1249.720 145.140 ;
        RECT 1249.920 144.880 1250.180 145.140 ;
        RECT 1249.920 48.320 1250.180 48.580 ;
        RECT 1250.380 48.320 1250.640 48.580 ;
        RECT 204.800 39.820 205.060 40.080 ;
        RECT 1249.920 39.820 1250.180 40.080 ;
      LAYER met2 ;
        RECT 1253.980 1700.410 1254.260 1704.000 ;
        RECT 1251.820 1700.270 1254.260 1700.410 ;
        RECT 1251.820 1678.650 1251.960 1700.270 ;
        RECT 1253.980 1700.000 1254.260 1700.270 ;
        RECT 1249.980 1678.510 1251.960 1678.650 ;
        RECT 1249.980 1608.530 1250.120 1678.510 ;
        RECT 1249.920 1608.210 1250.180 1608.530 ;
        RECT 1249.920 1587.130 1250.180 1587.450 ;
        RECT 1249.980 1586.850 1250.120 1587.130 ;
        RECT 1249.980 1586.710 1250.580 1586.850 ;
        RECT 1250.440 1562.970 1250.580 1586.710 ;
        RECT 1249.460 1562.650 1249.720 1562.970 ;
        RECT 1250.380 1562.650 1250.640 1562.970 ;
        RECT 1249.520 1521.570 1249.660 1562.650 ;
        RECT 1249.520 1521.430 1250.120 1521.570 ;
        RECT 1249.980 1497.350 1250.120 1521.430 ;
        RECT 1249.920 1497.030 1250.180 1497.350 ;
        RECT 1249.920 1449.090 1250.180 1449.410 ;
        RECT 1249.980 1365.430 1250.120 1449.090 ;
        RECT 1249.920 1365.110 1250.180 1365.430 ;
        RECT 1249.920 1364.430 1250.180 1364.750 ;
        RECT 1249.980 1268.870 1250.120 1364.430 ;
        RECT 1249.920 1268.550 1250.180 1268.870 ;
        RECT 1249.920 1267.870 1250.180 1268.190 ;
        RECT 1249.980 882.630 1250.120 1267.870 ;
        RECT 1249.920 882.310 1250.180 882.630 ;
        RECT 1249.920 881.630 1250.180 881.950 ;
        RECT 1249.980 786.490 1250.120 881.630 ;
        RECT 1249.520 786.350 1250.120 786.490 ;
        RECT 1249.520 785.130 1249.660 786.350 ;
        RECT 1249.520 784.990 1250.120 785.130 ;
        RECT 1249.980 677.010 1250.120 784.990 ;
        RECT 1249.520 676.870 1250.120 677.010 ;
        RECT 1249.520 676.330 1249.660 676.870 ;
        RECT 1249.520 676.190 1250.120 676.330 ;
        RECT 1249.980 629.525 1250.120 676.190 ;
        RECT 1249.910 629.155 1250.190 629.525 ;
        RECT 1249.910 627.795 1250.190 628.165 ;
        RECT 1249.980 620.830 1250.120 627.795 ;
        RECT 1249.920 620.510 1250.180 620.830 ;
        RECT 1249.920 572.570 1250.180 572.890 ;
        RECT 1249.980 427.710 1250.120 572.570 ;
        RECT 1249.920 427.390 1250.180 427.710 ;
        RECT 1249.920 396.450 1250.180 396.770 ;
        RECT 1249.980 331.150 1250.120 396.450 ;
        RECT 1249.460 330.830 1249.720 331.150 ;
        RECT 1249.920 330.830 1250.180 331.150 ;
        RECT 1249.520 324.350 1249.660 330.830 ;
        RECT 1249.460 324.030 1249.720 324.350 ;
        RECT 1249.460 282.550 1249.720 282.870 ;
        RECT 1249.520 256.010 1249.660 282.550 ;
        RECT 1249.460 255.690 1249.720 256.010 ;
        RECT 1249.460 234.950 1249.720 235.270 ;
        RECT 1249.520 234.590 1249.660 234.950 ;
        RECT 1249.460 234.270 1249.720 234.590 ;
        RECT 1249.460 186.330 1249.720 186.650 ;
        RECT 1249.520 145.170 1249.660 186.330 ;
        RECT 1249.460 144.850 1249.720 145.170 ;
        RECT 1249.920 144.850 1250.180 145.170 ;
        RECT 1249.980 144.570 1250.120 144.850 ;
        RECT 1249.980 144.430 1250.580 144.570 ;
        RECT 1250.440 96.800 1250.580 144.430 ;
        RECT 1250.440 96.660 1251.040 96.800 ;
        RECT 1250.900 95.610 1251.040 96.660 ;
        RECT 1250.440 95.470 1251.040 95.610 ;
        RECT 1250.440 48.610 1250.580 95.470 ;
        RECT 1249.920 48.290 1250.180 48.610 ;
        RECT 1250.380 48.290 1250.640 48.610 ;
        RECT 1249.980 40.110 1250.120 48.290 ;
        RECT 204.800 39.790 205.060 40.110 ;
        RECT 1249.920 39.790 1250.180 40.110 ;
        RECT 204.860 2.400 205.000 39.790 ;
        RECT 204.650 -4.800 205.210 2.400 ;
      LAYER via2 ;
        RECT 1249.910 629.200 1250.190 629.480 ;
        RECT 1249.910 627.840 1250.190 628.120 ;
      LAYER met3 ;
        RECT 1249.885 629.500 1250.215 629.505 ;
        RECT 1249.630 629.490 1250.215 629.500 ;
        RECT 1249.430 629.190 1250.215 629.490 ;
        RECT 1249.630 629.180 1250.215 629.190 ;
        RECT 1249.885 629.175 1250.215 629.180 ;
        RECT 1249.885 628.140 1250.215 628.145 ;
        RECT 1249.630 628.130 1250.215 628.140 ;
        RECT 1249.630 627.830 1250.440 628.130 ;
        RECT 1249.630 627.820 1250.215 627.830 ;
        RECT 1249.885 627.815 1250.215 627.820 ;
      LAYER via3 ;
        RECT 1249.660 629.180 1249.980 629.500 ;
        RECT 1249.660 627.820 1249.980 628.140 ;
      LAYER met4 ;
        RECT 1249.655 629.175 1249.985 629.505 ;
        RECT 1249.670 628.145 1249.970 629.175 ;
        RECT 1249.655 627.815 1249.985 628.145 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 222.710 40.360 223.030 40.420 ;
        RECT 1263.230 40.360 1263.550 40.420 ;
        RECT 222.710 40.220 1263.550 40.360 ;
        RECT 222.710 40.160 223.030 40.220 ;
        RECT 1263.230 40.160 1263.550 40.220 ;
      LAYER via ;
        RECT 222.740 40.160 223.000 40.420 ;
        RECT 1263.260 40.160 1263.520 40.420 ;
      LAYER met2 ;
        RECT 1263.180 1700.000 1263.460 1704.000 ;
        RECT 1263.320 40.450 1263.460 1700.000 ;
        RECT 222.740 40.130 223.000 40.450 ;
        RECT 1263.260 40.130 1263.520 40.450 ;
        RECT 222.800 2.400 222.940 40.130 ;
        RECT 222.590 -4.800 223.150 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1153.290 1678.140 1153.610 1678.200 ;
        RECT 1157.430 1678.140 1157.750 1678.200 ;
        RECT 1153.290 1678.000 1157.750 1678.140 ;
        RECT 1153.290 1677.940 1153.610 1678.000 ;
        RECT 1157.430 1677.940 1157.750 1678.000 ;
        RECT 20.310 37.980 20.630 38.040 ;
        RECT 1153.290 37.980 1153.610 38.040 ;
        RECT 20.310 37.840 1153.610 37.980 ;
        RECT 20.310 37.780 20.630 37.840 ;
        RECT 1153.290 37.780 1153.610 37.840 ;
      LAYER via ;
        RECT 1153.320 1677.940 1153.580 1678.200 ;
        RECT 1157.460 1677.940 1157.720 1678.200 ;
        RECT 20.340 37.780 20.600 38.040 ;
        RECT 1153.320 37.780 1153.580 38.040 ;
      LAYER met2 ;
        RECT 1158.760 1700.410 1159.040 1704.000 ;
        RECT 1157.520 1700.270 1159.040 1700.410 ;
        RECT 1157.520 1678.230 1157.660 1700.270 ;
        RECT 1158.760 1700.000 1159.040 1700.270 ;
        RECT 1153.320 1677.910 1153.580 1678.230 ;
        RECT 1157.460 1677.910 1157.720 1678.230 ;
        RECT 1153.380 38.070 1153.520 1677.910 ;
        RECT 20.340 37.750 20.600 38.070 ;
        RECT 1153.320 37.750 1153.580 38.070 ;
        RECT 20.400 2.400 20.540 37.750 ;
        RECT 20.190 -4.800 20.750 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1167.090 1594.160 1167.410 1594.220 ;
        RECT 1167.550 1594.160 1167.870 1594.220 ;
        RECT 1167.090 1594.020 1167.870 1594.160 ;
        RECT 1167.090 1593.960 1167.410 1594.020 ;
        RECT 1167.550 1593.960 1167.870 1594.020 ;
        RECT 1166.630 1511.200 1166.950 1511.260 ;
        RECT 1167.550 1511.200 1167.870 1511.260 ;
        RECT 1166.630 1511.060 1167.870 1511.200 ;
        RECT 1166.630 1511.000 1166.950 1511.060 ;
        RECT 1167.550 1511.000 1167.870 1511.060 ;
        RECT 1166.630 1414.640 1166.950 1414.700 ;
        RECT 1167.550 1414.640 1167.870 1414.700 ;
        RECT 1166.630 1414.500 1167.870 1414.640 ;
        RECT 1166.630 1414.440 1166.950 1414.500 ;
        RECT 1167.550 1414.440 1167.870 1414.500 ;
        RECT 1166.630 1318.080 1166.950 1318.140 ;
        RECT 1167.550 1318.080 1167.870 1318.140 ;
        RECT 1166.630 1317.940 1167.870 1318.080 ;
        RECT 1166.630 1317.880 1166.950 1317.940 ;
        RECT 1167.550 1317.880 1167.870 1317.940 ;
        RECT 1166.630 1221.520 1166.950 1221.580 ;
        RECT 1167.550 1221.520 1167.870 1221.580 ;
        RECT 1166.630 1221.380 1167.870 1221.520 ;
        RECT 1166.630 1221.320 1166.950 1221.380 ;
        RECT 1167.550 1221.320 1167.870 1221.380 ;
        RECT 1166.630 1124.960 1166.950 1125.020 ;
        RECT 1167.550 1124.960 1167.870 1125.020 ;
        RECT 1166.630 1124.820 1167.870 1124.960 ;
        RECT 1166.630 1124.760 1166.950 1124.820 ;
        RECT 1167.550 1124.760 1167.870 1124.820 ;
        RECT 1166.630 1028.400 1166.950 1028.460 ;
        RECT 1167.550 1028.400 1167.870 1028.460 ;
        RECT 1166.630 1028.260 1167.870 1028.400 ;
        RECT 1166.630 1028.200 1166.950 1028.260 ;
        RECT 1167.550 1028.200 1167.870 1028.260 ;
        RECT 1166.630 931.840 1166.950 931.900 ;
        RECT 1167.550 931.840 1167.870 931.900 ;
        RECT 1166.630 931.700 1167.870 931.840 ;
        RECT 1166.630 931.640 1166.950 931.700 ;
        RECT 1167.550 931.640 1167.870 931.700 ;
        RECT 1166.630 835.280 1166.950 835.340 ;
        RECT 1167.550 835.280 1167.870 835.340 ;
        RECT 1166.630 835.140 1167.870 835.280 ;
        RECT 1166.630 835.080 1166.950 835.140 ;
        RECT 1167.550 835.080 1167.870 835.140 ;
        RECT 1166.630 738.380 1166.950 738.440 ;
        RECT 1167.550 738.380 1167.870 738.440 ;
        RECT 1166.630 738.240 1167.870 738.380 ;
        RECT 1166.630 738.180 1166.950 738.240 ;
        RECT 1167.550 738.180 1167.870 738.240 ;
        RECT 1166.630 641.820 1166.950 641.880 ;
        RECT 1167.550 641.820 1167.870 641.880 ;
        RECT 1166.630 641.680 1167.870 641.820 ;
        RECT 1166.630 641.620 1166.950 641.680 ;
        RECT 1167.550 641.620 1167.870 641.680 ;
        RECT 1166.630 545.260 1166.950 545.320 ;
        RECT 1167.550 545.260 1167.870 545.320 ;
        RECT 1166.630 545.120 1167.870 545.260 ;
        RECT 1166.630 545.060 1166.950 545.120 ;
        RECT 1167.550 545.060 1167.870 545.120 ;
        RECT 1166.630 448.700 1166.950 448.760 ;
        RECT 1167.550 448.700 1167.870 448.760 ;
        RECT 1166.630 448.560 1167.870 448.700 ;
        RECT 1166.630 448.500 1166.950 448.560 ;
        RECT 1167.550 448.500 1167.870 448.560 ;
        RECT 1167.090 241.640 1167.410 241.700 ;
        RECT 1167.550 241.640 1167.870 241.700 ;
        RECT 1167.090 241.500 1167.870 241.640 ;
        RECT 1167.090 241.440 1167.410 241.500 ;
        RECT 1167.550 241.440 1167.870 241.500 ;
        RECT 44.230 38.320 44.550 38.380 ;
        RECT 1166.630 38.320 1166.950 38.380 ;
        RECT 44.230 38.180 1166.950 38.320 ;
        RECT 44.230 38.120 44.550 38.180 ;
        RECT 1166.630 38.120 1166.950 38.180 ;
      LAYER via ;
        RECT 1167.120 1593.960 1167.380 1594.220 ;
        RECT 1167.580 1593.960 1167.840 1594.220 ;
        RECT 1166.660 1511.000 1166.920 1511.260 ;
        RECT 1167.580 1511.000 1167.840 1511.260 ;
        RECT 1166.660 1414.440 1166.920 1414.700 ;
        RECT 1167.580 1414.440 1167.840 1414.700 ;
        RECT 1166.660 1317.880 1166.920 1318.140 ;
        RECT 1167.580 1317.880 1167.840 1318.140 ;
        RECT 1166.660 1221.320 1166.920 1221.580 ;
        RECT 1167.580 1221.320 1167.840 1221.580 ;
        RECT 1166.660 1124.760 1166.920 1125.020 ;
        RECT 1167.580 1124.760 1167.840 1125.020 ;
        RECT 1166.660 1028.200 1166.920 1028.460 ;
        RECT 1167.580 1028.200 1167.840 1028.460 ;
        RECT 1166.660 931.640 1166.920 931.900 ;
        RECT 1167.580 931.640 1167.840 931.900 ;
        RECT 1166.660 835.080 1166.920 835.340 ;
        RECT 1167.580 835.080 1167.840 835.340 ;
        RECT 1166.660 738.180 1166.920 738.440 ;
        RECT 1167.580 738.180 1167.840 738.440 ;
        RECT 1166.660 641.620 1166.920 641.880 ;
        RECT 1167.580 641.620 1167.840 641.880 ;
        RECT 1166.660 545.060 1166.920 545.320 ;
        RECT 1167.580 545.060 1167.840 545.320 ;
        RECT 1166.660 448.500 1166.920 448.760 ;
        RECT 1167.580 448.500 1167.840 448.760 ;
        RECT 1167.120 241.440 1167.380 241.700 ;
        RECT 1167.580 241.440 1167.840 241.700 ;
        RECT 44.260 38.120 44.520 38.380 ;
        RECT 1166.660 38.120 1166.920 38.380 ;
      LAYER met2 ;
        RECT 1171.180 1700.410 1171.460 1704.000 ;
        RECT 1169.020 1700.270 1171.460 1700.410 ;
        RECT 1169.020 1677.970 1169.160 1700.270 ;
        RECT 1171.180 1700.000 1171.460 1700.270 ;
        RECT 1167.640 1677.830 1169.160 1677.970 ;
        RECT 1167.640 1594.250 1167.780 1677.830 ;
        RECT 1167.120 1593.930 1167.380 1594.250 ;
        RECT 1167.580 1593.930 1167.840 1594.250 ;
        RECT 1167.180 1593.650 1167.320 1593.930 ;
        RECT 1167.180 1593.510 1167.780 1593.650 ;
        RECT 1167.640 1511.290 1167.780 1593.510 ;
        RECT 1166.660 1510.970 1166.920 1511.290 ;
        RECT 1167.580 1510.970 1167.840 1511.290 ;
        RECT 1166.720 1510.690 1166.860 1510.970 ;
        RECT 1166.720 1510.550 1167.320 1510.690 ;
        RECT 1167.180 1463.090 1167.320 1510.550 ;
        RECT 1167.180 1462.950 1167.780 1463.090 ;
        RECT 1167.640 1414.730 1167.780 1462.950 ;
        RECT 1166.660 1414.410 1166.920 1414.730 ;
        RECT 1167.580 1414.410 1167.840 1414.730 ;
        RECT 1166.720 1414.130 1166.860 1414.410 ;
        RECT 1166.720 1413.990 1167.320 1414.130 ;
        RECT 1167.180 1366.530 1167.320 1413.990 ;
        RECT 1167.180 1366.390 1167.780 1366.530 ;
        RECT 1167.640 1318.170 1167.780 1366.390 ;
        RECT 1166.660 1317.850 1166.920 1318.170 ;
        RECT 1167.580 1317.850 1167.840 1318.170 ;
        RECT 1166.720 1317.570 1166.860 1317.850 ;
        RECT 1166.720 1317.430 1167.320 1317.570 ;
        RECT 1167.180 1269.970 1167.320 1317.430 ;
        RECT 1167.180 1269.830 1167.780 1269.970 ;
        RECT 1167.640 1221.610 1167.780 1269.830 ;
        RECT 1166.660 1221.290 1166.920 1221.610 ;
        RECT 1167.580 1221.290 1167.840 1221.610 ;
        RECT 1166.720 1221.010 1166.860 1221.290 ;
        RECT 1166.720 1220.870 1167.320 1221.010 ;
        RECT 1167.180 1173.410 1167.320 1220.870 ;
        RECT 1167.180 1173.270 1167.780 1173.410 ;
        RECT 1167.640 1125.050 1167.780 1173.270 ;
        RECT 1166.660 1124.730 1166.920 1125.050 ;
        RECT 1167.580 1124.730 1167.840 1125.050 ;
        RECT 1166.720 1124.450 1166.860 1124.730 ;
        RECT 1166.720 1124.310 1167.320 1124.450 ;
        RECT 1167.180 1076.850 1167.320 1124.310 ;
        RECT 1167.180 1076.710 1167.780 1076.850 ;
        RECT 1167.640 1028.490 1167.780 1076.710 ;
        RECT 1166.660 1028.170 1166.920 1028.490 ;
        RECT 1167.580 1028.170 1167.840 1028.490 ;
        RECT 1166.720 1027.890 1166.860 1028.170 ;
        RECT 1166.720 1027.750 1167.320 1027.890 ;
        RECT 1167.180 980.290 1167.320 1027.750 ;
        RECT 1167.180 980.150 1167.780 980.290 ;
        RECT 1167.640 931.930 1167.780 980.150 ;
        RECT 1166.660 931.610 1166.920 931.930 ;
        RECT 1167.580 931.610 1167.840 931.930 ;
        RECT 1166.720 883.050 1166.860 931.610 ;
        RECT 1166.720 882.910 1167.780 883.050 ;
        RECT 1167.640 835.370 1167.780 882.910 ;
        RECT 1166.660 835.050 1166.920 835.370 ;
        RECT 1167.580 835.050 1167.840 835.370 ;
        RECT 1166.720 786.490 1166.860 835.050 ;
        RECT 1166.720 786.350 1167.780 786.490 ;
        RECT 1167.640 738.470 1167.780 786.350 ;
        RECT 1166.660 738.150 1166.920 738.470 ;
        RECT 1167.580 738.150 1167.840 738.470 ;
        RECT 1166.720 689.930 1166.860 738.150 ;
        RECT 1166.720 689.790 1167.780 689.930 ;
        RECT 1167.640 641.910 1167.780 689.790 ;
        RECT 1166.660 641.590 1166.920 641.910 ;
        RECT 1167.580 641.590 1167.840 641.910 ;
        RECT 1166.720 593.370 1166.860 641.590 ;
        RECT 1166.720 593.230 1167.780 593.370 ;
        RECT 1167.640 545.350 1167.780 593.230 ;
        RECT 1166.660 545.030 1166.920 545.350 ;
        RECT 1167.580 545.030 1167.840 545.350 ;
        RECT 1166.720 496.810 1166.860 545.030 ;
        RECT 1166.720 496.670 1167.780 496.810 ;
        RECT 1167.640 448.790 1167.780 496.670 ;
        RECT 1166.660 448.470 1166.920 448.790 ;
        RECT 1167.580 448.470 1167.840 448.790 ;
        RECT 1166.720 400.250 1166.860 448.470 ;
        RECT 1166.720 400.110 1167.780 400.250 ;
        RECT 1167.640 241.730 1167.780 400.110 ;
        RECT 1167.120 241.410 1167.380 241.730 ;
        RECT 1167.580 241.410 1167.840 241.730 ;
        RECT 1167.180 207.130 1167.320 241.410 ;
        RECT 1167.180 206.990 1167.780 207.130 ;
        RECT 1167.640 158.850 1167.780 206.990 ;
        RECT 1166.720 158.710 1167.780 158.850 ;
        RECT 1166.720 158.170 1166.860 158.710 ;
        RECT 1166.720 158.030 1167.320 158.170 ;
        RECT 1167.180 41.720 1167.320 158.030 ;
        RECT 1166.720 41.580 1167.320 41.720 ;
        RECT 1166.720 38.410 1166.860 41.580 ;
        RECT 44.260 38.090 44.520 38.410 ;
        RECT 1166.660 38.090 1166.920 38.410 ;
        RECT 44.320 2.400 44.460 38.090 ;
        RECT 44.110 -4.800 44.670 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1270.665 1386.945 1270.835 1448.995 ;
        RECT 1270.665 1242.445 1270.835 1270.155 ;
        RECT 1270.665 1221.025 1270.835 1241.935 ;
        RECT 1270.665 834.785 1270.835 862.495 ;
        RECT 1272.045 717.825 1272.215 765.595 ;
        RECT 1271.125 620.925 1271.295 717.655 ;
        RECT 1271.125 469.285 1271.295 517.395 ;
        RECT 1270.665 338.045 1270.835 427.635 ;
      LAYER mcon ;
        RECT 1270.665 1448.825 1270.835 1448.995 ;
        RECT 1270.665 1269.985 1270.835 1270.155 ;
        RECT 1270.665 1241.765 1270.835 1241.935 ;
        RECT 1270.665 862.325 1270.835 862.495 ;
        RECT 1272.045 765.425 1272.215 765.595 ;
        RECT 1271.125 717.485 1271.295 717.655 ;
        RECT 1271.125 517.225 1271.295 517.395 ;
        RECT 1270.665 427.465 1270.835 427.635 ;
      LAYER met1 ;
        RECT 1271.050 1652.300 1271.370 1652.360 ;
        RECT 1273.810 1652.300 1274.130 1652.360 ;
        RECT 1271.050 1652.160 1274.130 1652.300 ;
        RECT 1271.050 1652.100 1271.370 1652.160 ;
        RECT 1273.810 1652.100 1274.130 1652.160 ;
        RECT 1270.590 1448.980 1270.910 1449.040 ;
        RECT 1270.395 1448.840 1270.910 1448.980 ;
        RECT 1270.590 1448.780 1270.910 1448.840 ;
        RECT 1270.605 1387.100 1270.895 1387.145 ;
        RECT 1271.050 1387.100 1271.370 1387.160 ;
        RECT 1270.605 1386.960 1271.370 1387.100 ;
        RECT 1270.605 1386.915 1270.895 1386.960 ;
        RECT 1271.050 1386.900 1271.370 1386.960 ;
        RECT 1270.605 1270.140 1270.895 1270.185 ;
        RECT 1271.050 1270.140 1271.370 1270.200 ;
        RECT 1270.605 1270.000 1271.370 1270.140 ;
        RECT 1270.605 1269.955 1270.895 1270.000 ;
        RECT 1271.050 1269.940 1271.370 1270.000 ;
        RECT 1270.590 1242.600 1270.910 1242.660 ;
        RECT 1270.395 1242.460 1270.910 1242.600 ;
        RECT 1270.590 1242.400 1270.910 1242.460 ;
        RECT 1270.590 1241.920 1270.910 1241.980 ;
        RECT 1270.395 1241.780 1270.910 1241.920 ;
        RECT 1270.590 1241.720 1270.910 1241.780 ;
        RECT 1270.590 1221.180 1270.910 1221.240 ;
        RECT 1270.395 1221.040 1270.910 1221.180 ;
        RECT 1270.590 1220.980 1270.910 1221.040 ;
        RECT 1271.050 1063.080 1271.370 1063.140 ;
        RECT 1270.680 1062.940 1271.370 1063.080 ;
        RECT 1270.680 1062.800 1270.820 1062.940 ;
        RECT 1271.050 1062.880 1271.370 1062.940 ;
        RECT 1270.590 1062.540 1270.910 1062.800 ;
        RECT 1270.590 869.620 1270.910 869.680 ;
        RECT 1271.510 869.620 1271.830 869.680 ;
        RECT 1270.590 869.480 1271.830 869.620 ;
        RECT 1270.590 869.420 1270.910 869.480 ;
        RECT 1271.510 869.420 1271.830 869.480 ;
        RECT 1270.590 862.480 1270.910 862.540 ;
        RECT 1270.395 862.340 1270.910 862.480 ;
        RECT 1270.590 862.280 1270.910 862.340 ;
        RECT 1270.590 834.940 1270.910 835.000 ;
        RECT 1270.395 834.800 1270.910 834.940 ;
        RECT 1270.590 834.740 1270.910 834.800 ;
        RECT 1270.590 766.260 1270.910 766.320 ;
        RECT 1271.970 766.260 1272.290 766.320 ;
        RECT 1270.590 766.120 1272.290 766.260 ;
        RECT 1270.590 766.060 1270.910 766.120 ;
        RECT 1271.970 766.060 1272.290 766.120 ;
        RECT 1271.970 765.580 1272.290 765.640 ;
        RECT 1271.775 765.440 1272.290 765.580 ;
        RECT 1271.970 765.380 1272.290 765.440 ;
        RECT 1270.590 717.980 1270.910 718.040 ;
        RECT 1271.985 717.980 1272.275 718.025 ;
        RECT 1270.590 717.840 1272.275 717.980 ;
        RECT 1270.590 717.780 1270.910 717.840 ;
        RECT 1271.985 717.795 1272.275 717.840 ;
        RECT 1271.050 717.640 1271.370 717.700 ;
        RECT 1270.855 717.500 1271.370 717.640 ;
        RECT 1271.050 717.440 1271.370 717.500 ;
        RECT 1271.050 621.080 1271.370 621.140 ;
        RECT 1270.855 620.940 1271.370 621.080 ;
        RECT 1271.050 620.880 1271.370 620.940 ;
        RECT 1270.590 579.600 1270.910 579.660 ;
        RECT 1271.050 579.600 1271.370 579.660 ;
        RECT 1270.590 579.460 1271.370 579.600 ;
        RECT 1270.590 579.400 1270.910 579.460 ;
        RECT 1271.050 579.400 1271.370 579.460 ;
        RECT 1270.590 572.460 1270.910 572.520 ;
        RECT 1271.050 572.460 1271.370 572.520 ;
        RECT 1270.590 572.320 1271.370 572.460 ;
        RECT 1270.590 572.260 1270.910 572.320 ;
        RECT 1271.050 572.260 1271.370 572.320 ;
        RECT 1271.050 517.380 1271.370 517.440 ;
        RECT 1270.855 517.240 1271.370 517.380 ;
        RECT 1271.050 517.180 1271.370 517.240 ;
        RECT 1271.050 469.440 1271.370 469.500 ;
        RECT 1270.855 469.300 1271.370 469.440 ;
        RECT 1271.050 469.240 1271.370 469.300 ;
        RECT 1270.605 427.620 1270.895 427.665 ;
        RECT 1271.050 427.620 1271.370 427.680 ;
        RECT 1270.605 427.480 1271.370 427.620 ;
        RECT 1270.605 427.435 1270.895 427.480 ;
        RECT 1271.050 427.420 1271.370 427.480 ;
        RECT 1270.590 338.200 1270.910 338.260 ;
        RECT 1270.395 338.060 1270.910 338.200 ;
        RECT 1270.590 338.000 1270.910 338.060 ;
        RECT 1271.050 144.740 1271.370 144.800 ;
        RECT 1271.510 144.740 1271.830 144.800 ;
        RECT 1271.050 144.600 1271.830 144.740 ;
        RECT 1271.050 144.540 1271.370 144.600 ;
        RECT 1271.510 144.540 1271.830 144.600 ;
        RECT 1271.510 96.260 1271.830 96.520 ;
        RECT 1271.600 95.840 1271.740 96.260 ;
        RECT 1271.510 95.580 1271.830 95.840 ;
        RECT 1270.130 48.520 1270.450 48.580 ;
        RECT 1271.510 48.520 1271.830 48.580 ;
        RECT 1270.130 48.380 1271.830 48.520 ;
        RECT 1270.130 48.320 1270.450 48.380 ;
        RECT 1271.510 48.320 1271.830 48.380 ;
        RECT 246.630 40.700 246.950 40.760 ;
        RECT 1270.130 40.700 1270.450 40.760 ;
        RECT 246.630 40.560 1270.450 40.700 ;
        RECT 246.630 40.500 246.950 40.560 ;
        RECT 1270.130 40.500 1270.450 40.560 ;
      LAYER via ;
        RECT 1271.080 1652.100 1271.340 1652.360 ;
        RECT 1273.840 1652.100 1274.100 1652.360 ;
        RECT 1270.620 1448.780 1270.880 1449.040 ;
        RECT 1271.080 1386.900 1271.340 1387.160 ;
        RECT 1271.080 1269.940 1271.340 1270.200 ;
        RECT 1270.620 1242.400 1270.880 1242.660 ;
        RECT 1270.620 1241.720 1270.880 1241.980 ;
        RECT 1270.620 1220.980 1270.880 1221.240 ;
        RECT 1271.080 1062.880 1271.340 1063.140 ;
        RECT 1270.620 1062.540 1270.880 1062.800 ;
        RECT 1270.620 869.420 1270.880 869.680 ;
        RECT 1271.540 869.420 1271.800 869.680 ;
        RECT 1270.620 862.280 1270.880 862.540 ;
        RECT 1270.620 834.740 1270.880 835.000 ;
        RECT 1270.620 766.060 1270.880 766.320 ;
        RECT 1272.000 766.060 1272.260 766.320 ;
        RECT 1272.000 765.380 1272.260 765.640 ;
        RECT 1270.620 717.780 1270.880 718.040 ;
        RECT 1271.080 717.440 1271.340 717.700 ;
        RECT 1271.080 620.880 1271.340 621.140 ;
        RECT 1270.620 579.400 1270.880 579.660 ;
        RECT 1271.080 579.400 1271.340 579.660 ;
        RECT 1270.620 572.260 1270.880 572.520 ;
        RECT 1271.080 572.260 1271.340 572.520 ;
        RECT 1271.080 517.180 1271.340 517.440 ;
        RECT 1271.080 469.240 1271.340 469.500 ;
        RECT 1271.080 427.420 1271.340 427.680 ;
        RECT 1270.620 338.000 1270.880 338.260 ;
        RECT 1271.080 144.540 1271.340 144.800 ;
        RECT 1271.540 144.540 1271.800 144.800 ;
        RECT 1271.540 96.260 1271.800 96.520 ;
        RECT 1271.540 95.580 1271.800 95.840 ;
        RECT 1270.160 48.320 1270.420 48.580 ;
        RECT 1271.540 48.320 1271.800 48.580 ;
        RECT 246.660 40.500 246.920 40.760 ;
        RECT 1270.160 40.500 1270.420 40.760 ;
      LAYER met2 ;
        RECT 1275.140 1700.410 1275.420 1704.000 ;
        RECT 1273.900 1700.270 1275.420 1700.410 ;
        RECT 1273.900 1652.390 1274.040 1700.270 ;
        RECT 1275.140 1700.000 1275.420 1700.270 ;
        RECT 1271.080 1652.070 1271.340 1652.390 ;
        RECT 1273.840 1652.070 1274.100 1652.390 ;
        RECT 1271.140 1608.610 1271.280 1652.070 ;
        RECT 1271.140 1608.470 1271.740 1608.610 ;
        RECT 1271.600 1607.250 1271.740 1608.470 ;
        RECT 1270.680 1607.110 1271.740 1607.250 ;
        RECT 1270.680 1593.650 1270.820 1607.110 ;
        RECT 1270.680 1593.510 1271.280 1593.650 ;
        RECT 1271.140 1463.090 1271.280 1593.510 ;
        RECT 1270.680 1462.950 1271.280 1463.090 ;
        RECT 1270.680 1449.070 1270.820 1462.950 ;
        RECT 1270.620 1448.750 1270.880 1449.070 ;
        RECT 1271.080 1386.870 1271.340 1387.190 ;
        RECT 1271.140 1338.765 1271.280 1386.870 ;
        RECT 1270.150 1338.395 1270.430 1338.765 ;
        RECT 1271.070 1338.395 1271.350 1338.765 ;
        RECT 1270.220 1290.485 1270.360 1338.395 ;
        RECT 1270.150 1290.115 1270.430 1290.485 ;
        RECT 1271.070 1290.115 1271.350 1290.485 ;
        RECT 1271.140 1270.230 1271.280 1290.115 ;
        RECT 1271.080 1269.910 1271.340 1270.230 ;
        RECT 1270.620 1242.370 1270.880 1242.690 ;
        RECT 1270.680 1242.010 1270.820 1242.370 ;
        RECT 1270.620 1241.690 1270.880 1242.010 ;
        RECT 1270.620 1220.950 1270.880 1221.270 ;
        RECT 1270.680 1193.810 1270.820 1220.950 ;
        RECT 1270.680 1193.670 1271.280 1193.810 ;
        RECT 1271.140 1063.170 1271.280 1193.670 ;
        RECT 1271.080 1062.850 1271.340 1063.170 ;
        RECT 1270.620 1062.510 1270.880 1062.830 ;
        RECT 1270.680 1038.770 1270.820 1062.510 ;
        RECT 1270.680 1038.630 1271.280 1038.770 ;
        RECT 1271.140 990.490 1271.280 1038.630 ;
        RECT 1270.680 990.350 1271.280 990.490 ;
        RECT 1270.680 966.125 1270.820 990.350 ;
        RECT 1270.610 965.755 1270.890 966.125 ;
        RECT 1271.530 965.755 1271.810 966.125 ;
        RECT 1271.600 869.710 1271.740 965.755 ;
        RECT 1270.620 869.390 1270.880 869.710 ;
        RECT 1271.540 869.390 1271.800 869.710 ;
        RECT 1270.680 862.570 1270.820 869.390 ;
        RECT 1270.620 862.250 1270.880 862.570 ;
        RECT 1270.620 834.710 1270.880 835.030 ;
        RECT 1270.680 766.350 1270.820 834.710 ;
        RECT 1270.620 766.030 1270.880 766.350 ;
        RECT 1272.000 766.030 1272.260 766.350 ;
        RECT 1272.060 765.670 1272.200 766.030 ;
        RECT 1272.000 765.350 1272.260 765.670 ;
        RECT 1270.620 717.810 1270.880 718.070 ;
        RECT 1270.620 717.750 1271.280 717.810 ;
        RECT 1270.680 717.730 1271.280 717.750 ;
        RECT 1270.680 717.670 1271.340 717.730 ;
        RECT 1271.080 717.410 1271.340 717.670 ;
        RECT 1271.080 620.850 1271.340 621.170 ;
        RECT 1271.140 579.770 1271.280 620.850 ;
        RECT 1270.680 579.690 1271.280 579.770 ;
        RECT 1270.620 579.630 1271.340 579.690 ;
        RECT 1270.620 579.370 1270.880 579.630 ;
        RECT 1271.080 579.370 1271.340 579.630 ;
        RECT 1270.680 579.215 1270.820 579.370 ;
        RECT 1271.140 572.550 1271.280 579.370 ;
        RECT 1270.620 572.230 1270.880 572.550 ;
        RECT 1271.080 572.230 1271.340 572.550 ;
        RECT 1270.680 524.690 1270.820 572.230 ;
        RECT 1270.680 524.550 1271.280 524.690 ;
        RECT 1271.140 517.470 1271.280 524.550 ;
        RECT 1271.080 517.150 1271.340 517.470 ;
        RECT 1271.080 469.210 1271.340 469.530 ;
        RECT 1271.140 427.710 1271.280 469.210 ;
        RECT 1271.080 427.390 1271.340 427.710 ;
        RECT 1270.620 337.970 1270.880 338.290 ;
        RECT 1270.680 304.370 1270.820 337.970 ;
        RECT 1270.680 304.230 1271.280 304.370 ;
        RECT 1271.140 303.520 1271.280 304.230 ;
        RECT 1270.680 303.380 1271.280 303.520 ;
        RECT 1270.680 265.610 1270.820 303.380 ;
        RECT 1270.680 265.470 1271.280 265.610 ;
        RECT 1271.140 144.830 1271.280 265.470 ;
        RECT 1271.080 144.510 1271.340 144.830 ;
        RECT 1271.540 144.510 1271.800 144.830 ;
        RECT 1271.600 96.550 1271.740 144.510 ;
        RECT 1271.540 96.230 1271.800 96.550 ;
        RECT 1271.540 95.550 1271.800 95.870 ;
        RECT 1271.600 48.610 1271.740 95.550 ;
        RECT 1270.160 48.290 1270.420 48.610 ;
        RECT 1271.540 48.290 1271.800 48.610 ;
        RECT 1270.220 40.790 1270.360 48.290 ;
        RECT 246.660 40.470 246.920 40.790 ;
        RECT 1270.160 40.470 1270.420 40.790 ;
        RECT 246.720 2.400 246.860 40.470 ;
        RECT 246.510 -4.800 247.070 2.400 ;
      LAYER via2 ;
        RECT 1270.150 1338.440 1270.430 1338.720 ;
        RECT 1271.070 1338.440 1271.350 1338.720 ;
        RECT 1270.150 1290.160 1270.430 1290.440 ;
        RECT 1271.070 1290.160 1271.350 1290.440 ;
        RECT 1270.610 965.800 1270.890 966.080 ;
        RECT 1271.530 965.800 1271.810 966.080 ;
      LAYER met3 ;
        RECT 1270.125 1338.730 1270.455 1338.745 ;
        RECT 1271.045 1338.730 1271.375 1338.745 ;
        RECT 1270.125 1338.430 1271.375 1338.730 ;
        RECT 1270.125 1338.415 1270.455 1338.430 ;
        RECT 1271.045 1338.415 1271.375 1338.430 ;
        RECT 1270.125 1290.450 1270.455 1290.465 ;
        RECT 1271.045 1290.450 1271.375 1290.465 ;
        RECT 1270.125 1290.150 1271.375 1290.450 ;
        RECT 1270.125 1290.135 1270.455 1290.150 ;
        RECT 1271.045 1290.135 1271.375 1290.150 ;
        RECT 1270.585 966.090 1270.915 966.105 ;
        RECT 1271.505 966.090 1271.835 966.105 ;
        RECT 1270.585 965.790 1271.835 966.090 ;
        RECT 1270.585 965.775 1270.915 965.790 ;
        RECT 1271.505 965.775 1271.835 965.790 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 264.110 41.040 264.430 41.100 ;
        RECT 1283.930 41.040 1284.250 41.100 ;
        RECT 264.110 40.900 1284.250 41.040 ;
        RECT 264.110 40.840 264.430 40.900 ;
        RECT 1283.930 40.840 1284.250 40.900 ;
      LAYER via ;
        RECT 264.140 40.840 264.400 41.100 ;
        RECT 1283.960 40.840 1284.220 41.100 ;
      LAYER met2 ;
        RECT 1284.340 1700.410 1284.620 1704.000 ;
        RECT 1284.020 1700.270 1284.620 1700.410 ;
        RECT 1284.020 41.130 1284.160 1700.270 ;
        RECT 1284.340 1700.000 1284.620 1700.270 ;
        RECT 264.140 40.810 264.400 41.130 ;
        RECT 1283.960 40.810 1284.220 41.130 ;
        RECT 264.200 2.400 264.340 40.810 ;
        RECT 263.990 -4.800 264.550 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 282.050 41.380 282.370 41.440 ;
        RECT 1291.750 41.380 1292.070 41.440 ;
        RECT 282.050 41.240 1292.070 41.380 ;
        RECT 282.050 41.180 282.370 41.240 ;
        RECT 1291.750 41.180 1292.070 41.240 ;
      LAYER via ;
        RECT 282.080 41.180 282.340 41.440 ;
        RECT 1291.780 41.180 1292.040 41.440 ;
      LAYER met2 ;
        RECT 1293.540 1700.410 1293.820 1704.000 ;
        RECT 1291.840 1700.270 1293.820 1700.410 ;
        RECT 1291.840 41.470 1291.980 1700.270 ;
        RECT 1293.540 1700.000 1293.820 1700.270 ;
        RECT 282.080 41.150 282.340 41.470 ;
        RECT 1291.780 41.150 1292.040 41.470 ;
        RECT 282.140 2.400 282.280 41.150 ;
        RECT 281.930 -4.800 282.490 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1298.265 1594.005 1298.435 1608.115 ;
        RECT 1298.265 1386.945 1298.435 1448.995 ;
        RECT 1298.265 1242.445 1298.435 1270.155 ;
        RECT 1298.265 1110.865 1298.435 1158.975 ;
        RECT 1298.265 1014.305 1298.435 1062.415 ;
        RECT 1298.265 814.385 1298.435 862.495 ;
        RECT 1298.265 668.865 1298.435 717.655 ;
        RECT 1298.265 355.385 1298.435 420.835 ;
      LAYER mcon ;
        RECT 1298.265 1607.945 1298.435 1608.115 ;
        RECT 1298.265 1448.825 1298.435 1448.995 ;
        RECT 1298.265 1269.985 1298.435 1270.155 ;
        RECT 1298.265 1158.805 1298.435 1158.975 ;
        RECT 1298.265 1062.245 1298.435 1062.415 ;
        RECT 1298.265 862.325 1298.435 862.495 ;
        RECT 1298.265 717.485 1298.435 717.655 ;
        RECT 1298.265 420.665 1298.435 420.835 ;
      LAYER met1 ;
        RECT 1298.190 1666.580 1298.510 1666.640 ;
        RECT 1301.410 1666.580 1301.730 1666.640 ;
        RECT 1298.190 1666.440 1301.730 1666.580 ;
        RECT 1298.190 1666.380 1298.510 1666.440 ;
        RECT 1301.410 1666.380 1301.730 1666.440 ;
        RECT 1298.190 1608.100 1298.510 1608.160 ;
        RECT 1297.995 1607.960 1298.510 1608.100 ;
        RECT 1298.190 1607.900 1298.510 1607.960 ;
        RECT 1298.190 1594.160 1298.510 1594.220 ;
        RECT 1297.995 1594.020 1298.510 1594.160 ;
        RECT 1298.190 1593.960 1298.510 1594.020 ;
        RECT 1298.190 1448.980 1298.510 1449.040 ;
        RECT 1297.995 1448.840 1298.510 1448.980 ;
        RECT 1298.190 1448.780 1298.510 1448.840 ;
        RECT 1298.205 1387.100 1298.495 1387.145 ;
        RECT 1298.650 1387.100 1298.970 1387.160 ;
        RECT 1298.205 1386.960 1298.970 1387.100 ;
        RECT 1298.205 1386.915 1298.495 1386.960 ;
        RECT 1298.650 1386.900 1298.970 1386.960 ;
        RECT 1298.205 1270.140 1298.495 1270.185 ;
        RECT 1298.650 1270.140 1298.970 1270.200 ;
        RECT 1298.205 1270.000 1298.970 1270.140 ;
        RECT 1298.205 1269.955 1298.495 1270.000 ;
        RECT 1298.650 1269.940 1298.970 1270.000 ;
        RECT 1298.190 1242.600 1298.510 1242.660 ;
        RECT 1297.995 1242.460 1298.510 1242.600 ;
        RECT 1298.190 1242.400 1298.510 1242.460 ;
        RECT 1296.810 1241.920 1297.130 1241.980 ;
        RECT 1298.190 1241.920 1298.510 1241.980 ;
        RECT 1296.810 1241.780 1298.510 1241.920 ;
        RECT 1296.810 1241.720 1297.130 1241.780 ;
        RECT 1298.190 1241.720 1298.510 1241.780 ;
        RECT 1298.190 1158.960 1298.510 1159.020 ;
        RECT 1297.995 1158.820 1298.510 1158.960 ;
        RECT 1298.190 1158.760 1298.510 1158.820 ;
        RECT 1298.205 1111.020 1298.495 1111.065 ;
        RECT 1298.650 1111.020 1298.970 1111.080 ;
        RECT 1298.205 1110.880 1298.970 1111.020 ;
        RECT 1298.205 1110.835 1298.495 1110.880 ;
        RECT 1298.650 1110.820 1298.970 1110.880 ;
        RECT 1298.650 1087.220 1298.970 1087.280 ;
        RECT 1298.280 1087.080 1298.970 1087.220 ;
        RECT 1298.280 1086.940 1298.420 1087.080 ;
        RECT 1298.650 1087.020 1298.970 1087.080 ;
        RECT 1298.190 1086.680 1298.510 1086.940 ;
        RECT 1298.190 1062.400 1298.510 1062.460 ;
        RECT 1297.995 1062.260 1298.510 1062.400 ;
        RECT 1298.190 1062.200 1298.510 1062.260 ;
        RECT 1298.205 1014.460 1298.495 1014.505 ;
        RECT 1298.650 1014.460 1298.970 1014.520 ;
        RECT 1298.205 1014.320 1298.970 1014.460 ;
        RECT 1298.205 1014.275 1298.495 1014.320 ;
        RECT 1298.650 1014.260 1298.970 1014.320 ;
        RECT 1298.650 990.660 1298.970 990.720 ;
        RECT 1298.280 990.520 1298.970 990.660 ;
        RECT 1298.280 990.380 1298.420 990.520 ;
        RECT 1298.650 990.460 1298.970 990.520 ;
        RECT 1298.190 990.120 1298.510 990.380 ;
        RECT 1298.650 869.620 1298.970 869.680 ;
        RECT 1299.110 869.620 1299.430 869.680 ;
        RECT 1298.650 869.480 1299.430 869.620 ;
        RECT 1298.650 869.420 1298.970 869.480 ;
        RECT 1299.110 869.420 1299.430 869.480 ;
        RECT 1298.205 862.480 1298.495 862.525 ;
        RECT 1298.650 862.480 1298.970 862.540 ;
        RECT 1298.205 862.340 1298.970 862.480 ;
        RECT 1298.205 862.295 1298.495 862.340 ;
        RECT 1298.650 862.280 1298.970 862.340 ;
        RECT 1298.190 814.540 1298.510 814.600 ;
        RECT 1297.995 814.400 1298.510 814.540 ;
        RECT 1298.190 814.340 1298.510 814.400 ;
        RECT 1298.205 717.640 1298.495 717.685 ;
        RECT 1298.650 717.640 1298.970 717.700 ;
        RECT 1298.205 717.500 1298.970 717.640 ;
        RECT 1298.205 717.455 1298.495 717.500 ;
        RECT 1298.650 717.440 1298.970 717.500 ;
        RECT 1298.205 669.020 1298.495 669.065 ;
        RECT 1298.650 669.020 1298.970 669.080 ;
        RECT 1298.205 668.880 1298.970 669.020 ;
        RECT 1298.205 668.835 1298.495 668.880 ;
        RECT 1298.650 668.820 1298.970 668.880 ;
        RECT 1298.650 621.560 1298.970 621.820 ;
        RECT 1298.740 621.140 1298.880 621.560 ;
        RECT 1298.650 620.880 1298.970 621.140 ;
        RECT 1298.650 613.940 1298.970 614.000 ;
        RECT 1299.110 613.940 1299.430 614.000 ;
        RECT 1298.650 613.800 1299.430 613.940 ;
        RECT 1298.650 613.740 1298.970 613.800 ;
        RECT 1299.110 613.740 1299.430 613.800 ;
        RECT 1298.190 476.240 1298.510 476.300 ;
        RECT 1299.110 476.240 1299.430 476.300 ;
        RECT 1298.190 476.100 1299.430 476.240 ;
        RECT 1298.190 476.040 1298.510 476.100 ;
        RECT 1299.110 476.040 1299.430 476.100 ;
        RECT 1298.190 448.500 1298.510 448.760 ;
        RECT 1298.280 448.020 1298.420 448.500 ;
        RECT 1298.650 448.020 1298.970 448.080 ;
        RECT 1298.280 447.880 1298.970 448.020 ;
        RECT 1298.650 447.820 1298.970 447.880 ;
        RECT 1298.205 420.820 1298.495 420.865 ;
        RECT 1298.650 420.820 1298.970 420.880 ;
        RECT 1298.205 420.680 1298.970 420.820 ;
        RECT 1298.205 420.635 1298.495 420.680 ;
        RECT 1298.650 420.620 1298.970 420.680 ;
        RECT 1298.190 355.540 1298.510 355.600 ;
        RECT 1297.995 355.400 1298.510 355.540 ;
        RECT 1298.190 355.340 1298.510 355.400 ;
        RECT 1298.190 304.000 1298.510 304.260 ;
        RECT 1298.280 303.580 1298.420 304.000 ;
        RECT 1298.190 303.320 1298.510 303.580 ;
        RECT 1297.730 144.740 1298.050 144.800 ;
        RECT 1298.650 144.740 1298.970 144.800 ;
        RECT 1297.730 144.600 1298.970 144.740 ;
        RECT 1297.730 144.540 1298.050 144.600 ;
        RECT 1298.650 144.540 1298.970 144.600 ;
        RECT 299.990 16.900 300.310 16.960 ;
        RECT 303.210 16.900 303.530 16.960 ;
        RECT 299.990 16.760 303.530 16.900 ;
        RECT 299.990 16.700 300.310 16.760 ;
        RECT 303.210 16.700 303.530 16.760 ;
      LAYER via ;
        RECT 1298.220 1666.380 1298.480 1666.640 ;
        RECT 1301.440 1666.380 1301.700 1666.640 ;
        RECT 1298.220 1607.900 1298.480 1608.160 ;
        RECT 1298.220 1593.960 1298.480 1594.220 ;
        RECT 1298.220 1448.780 1298.480 1449.040 ;
        RECT 1298.680 1386.900 1298.940 1387.160 ;
        RECT 1298.680 1269.940 1298.940 1270.200 ;
        RECT 1298.220 1242.400 1298.480 1242.660 ;
        RECT 1296.840 1241.720 1297.100 1241.980 ;
        RECT 1298.220 1241.720 1298.480 1241.980 ;
        RECT 1298.220 1158.760 1298.480 1159.020 ;
        RECT 1298.680 1110.820 1298.940 1111.080 ;
        RECT 1298.680 1087.020 1298.940 1087.280 ;
        RECT 1298.220 1086.680 1298.480 1086.940 ;
        RECT 1298.220 1062.200 1298.480 1062.460 ;
        RECT 1298.680 1014.260 1298.940 1014.520 ;
        RECT 1298.680 990.460 1298.940 990.720 ;
        RECT 1298.220 990.120 1298.480 990.380 ;
        RECT 1298.680 869.420 1298.940 869.680 ;
        RECT 1299.140 869.420 1299.400 869.680 ;
        RECT 1298.680 862.280 1298.940 862.540 ;
        RECT 1298.220 814.340 1298.480 814.600 ;
        RECT 1298.680 717.440 1298.940 717.700 ;
        RECT 1298.680 668.820 1298.940 669.080 ;
        RECT 1298.680 621.560 1298.940 621.820 ;
        RECT 1298.680 620.880 1298.940 621.140 ;
        RECT 1298.680 613.740 1298.940 614.000 ;
        RECT 1299.140 613.740 1299.400 614.000 ;
        RECT 1298.220 476.040 1298.480 476.300 ;
        RECT 1299.140 476.040 1299.400 476.300 ;
        RECT 1298.220 448.500 1298.480 448.760 ;
        RECT 1298.680 447.820 1298.940 448.080 ;
        RECT 1298.680 420.620 1298.940 420.880 ;
        RECT 1298.220 355.340 1298.480 355.600 ;
        RECT 1298.220 304.000 1298.480 304.260 ;
        RECT 1298.220 303.320 1298.480 303.580 ;
        RECT 1297.760 144.540 1298.020 144.800 ;
        RECT 1298.680 144.540 1298.940 144.800 ;
        RECT 300.020 16.700 300.280 16.960 ;
        RECT 303.240 16.700 303.500 16.960 ;
      LAYER met2 ;
        RECT 1302.740 1700.410 1303.020 1704.000 ;
        RECT 1301.500 1700.270 1303.020 1700.410 ;
        RECT 1301.500 1666.670 1301.640 1700.270 ;
        RECT 1302.740 1700.000 1303.020 1700.270 ;
        RECT 1298.220 1666.350 1298.480 1666.670 ;
        RECT 1301.440 1666.350 1301.700 1666.670 ;
        RECT 1298.280 1608.190 1298.420 1666.350 ;
        RECT 1298.220 1607.870 1298.480 1608.190 ;
        RECT 1298.220 1593.930 1298.480 1594.250 ;
        RECT 1298.280 1593.650 1298.420 1593.930 ;
        RECT 1298.280 1593.510 1298.880 1593.650 ;
        RECT 1298.740 1463.090 1298.880 1593.510 ;
        RECT 1298.280 1462.950 1298.880 1463.090 ;
        RECT 1298.280 1449.070 1298.420 1462.950 ;
        RECT 1298.220 1448.750 1298.480 1449.070 ;
        RECT 1298.680 1386.870 1298.940 1387.190 ;
        RECT 1298.740 1338.765 1298.880 1386.870 ;
        RECT 1297.750 1338.395 1298.030 1338.765 ;
        RECT 1298.670 1338.395 1298.950 1338.765 ;
        RECT 1297.820 1290.485 1297.960 1338.395 ;
        RECT 1297.750 1290.115 1298.030 1290.485 ;
        RECT 1298.670 1290.115 1298.950 1290.485 ;
        RECT 1298.740 1270.230 1298.880 1290.115 ;
        RECT 1298.680 1269.910 1298.940 1270.230 ;
        RECT 1298.220 1242.370 1298.480 1242.690 ;
        RECT 1298.280 1242.010 1298.420 1242.370 ;
        RECT 1296.840 1241.690 1297.100 1242.010 ;
        RECT 1298.220 1241.690 1298.480 1242.010 ;
        RECT 1296.900 1193.925 1297.040 1241.690 ;
        RECT 1296.830 1193.555 1297.110 1193.925 ;
        RECT 1297.750 1193.555 1298.030 1193.925 ;
        RECT 1297.820 1182.930 1297.960 1193.555 ;
        RECT 1297.820 1182.790 1298.420 1182.930 ;
        RECT 1298.280 1159.050 1298.420 1182.790 ;
        RECT 1298.220 1158.730 1298.480 1159.050 ;
        RECT 1298.680 1110.790 1298.940 1111.110 ;
        RECT 1298.740 1087.310 1298.880 1110.790 ;
        RECT 1298.680 1086.990 1298.940 1087.310 ;
        RECT 1298.220 1086.650 1298.480 1086.970 ;
        RECT 1298.280 1062.490 1298.420 1086.650 ;
        RECT 1298.220 1062.170 1298.480 1062.490 ;
        RECT 1298.680 1014.230 1298.940 1014.550 ;
        RECT 1298.740 990.750 1298.880 1014.230 ;
        RECT 1298.680 990.430 1298.940 990.750 ;
        RECT 1298.220 990.090 1298.480 990.410 ;
        RECT 1298.280 966.125 1298.420 990.090 ;
        RECT 1298.210 965.755 1298.490 966.125 ;
        RECT 1299.130 965.755 1299.410 966.125 ;
        RECT 1299.200 869.710 1299.340 965.755 ;
        RECT 1298.680 869.390 1298.940 869.710 ;
        RECT 1299.140 869.390 1299.400 869.710 ;
        RECT 1298.740 862.570 1298.880 869.390 ;
        RECT 1298.680 862.250 1298.940 862.570 ;
        RECT 1298.220 814.310 1298.480 814.630 ;
        RECT 1298.280 748.410 1298.420 814.310 ;
        RECT 1298.280 748.270 1298.880 748.410 ;
        RECT 1298.740 717.730 1298.880 748.270 ;
        RECT 1298.680 717.410 1298.940 717.730 ;
        RECT 1298.680 668.790 1298.940 669.110 ;
        RECT 1298.740 621.850 1298.880 668.790 ;
        RECT 1298.680 621.530 1298.940 621.850 ;
        RECT 1298.680 620.850 1298.940 621.170 ;
        RECT 1298.740 614.030 1298.880 620.850 ;
        RECT 1298.680 613.710 1298.940 614.030 ;
        RECT 1299.140 613.710 1299.400 614.030 ;
        RECT 1299.200 476.330 1299.340 613.710 ;
        RECT 1298.220 476.010 1298.480 476.330 ;
        RECT 1299.140 476.010 1299.400 476.330 ;
        RECT 1298.280 448.790 1298.420 476.010 ;
        RECT 1298.220 448.470 1298.480 448.790 ;
        RECT 1298.680 447.790 1298.940 448.110 ;
        RECT 1298.740 420.910 1298.880 447.790 ;
        RECT 1298.680 420.590 1298.940 420.910 ;
        RECT 1298.220 355.310 1298.480 355.630 ;
        RECT 1298.280 304.290 1298.420 355.310 ;
        RECT 1298.220 303.970 1298.480 304.290 ;
        RECT 1298.220 303.290 1298.480 303.610 ;
        RECT 1298.280 265.610 1298.420 303.290 ;
        RECT 1298.280 265.470 1298.880 265.610 ;
        RECT 1298.740 144.830 1298.880 265.470 ;
        RECT 1297.760 144.510 1298.020 144.830 ;
        RECT 1298.680 144.510 1298.940 144.830 ;
        RECT 1297.820 96.970 1297.960 144.510 ;
        RECT 1297.820 96.830 1298.420 96.970 ;
        RECT 1298.280 62.970 1298.420 96.830 ;
        RECT 1298.280 62.830 1298.880 62.970 ;
        RECT 1298.740 51.525 1298.880 62.830 ;
        RECT 303.230 51.155 303.510 51.525 ;
        RECT 1298.670 51.155 1298.950 51.525 ;
        RECT 303.300 16.990 303.440 51.155 ;
        RECT 300.020 16.670 300.280 16.990 ;
        RECT 303.240 16.670 303.500 16.990 ;
        RECT 300.080 2.400 300.220 16.670 ;
        RECT 299.870 -4.800 300.430 2.400 ;
      LAYER via2 ;
        RECT 1297.750 1338.440 1298.030 1338.720 ;
        RECT 1298.670 1338.440 1298.950 1338.720 ;
        RECT 1297.750 1290.160 1298.030 1290.440 ;
        RECT 1298.670 1290.160 1298.950 1290.440 ;
        RECT 1296.830 1193.600 1297.110 1193.880 ;
        RECT 1297.750 1193.600 1298.030 1193.880 ;
        RECT 1298.210 965.800 1298.490 966.080 ;
        RECT 1299.130 965.800 1299.410 966.080 ;
        RECT 303.230 51.200 303.510 51.480 ;
        RECT 1298.670 51.200 1298.950 51.480 ;
      LAYER met3 ;
        RECT 1297.725 1338.730 1298.055 1338.745 ;
        RECT 1298.645 1338.730 1298.975 1338.745 ;
        RECT 1297.725 1338.430 1298.975 1338.730 ;
        RECT 1297.725 1338.415 1298.055 1338.430 ;
        RECT 1298.645 1338.415 1298.975 1338.430 ;
        RECT 1297.725 1290.450 1298.055 1290.465 ;
        RECT 1298.645 1290.450 1298.975 1290.465 ;
        RECT 1297.725 1290.150 1298.975 1290.450 ;
        RECT 1297.725 1290.135 1298.055 1290.150 ;
        RECT 1298.645 1290.135 1298.975 1290.150 ;
        RECT 1296.805 1193.890 1297.135 1193.905 ;
        RECT 1297.725 1193.890 1298.055 1193.905 ;
        RECT 1296.805 1193.590 1298.055 1193.890 ;
        RECT 1296.805 1193.575 1297.135 1193.590 ;
        RECT 1297.725 1193.575 1298.055 1193.590 ;
        RECT 1298.185 966.090 1298.515 966.105 ;
        RECT 1299.105 966.090 1299.435 966.105 ;
        RECT 1298.185 965.790 1299.435 966.090 ;
        RECT 1298.185 965.775 1298.515 965.790 ;
        RECT 1299.105 965.775 1299.435 965.790 ;
        RECT 303.205 51.490 303.535 51.505 ;
        RECT 1298.645 51.490 1298.975 51.505 ;
        RECT 303.205 51.190 1298.975 51.490 ;
        RECT 303.205 51.175 303.535 51.190 ;
        RECT 1298.645 51.175 1298.975 51.190 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 323.910 51.580 324.230 51.640 ;
        RECT 1311.530 51.580 1311.850 51.640 ;
        RECT 323.910 51.440 1311.850 51.580 ;
        RECT 323.910 51.380 324.230 51.440 ;
        RECT 1311.530 51.380 1311.850 51.440 ;
        RECT 317.930 16.900 318.250 16.960 ;
        RECT 323.910 16.900 324.230 16.960 ;
        RECT 317.930 16.760 324.230 16.900 ;
        RECT 317.930 16.700 318.250 16.760 ;
        RECT 323.910 16.700 324.230 16.760 ;
      LAYER via ;
        RECT 323.940 51.380 324.200 51.640 ;
        RECT 1311.560 51.380 1311.820 51.640 ;
        RECT 317.960 16.700 318.220 16.960 ;
        RECT 323.940 16.700 324.200 16.960 ;
      LAYER met2 ;
        RECT 1311.940 1700.410 1312.220 1704.000 ;
        RECT 1311.620 1700.270 1312.220 1700.410 ;
        RECT 1311.620 51.670 1311.760 1700.270 ;
        RECT 1311.940 1700.000 1312.220 1700.270 ;
        RECT 323.940 51.350 324.200 51.670 ;
        RECT 1311.560 51.350 1311.820 51.670 ;
        RECT 324.000 16.990 324.140 51.350 ;
        RECT 317.960 16.670 318.220 16.990 ;
        RECT 323.940 16.670 324.200 16.990 ;
        RECT 318.020 2.400 318.160 16.670 ;
        RECT 317.810 -4.800 318.370 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 335.870 26.420 336.190 26.480 ;
        RECT 1318.890 26.420 1319.210 26.480 ;
        RECT 335.870 26.280 1319.210 26.420 ;
        RECT 335.870 26.220 336.190 26.280 ;
        RECT 1318.890 26.220 1319.210 26.280 ;
      LAYER via ;
        RECT 335.900 26.220 336.160 26.480 ;
        RECT 1318.920 26.220 1319.180 26.480 ;
      LAYER met2 ;
        RECT 1321.140 1700.410 1321.420 1704.000 ;
        RECT 1318.980 1700.270 1321.420 1700.410 ;
        RECT 1318.980 26.510 1319.120 1700.270 ;
        RECT 1321.140 1700.000 1321.420 1700.270 ;
        RECT 335.900 26.190 336.160 26.510 ;
        RECT 1318.920 26.190 1319.180 26.510 ;
        RECT 335.960 2.400 336.100 26.190 ;
        RECT 335.750 -4.800 336.310 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1325.865 1442.025 1326.035 1490.475 ;
        RECT 1326.325 1256.045 1326.495 1304.155 ;
        RECT 1326.325 1014.305 1326.495 1028.415 ;
        RECT 1325.865 773.245 1326.035 821.015 ;
      LAYER mcon ;
        RECT 1325.865 1490.305 1326.035 1490.475 ;
        RECT 1326.325 1303.985 1326.495 1304.155 ;
        RECT 1326.325 1028.245 1326.495 1028.415 ;
        RECT 1325.865 820.845 1326.035 821.015 ;
      LAYER met1 ;
        RECT 1326.250 1642.440 1326.570 1642.500 ;
        RECT 1328.090 1642.440 1328.410 1642.500 ;
        RECT 1326.250 1642.300 1328.410 1642.440 ;
        RECT 1326.250 1642.240 1326.570 1642.300 ;
        RECT 1328.090 1642.240 1328.410 1642.300 ;
        RECT 1325.790 1497.600 1326.110 1497.660 ;
        RECT 1326.250 1497.600 1326.570 1497.660 ;
        RECT 1325.790 1497.460 1326.570 1497.600 ;
        RECT 1325.790 1497.400 1326.110 1497.460 ;
        RECT 1326.250 1497.400 1326.570 1497.460 ;
        RECT 1325.805 1490.460 1326.095 1490.505 ;
        RECT 1326.250 1490.460 1326.570 1490.520 ;
        RECT 1325.805 1490.320 1326.570 1490.460 ;
        RECT 1325.805 1490.275 1326.095 1490.320 ;
        RECT 1326.250 1490.260 1326.570 1490.320 ;
        RECT 1325.790 1442.180 1326.110 1442.240 ;
        RECT 1325.595 1442.040 1326.110 1442.180 ;
        RECT 1325.790 1441.980 1326.110 1442.040 ;
        RECT 1325.330 1401.040 1325.650 1401.100 ;
        RECT 1326.250 1401.040 1326.570 1401.100 ;
        RECT 1325.330 1400.900 1326.570 1401.040 ;
        RECT 1325.330 1400.840 1325.650 1400.900 ;
        RECT 1326.250 1400.840 1326.570 1400.900 ;
        RECT 1326.250 1304.140 1326.570 1304.200 ;
        RECT 1326.055 1304.000 1326.570 1304.140 ;
        RECT 1326.250 1303.940 1326.570 1304.000 ;
        RECT 1326.250 1256.200 1326.570 1256.260 ;
        RECT 1326.055 1256.060 1326.570 1256.200 ;
        RECT 1326.250 1256.000 1326.570 1256.060 ;
        RECT 1325.790 1221.660 1326.110 1221.920 ;
        RECT 1325.880 1220.900 1326.020 1221.660 ;
        RECT 1325.790 1220.640 1326.110 1220.900 ;
        RECT 1325.790 1159.980 1326.110 1160.040 ;
        RECT 1325.790 1159.840 1326.480 1159.980 ;
        RECT 1325.790 1159.780 1326.110 1159.840 ;
        RECT 1326.340 1159.360 1326.480 1159.840 ;
        RECT 1326.250 1159.100 1326.570 1159.360 ;
        RECT 1325.790 1063.420 1326.110 1063.480 ;
        RECT 1325.790 1063.280 1326.480 1063.420 ;
        RECT 1325.790 1063.220 1326.110 1063.280 ;
        RECT 1326.340 1062.800 1326.480 1063.280 ;
        RECT 1326.250 1062.540 1326.570 1062.800 ;
        RECT 1326.250 1028.400 1326.570 1028.460 ;
        RECT 1326.055 1028.260 1326.570 1028.400 ;
        RECT 1326.250 1028.200 1326.570 1028.260 ;
        RECT 1326.250 1014.460 1326.570 1014.520 ;
        RECT 1326.055 1014.320 1326.570 1014.460 ;
        RECT 1326.250 1014.260 1326.570 1014.320 ;
        RECT 1326.250 966.520 1326.570 966.580 ;
        RECT 1325.880 966.380 1326.570 966.520 ;
        RECT 1325.880 966.240 1326.020 966.380 ;
        RECT 1326.250 966.320 1326.570 966.380 ;
        RECT 1325.790 965.980 1326.110 966.240 ;
        RECT 1325.790 910.760 1326.110 910.820 ;
        RECT 1326.250 910.760 1326.570 910.820 ;
        RECT 1325.790 910.620 1326.570 910.760 ;
        RECT 1325.790 910.560 1326.110 910.620 ;
        RECT 1326.250 910.560 1326.570 910.620 ;
        RECT 1325.805 821.000 1326.095 821.045 ;
        RECT 1326.250 821.000 1326.570 821.060 ;
        RECT 1325.805 820.860 1326.570 821.000 ;
        RECT 1325.805 820.815 1326.095 820.860 ;
        RECT 1326.250 820.800 1326.570 820.860 ;
        RECT 1325.790 773.400 1326.110 773.460 ;
        RECT 1325.595 773.260 1326.110 773.400 ;
        RECT 1325.790 773.200 1326.110 773.260 ;
        RECT 1325.790 738.520 1326.110 738.780 ;
        RECT 1325.880 738.100 1326.020 738.520 ;
        RECT 1325.790 737.840 1326.110 738.100 ;
        RECT 1325.330 603.740 1325.650 603.800 ;
        RECT 1326.250 603.740 1326.570 603.800 ;
        RECT 1325.330 603.600 1326.570 603.740 ;
        RECT 1325.330 603.540 1325.650 603.600 ;
        RECT 1326.250 603.540 1326.570 603.600 ;
        RECT 1325.790 331.400 1326.110 331.460 ;
        RECT 1326.250 331.400 1326.570 331.460 ;
        RECT 1325.790 331.260 1326.570 331.400 ;
        RECT 1325.790 331.200 1326.110 331.260 ;
        RECT 1326.250 331.200 1326.570 331.260 ;
        RECT 1325.790 144.740 1326.110 144.800 ;
        RECT 1326.250 144.740 1326.570 144.800 ;
        RECT 1325.790 144.600 1326.570 144.740 ;
        RECT 1325.790 144.540 1326.110 144.600 ;
        RECT 1326.250 144.540 1326.570 144.600 ;
        RECT 358.410 72.660 358.730 72.720 ;
        RECT 1325.790 72.660 1326.110 72.720 ;
        RECT 358.410 72.520 1326.110 72.660 ;
        RECT 358.410 72.460 358.730 72.520 ;
        RECT 1325.790 72.460 1326.110 72.520 ;
        RECT 353.350 16.900 353.670 16.960 ;
        RECT 358.410 16.900 358.730 16.960 ;
        RECT 353.350 16.760 358.730 16.900 ;
        RECT 353.350 16.700 353.670 16.760 ;
        RECT 358.410 16.700 358.730 16.760 ;
      LAYER via ;
        RECT 1326.280 1642.240 1326.540 1642.500 ;
        RECT 1328.120 1642.240 1328.380 1642.500 ;
        RECT 1325.820 1497.400 1326.080 1497.660 ;
        RECT 1326.280 1497.400 1326.540 1497.660 ;
        RECT 1326.280 1490.260 1326.540 1490.520 ;
        RECT 1325.820 1441.980 1326.080 1442.240 ;
        RECT 1325.360 1400.840 1325.620 1401.100 ;
        RECT 1326.280 1400.840 1326.540 1401.100 ;
        RECT 1326.280 1303.940 1326.540 1304.200 ;
        RECT 1326.280 1256.000 1326.540 1256.260 ;
        RECT 1325.820 1221.660 1326.080 1221.920 ;
        RECT 1325.820 1220.640 1326.080 1220.900 ;
        RECT 1325.820 1159.780 1326.080 1160.040 ;
        RECT 1326.280 1159.100 1326.540 1159.360 ;
        RECT 1325.820 1063.220 1326.080 1063.480 ;
        RECT 1326.280 1062.540 1326.540 1062.800 ;
        RECT 1326.280 1028.200 1326.540 1028.460 ;
        RECT 1326.280 1014.260 1326.540 1014.520 ;
        RECT 1326.280 966.320 1326.540 966.580 ;
        RECT 1325.820 965.980 1326.080 966.240 ;
        RECT 1325.820 910.560 1326.080 910.820 ;
        RECT 1326.280 910.560 1326.540 910.820 ;
        RECT 1326.280 820.800 1326.540 821.060 ;
        RECT 1325.820 773.200 1326.080 773.460 ;
        RECT 1325.820 738.520 1326.080 738.780 ;
        RECT 1325.820 737.840 1326.080 738.100 ;
        RECT 1325.360 603.540 1325.620 603.800 ;
        RECT 1326.280 603.540 1326.540 603.800 ;
        RECT 1325.820 331.200 1326.080 331.460 ;
        RECT 1326.280 331.200 1326.540 331.460 ;
        RECT 1325.820 144.540 1326.080 144.800 ;
        RECT 1326.280 144.540 1326.540 144.800 ;
        RECT 358.440 72.460 358.700 72.720 ;
        RECT 1325.820 72.460 1326.080 72.720 ;
        RECT 353.380 16.700 353.640 16.960 ;
        RECT 358.440 16.700 358.700 16.960 ;
      LAYER met2 ;
        RECT 1330.340 1700.410 1330.620 1704.000 ;
        RECT 1328.180 1700.270 1330.620 1700.410 ;
        RECT 1328.180 1642.530 1328.320 1700.270 ;
        RECT 1330.340 1700.000 1330.620 1700.270 ;
        RECT 1326.280 1642.210 1326.540 1642.530 ;
        RECT 1328.120 1642.210 1328.380 1642.530 ;
        RECT 1326.340 1559.650 1326.480 1642.210 ;
        RECT 1325.880 1559.510 1326.480 1559.650 ;
        RECT 1325.880 1497.690 1326.020 1559.510 ;
        RECT 1325.820 1497.370 1326.080 1497.690 ;
        RECT 1326.280 1497.370 1326.540 1497.690 ;
        RECT 1326.340 1490.550 1326.480 1497.370 ;
        RECT 1326.280 1490.230 1326.540 1490.550 ;
        RECT 1325.820 1441.950 1326.080 1442.270 ;
        RECT 1325.880 1402.570 1326.020 1441.950 ;
        RECT 1325.880 1402.430 1326.480 1402.570 ;
        RECT 1326.340 1401.130 1326.480 1402.430 ;
        RECT 1325.360 1400.810 1325.620 1401.130 ;
        RECT 1326.280 1400.810 1326.540 1401.130 ;
        RECT 1325.420 1393.845 1325.560 1400.810 ;
        RECT 1325.350 1393.475 1325.630 1393.845 ;
        RECT 1326.730 1393.475 1327.010 1393.845 ;
        RECT 1326.800 1317.570 1326.940 1393.475 ;
        RECT 1326.340 1317.430 1326.940 1317.570 ;
        RECT 1326.340 1304.230 1326.480 1317.430 ;
        RECT 1326.280 1303.910 1326.540 1304.230 ;
        RECT 1326.280 1256.200 1326.540 1256.290 ;
        RECT 1325.880 1256.060 1326.540 1256.200 ;
        RECT 1325.880 1221.950 1326.020 1256.060 ;
        RECT 1326.280 1255.970 1326.540 1256.060 ;
        RECT 1325.820 1221.630 1326.080 1221.950 ;
        RECT 1325.820 1220.610 1326.080 1220.930 ;
        RECT 1325.880 1160.070 1326.020 1220.610 ;
        RECT 1325.820 1159.750 1326.080 1160.070 ;
        RECT 1326.280 1159.070 1326.540 1159.390 ;
        RECT 1326.340 1134.650 1326.480 1159.070 ;
        RECT 1325.880 1134.510 1326.480 1134.650 ;
        RECT 1325.880 1063.510 1326.020 1134.510 ;
        RECT 1325.820 1063.190 1326.080 1063.510 ;
        RECT 1326.280 1062.510 1326.540 1062.830 ;
        RECT 1326.340 1028.490 1326.480 1062.510 ;
        RECT 1326.280 1028.170 1326.540 1028.490 ;
        RECT 1326.280 1014.230 1326.540 1014.550 ;
        RECT 1326.340 966.610 1326.480 1014.230 ;
        RECT 1326.280 966.290 1326.540 966.610 ;
        RECT 1325.820 966.010 1326.080 966.270 ;
        RECT 1325.420 965.950 1326.080 966.010 ;
        RECT 1325.420 965.870 1326.020 965.950 ;
        RECT 1325.420 931.330 1325.560 965.870 ;
        RECT 1325.420 931.190 1326.020 931.330 ;
        RECT 1325.880 910.850 1326.020 931.190 ;
        RECT 1325.820 910.530 1326.080 910.850 ;
        RECT 1326.280 910.530 1326.540 910.850 ;
        RECT 1326.340 886.565 1326.480 910.530 ;
        RECT 1326.270 886.195 1326.550 886.565 ;
        RECT 1326.270 820.915 1326.550 821.285 ;
        RECT 1326.280 820.770 1326.540 820.915 ;
        RECT 1325.820 773.170 1326.080 773.490 ;
        RECT 1325.880 738.810 1326.020 773.170 ;
        RECT 1325.820 738.490 1326.080 738.810 ;
        RECT 1325.820 737.810 1326.080 738.130 ;
        RECT 1325.880 677.125 1326.020 737.810 ;
        RECT 1325.810 676.755 1326.090 677.125 ;
        RECT 1325.810 676.075 1326.090 676.445 ;
        RECT 1325.880 628.050 1326.020 676.075 ;
        RECT 1325.880 627.910 1326.480 628.050 ;
        RECT 1326.340 603.830 1326.480 627.910 ;
        RECT 1325.360 603.510 1325.620 603.830 ;
        RECT 1326.280 603.510 1326.540 603.830 ;
        RECT 1325.420 579.885 1325.560 603.510 ;
        RECT 1325.350 579.515 1325.630 579.885 ;
        RECT 1326.270 579.515 1326.550 579.885 ;
        RECT 1326.340 500.210 1326.480 579.515 ;
        RECT 1325.880 500.070 1326.480 500.210 ;
        RECT 1325.880 387.330 1326.020 500.070 ;
        RECT 1325.880 387.190 1326.480 387.330 ;
        RECT 1326.340 386.480 1326.480 387.190 ;
        RECT 1325.880 386.340 1326.480 386.480 ;
        RECT 1325.880 331.490 1326.020 386.340 ;
        RECT 1325.820 331.170 1326.080 331.490 ;
        RECT 1326.280 331.170 1326.540 331.490 ;
        RECT 1326.340 144.830 1326.480 331.170 ;
        RECT 1325.820 144.510 1326.080 144.830 ;
        RECT 1326.280 144.510 1326.540 144.830 ;
        RECT 1325.880 72.750 1326.020 144.510 ;
        RECT 358.440 72.430 358.700 72.750 ;
        RECT 1325.820 72.430 1326.080 72.750 ;
        RECT 358.500 16.990 358.640 72.430 ;
        RECT 353.380 16.670 353.640 16.990 ;
        RECT 358.440 16.670 358.700 16.990 ;
        RECT 353.440 2.400 353.580 16.670 ;
        RECT 353.230 -4.800 353.790 2.400 ;
      LAYER via2 ;
        RECT 1325.350 1393.520 1325.630 1393.800 ;
        RECT 1326.730 1393.520 1327.010 1393.800 ;
        RECT 1326.270 886.240 1326.550 886.520 ;
        RECT 1326.270 820.960 1326.550 821.240 ;
        RECT 1325.810 676.800 1326.090 677.080 ;
        RECT 1325.810 676.120 1326.090 676.400 ;
        RECT 1325.350 579.560 1325.630 579.840 ;
        RECT 1326.270 579.560 1326.550 579.840 ;
      LAYER met3 ;
        RECT 1325.325 1393.810 1325.655 1393.825 ;
        RECT 1326.705 1393.810 1327.035 1393.825 ;
        RECT 1325.325 1393.510 1327.035 1393.810 ;
        RECT 1325.325 1393.495 1325.655 1393.510 ;
        RECT 1326.705 1393.495 1327.035 1393.510 ;
        RECT 1326.245 886.540 1326.575 886.545 ;
        RECT 1325.990 886.530 1326.575 886.540 ;
        RECT 1325.990 886.230 1326.800 886.530 ;
        RECT 1325.990 886.220 1326.575 886.230 ;
        RECT 1326.245 886.215 1326.575 886.220 ;
        RECT 1326.245 821.260 1326.575 821.265 ;
        RECT 1325.990 821.250 1326.575 821.260 ;
        RECT 1325.790 820.950 1326.575 821.250 ;
        RECT 1325.990 820.940 1326.575 820.950 ;
        RECT 1326.245 820.935 1326.575 820.940 ;
        RECT 1325.785 677.090 1326.115 677.105 ;
        RECT 1325.785 676.775 1326.330 677.090 ;
        RECT 1326.030 676.425 1326.330 676.775 ;
        RECT 1325.785 676.110 1326.330 676.425 ;
        RECT 1325.785 676.095 1326.115 676.110 ;
        RECT 1325.325 579.850 1325.655 579.865 ;
        RECT 1326.245 579.850 1326.575 579.865 ;
        RECT 1325.325 579.550 1326.575 579.850 ;
        RECT 1325.325 579.535 1325.655 579.550 ;
        RECT 1326.245 579.535 1326.575 579.550 ;
      LAYER via3 ;
        RECT 1326.020 886.220 1326.340 886.540 ;
        RECT 1326.020 820.940 1326.340 821.260 ;
      LAYER met4 ;
        RECT 1326.015 886.215 1326.345 886.545 ;
        RECT 1326.030 821.265 1326.330 886.215 ;
        RECT 1326.015 820.935 1326.345 821.265 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 372.210 73.000 372.530 73.060 ;
        RECT 1339.130 73.000 1339.450 73.060 ;
        RECT 372.210 72.860 1339.450 73.000 ;
        RECT 372.210 72.800 372.530 72.860 ;
        RECT 1339.130 72.800 1339.450 72.860 ;
      LAYER via ;
        RECT 372.240 72.800 372.500 73.060 ;
        RECT 1339.160 72.800 1339.420 73.060 ;
      LAYER met2 ;
        RECT 1339.540 1700.410 1339.820 1704.000 ;
        RECT 1339.220 1700.270 1339.820 1700.410 ;
        RECT 1339.220 73.090 1339.360 1700.270 ;
        RECT 1339.540 1700.000 1339.820 1700.270 ;
        RECT 372.240 72.770 372.500 73.090 ;
        RECT 1339.160 72.770 1339.420 73.090 ;
        RECT 372.300 16.900 372.440 72.770 ;
        RECT 371.380 16.760 372.440 16.900 ;
        RECT 371.380 2.400 371.520 16.760 ;
        RECT 371.170 -4.800 371.730 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 392.910 73.340 393.230 73.400 ;
        RECT 1346.030 73.340 1346.350 73.400 ;
        RECT 392.910 73.200 1346.350 73.340 ;
        RECT 392.910 73.140 393.230 73.200 ;
        RECT 1346.030 73.140 1346.350 73.200 ;
        RECT 389.230 16.220 389.550 16.280 ;
        RECT 392.910 16.220 393.230 16.280 ;
        RECT 389.230 16.080 393.230 16.220 ;
        RECT 389.230 16.020 389.550 16.080 ;
        RECT 392.910 16.020 393.230 16.080 ;
      LAYER via ;
        RECT 392.940 73.140 393.200 73.400 ;
        RECT 1346.060 73.140 1346.320 73.400 ;
        RECT 389.260 16.020 389.520 16.280 ;
        RECT 392.940 16.020 393.200 16.280 ;
      LAYER met2 ;
        RECT 1348.740 1700.410 1349.020 1704.000 ;
        RECT 1346.120 1700.270 1349.020 1700.410 ;
        RECT 1346.120 73.430 1346.260 1700.270 ;
        RECT 1348.740 1700.000 1349.020 1700.270 ;
        RECT 392.940 73.110 393.200 73.430 ;
        RECT 1346.060 73.110 1346.320 73.430 ;
        RECT 393.000 16.310 393.140 73.110 ;
        RECT 389.260 15.990 389.520 16.310 ;
        RECT 392.940 15.990 393.200 16.310 ;
        RECT 389.320 2.400 389.460 15.990 ;
        RECT 389.110 -4.800 389.670 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1353.465 1497.445 1353.635 1545.555 ;
        RECT 1353.005 1304.325 1353.175 1393.575 ;
        RECT 1353.465 1062.245 1353.635 1077.035 ;
        RECT 1353.465 1027.905 1353.635 1055.615 ;
        RECT 1353.005 965.685 1353.175 980.475 ;
        RECT 1353.005 917.405 1353.175 959.055 ;
        RECT 1353.465 331.245 1353.635 379.355 ;
        RECT 1353.465 89.845 1353.635 137.955 ;
      LAYER mcon ;
        RECT 1353.465 1545.385 1353.635 1545.555 ;
        RECT 1353.005 1393.405 1353.175 1393.575 ;
        RECT 1353.465 1076.865 1353.635 1077.035 ;
        RECT 1353.465 1055.445 1353.635 1055.615 ;
        RECT 1353.005 980.305 1353.175 980.475 ;
        RECT 1353.005 958.885 1353.175 959.055 ;
        RECT 1353.465 379.185 1353.635 379.355 ;
        RECT 1353.465 137.785 1353.635 137.955 ;
      LAYER met1 ;
        RECT 1353.850 1642.440 1354.170 1642.500 ;
        RECT 1355.690 1642.440 1356.010 1642.500 ;
        RECT 1353.850 1642.300 1356.010 1642.440 ;
        RECT 1353.850 1642.240 1354.170 1642.300 ;
        RECT 1355.690 1642.240 1356.010 1642.300 ;
        RECT 1353.390 1545.540 1353.710 1545.600 ;
        RECT 1353.195 1545.400 1353.710 1545.540 ;
        RECT 1353.390 1545.340 1353.710 1545.400 ;
        RECT 1353.405 1497.600 1353.695 1497.645 ;
        RECT 1353.850 1497.600 1354.170 1497.660 ;
        RECT 1353.405 1497.460 1354.170 1497.600 ;
        RECT 1353.405 1497.415 1353.695 1497.460 ;
        RECT 1353.850 1497.400 1354.170 1497.460 ;
        RECT 1353.850 1490.460 1354.170 1490.520 ;
        RECT 1354.310 1490.460 1354.630 1490.520 ;
        RECT 1353.850 1490.320 1354.630 1490.460 ;
        RECT 1353.850 1490.260 1354.170 1490.320 ;
        RECT 1354.310 1490.260 1354.630 1490.320 ;
        RECT 1352.930 1400.700 1353.250 1400.760 ;
        RECT 1354.310 1400.700 1354.630 1400.760 ;
        RECT 1352.930 1400.560 1354.630 1400.700 ;
        RECT 1352.930 1400.500 1353.250 1400.560 ;
        RECT 1354.310 1400.500 1354.630 1400.560 ;
        RECT 1352.930 1393.560 1353.250 1393.620 ;
        RECT 1352.735 1393.420 1353.250 1393.560 ;
        RECT 1352.930 1393.360 1353.250 1393.420 ;
        RECT 1352.945 1304.480 1353.235 1304.525 ;
        RECT 1353.850 1304.480 1354.170 1304.540 ;
        RECT 1352.945 1304.340 1354.170 1304.480 ;
        RECT 1352.945 1304.295 1353.235 1304.340 ;
        RECT 1353.850 1304.280 1354.170 1304.340 ;
        RECT 1353.390 1256.200 1353.710 1256.260 ;
        RECT 1354.770 1256.200 1355.090 1256.260 ;
        RECT 1353.390 1256.060 1355.090 1256.200 ;
        RECT 1353.390 1256.000 1353.710 1256.060 ;
        RECT 1354.770 1256.000 1355.090 1256.060 ;
        RECT 1353.390 1221.320 1353.710 1221.580 ;
        RECT 1353.480 1220.840 1353.620 1221.320 ;
        RECT 1353.850 1220.840 1354.170 1220.900 ;
        RECT 1353.480 1220.700 1354.170 1220.840 ;
        RECT 1353.850 1220.640 1354.170 1220.700 ;
        RECT 1352.930 1152.500 1353.250 1152.560 ;
        RECT 1353.390 1152.500 1353.710 1152.560 ;
        RECT 1352.930 1152.360 1353.710 1152.500 ;
        RECT 1352.930 1152.300 1353.250 1152.360 ;
        RECT 1353.390 1152.300 1353.710 1152.360 ;
        RECT 1353.850 1124.960 1354.170 1125.020 ;
        RECT 1353.480 1124.820 1354.170 1124.960 ;
        RECT 1353.480 1124.680 1353.620 1124.820 ;
        RECT 1353.850 1124.760 1354.170 1124.820 ;
        RECT 1353.390 1124.420 1353.710 1124.680 ;
        RECT 1353.390 1077.020 1353.710 1077.080 ;
        RECT 1353.195 1076.880 1353.710 1077.020 ;
        RECT 1353.390 1076.820 1353.710 1076.880 ;
        RECT 1353.390 1062.400 1353.710 1062.460 ;
        RECT 1353.195 1062.260 1353.710 1062.400 ;
        RECT 1353.390 1062.200 1353.710 1062.260 ;
        RECT 1353.390 1055.600 1353.710 1055.660 ;
        RECT 1353.195 1055.460 1353.710 1055.600 ;
        RECT 1353.390 1055.400 1353.710 1055.460 ;
        RECT 1353.390 1028.060 1353.710 1028.120 ;
        RECT 1353.195 1027.920 1353.710 1028.060 ;
        RECT 1353.390 1027.860 1353.710 1027.920 ;
        RECT 1352.945 980.460 1353.235 980.505 ;
        RECT 1353.850 980.460 1354.170 980.520 ;
        RECT 1352.945 980.320 1354.170 980.460 ;
        RECT 1352.945 980.275 1353.235 980.320 ;
        RECT 1353.850 980.260 1354.170 980.320 ;
        RECT 1352.930 965.840 1353.250 965.900 ;
        RECT 1352.735 965.700 1353.250 965.840 ;
        RECT 1352.930 965.640 1353.250 965.700 ;
        RECT 1352.930 959.040 1353.250 959.100 ;
        RECT 1352.735 958.900 1353.250 959.040 ;
        RECT 1352.930 958.840 1353.250 958.900 ;
        RECT 1352.945 917.560 1353.235 917.605 ;
        RECT 1353.390 917.560 1353.710 917.620 ;
        RECT 1352.945 917.420 1353.710 917.560 ;
        RECT 1352.945 917.375 1353.235 917.420 ;
        RECT 1353.390 917.360 1353.710 917.420 ;
        RECT 1353.390 869.620 1353.710 869.680 ;
        RECT 1354.310 869.620 1354.630 869.680 ;
        RECT 1353.390 869.480 1354.630 869.620 ;
        RECT 1353.390 869.420 1353.710 869.480 ;
        RECT 1354.310 869.420 1354.630 869.480 ;
        RECT 1353.390 835.080 1353.710 835.340 ;
        RECT 1353.480 834.600 1353.620 835.080 ;
        RECT 1353.850 834.600 1354.170 834.660 ;
        RECT 1353.480 834.460 1354.170 834.600 ;
        RECT 1353.850 834.400 1354.170 834.460 ;
        RECT 1352.930 627.880 1353.250 627.940 ;
        RECT 1353.850 627.880 1354.170 627.940 ;
        RECT 1352.930 627.740 1354.170 627.880 ;
        RECT 1352.930 627.680 1353.250 627.740 ;
        RECT 1353.850 627.680 1354.170 627.740 ;
        RECT 1352.930 434.420 1353.250 434.480 ;
        RECT 1354.310 434.420 1354.630 434.480 ;
        RECT 1352.930 434.280 1354.630 434.420 ;
        RECT 1352.930 434.220 1353.250 434.280 ;
        RECT 1354.310 434.220 1354.630 434.280 ;
        RECT 1353.390 386.480 1353.710 386.540 ;
        RECT 1354.310 386.480 1354.630 386.540 ;
        RECT 1353.390 386.340 1354.630 386.480 ;
        RECT 1353.390 386.280 1353.710 386.340 ;
        RECT 1354.310 386.280 1354.630 386.340 ;
        RECT 1353.390 379.340 1353.710 379.400 ;
        RECT 1353.195 379.200 1353.710 379.340 ;
        RECT 1353.390 379.140 1353.710 379.200 ;
        RECT 1353.405 331.400 1353.695 331.445 ;
        RECT 1353.850 331.400 1354.170 331.460 ;
        RECT 1353.405 331.260 1354.170 331.400 ;
        RECT 1353.405 331.215 1353.695 331.260 ;
        RECT 1353.850 331.200 1354.170 331.260 ;
        RECT 1353.850 304.200 1354.170 304.260 ;
        RECT 1353.480 304.060 1354.170 304.200 ;
        RECT 1353.480 303.580 1353.620 304.060 ;
        RECT 1353.850 304.000 1354.170 304.060 ;
        RECT 1353.390 303.320 1353.710 303.580 ;
        RECT 1353.390 235.180 1353.710 235.240 ;
        RECT 1353.020 235.040 1353.710 235.180 ;
        RECT 1353.020 234.900 1353.160 235.040 ;
        RECT 1353.390 234.980 1353.710 235.040 ;
        RECT 1352.930 234.640 1353.250 234.900 ;
        RECT 1353.390 145.080 1353.710 145.140 ;
        RECT 1353.850 145.080 1354.170 145.140 ;
        RECT 1353.390 144.940 1354.170 145.080 ;
        RECT 1353.390 144.880 1353.710 144.940 ;
        RECT 1353.850 144.880 1354.170 144.940 ;
        RECT 1353.405 137.940 1353.695 137.985 ;
        RECT 1353.850 137.940 1354.170 138.000 ;
        RECT 1353.405 137.800 1354.170 137.940 ;
        RECT 1353.405 137.755 1353.695 137.800 ;
        RECT 1353.850 137.740 1354.170 137.800 ;
        RECT 1353.390 90.000 1353.710 90.060 ;
        RECT 1353.195 89.860 1353.710 90.000 ;
        RECT 1353.390 89.800 1353.710 89.860 ;
        RECT 413.610 73.680 413.930 73.740 ;
        RECT 1353.390 73.680 1353.710 73.740 ;
        RECT 413.610 73.540 1353.710 73.680 ;
        RECT 413.610 73.480 413.930 73.540 ;
        RECT 1353.390 73.480 1353.710 73.540 ;
        RECT 407.170 16.220 407.490 16.280 ;
        RECT 413.610 16.220 413.930 16.280 ;
        RECT 407.170 16.080 413.930 16.220 ;
        RECT 407.170 16.020 407.490 16.080 ;
        RECT 413.610 16.020 413.930 16.080 ;
      LAYER via ;
        RECT 1353.880 1642.240 1354.140 1642.500 ;
        RECT 1355.720 1642.240 1355.980 1642.500 ;
        RECT 1353.420 1545.340 1353.680 1545.600 ;
        RECT 1353.880 1497.400 1354.140 1497.660 ;
        RECT 1353.880 1490.260 1354.140 1490.520 ;
        RECT 1354.340 1490.260 1354.600 1490.520 ;
        RECT 1352.960 1400.500 1353.220 1400.760 ;
        RECT 1354.340 1400.500 1354.600 1400.760 ;
        RECT 1352.960 1393.360 1353.220 1393.620 ;
        RECT 1353.880 1304.280 1354.140 1304.540 ;
        RECT 1353.420 1256.000 1353.680 1256.260 ;
        RECT 1354.800 1256.000 1355.060 1256.260 ;
        RECT 1353.420 1221.320 1353.680 1221.580 ;
        RECT 1353.880 1220.640 1354.140 1220.900 ;
        RECT 1352.960 1152.300 1353.220 1152.560 ;
        RECT 1353.420 1152.300 1353.680 1152.560 ;
        RECT 1353.880 1124.760 1354.140 1125.020 ;
        RECT 1353.420 1124.420 1353.680 1124.680 ;
        RECT 1353.420 1076.820 1353.680 1077.080 ;
        RECT 1353.420 1062.200 1353.680 1062.460 ;
        RECT 1353.420 1055.400 1353.680 1055.660 ;
        RECT 1353.420 1027.860 1353.680 1028.120 ;
        RECT 1353.880 980.260 1354.140 980.520 ;
        RECT 1352.960 965.640 1353.220 965.900 ;
        RECT 1352.960 958.840 1353.220 959.100 ;
        RECT 1353.420 917.360 1353.680 917.620 ;
        RECT 1353.420 869.420 1353.680 869.680 ;
        RECT 1354.340 869.420 1354.600 869.680 ;
        RECT 1353.420 835.080 1353.680 835.340 ;
        RECT 1353.880 834.400 1354.140 834.660 ;
        RECT 1352.960 627.680 1353.220 627.940 ;
        RECT 1353.880 627.680 1354.140 627.940 ;
        RECT 1352.960 434.220 1353.220 434.480 ;
        RECT 1354.340 434.220 1354.600 434.480 ;
        RECT 1353.420 386.280 1353.680 386.540 ;
        RECT 1354.340 386.280 1354.600 386.540 ;
        RECT 1353.420 379.140 1353.680 379.400 ;
        RECT 1353.880 331.200 1354.140 331.460 ;
        RECT 1353.880 304.000 1354.140 304.260 ;
        RECT 1353.420 303.320 1353.680 303.580 ;
        RECT 1353.420 234.980 1353.680 235.240 ;
        RECT 1352.960 234.640 1353.220 234.900 ;
        RECT 1353.420 144.880 1353.680 145.140 ;
        RECT 1353.880 144.880 1354.140 145.140 ;
        RECT 1353.880 137.740 1354.140 138.000 ;
        RECT 1353.420 89.800 1353.680 90.060 ;
        RECT 413.640 73.480 413.900 73.740 ;
        RECT 1353.420 73.480 1353.680 73.740 ;
        RECT 407.200 16.020 407.460 16.280 ;
        RECT 413.640 16.020 413.900 16.280 ;
      LAYER met2 ;
        RECT 1357.940 1700.410 1358.220 1704.000 ;
        RECT 1355.780 1700.270 1358.220 1700.410 ;
        RECT 1355.780 1642.530 1355.920 1700.270 ;
        RECT 1357.940 1700.000 1358.220 1700.270 ;
        RECT 1353.880 1642.210 1354.140 1642.530 ;
        RECT 1355.720 1642.210 1355.980 1642.530 ;
        RECT 1353.940 1559.650 1354.080 1642.210 ;
        RECT 1353.480 1559.510 1354.080 1559.650 ;
        RECT 1353.480 1545.630 1353.620 1559.510 ;
        RECT 1353.420 1545.310 1353.680 1545.630 ;
        RECT 1353.880 1497.370 1354.140 1497.690 ;
        RECT 1353.940 1490.550 1354.080 1497.370 ;
        RECT 1353.880 1490.230 1354.140 1490.550 ;
        RECT 1354.340 1490.230 1354.600 1490.550 ;
        RECT 1354.400 1400.790 1354.540 1490.230 ;
        RECT 1352.960 1400.470 1353.220 1400.790 ;
        RECT 1354.340 1400.470 1354.600 1400.790 ;
        RECT 1353.020 1393.650 1353.160 1400.470 ;
        RECT 1352.960 1393.330 1353.220 1393.650 ;
        RECT 1353.880 1304.250 1354.140 1304.570 ;
        RECT 1353.940 1304.085 1354.080 1304.250 ;
        RECT 1353.870 1303.715 1354.150 1304.085 ;
        RECT 1354.790 1303.715 1355.070 1304.085 ;
        RECT 1354.860 1256.290 1355.000 1303.715 ;
        RECT 1353.420 1255.970 1353.680 1256.290 ;
        RECT 1354.800 1255.970 1355.060 1256.290 ;
        RECT 1353.480 1221.610 1353.620 1255.970 ;
        RECT 1353.420 1221.290 1353.680 1221.610 ;
        RECT 1353.880 1220.610 1354.140 1220.930 ;
        RECT 1353.940 1207.410 1354.080 1220.610 ;
        RECT 1353.480 1207.270 1354.080 1207.410 ;
        RECT 1353.480 1174.090 1353.620 1207.270 ;
        RECT 1353.020 1173.950 1353.620 1174.090 ;
        RECT 1353.020 1152.590 1353.160 1173.950 ;
        RECT 1352.960 1152.270 1353.220 1152.590 ;
        RECT 1353.420 1152.330 1353.680 1152.590 ;
        RECT 1353.420 1152.270 1354.080 1152.330 ;
        RECT 1353.480 1152.190 1354.080 1152.270 ;
        RECT 1353.940 1125.050 1354.080 1152.190 ;
        RECT 1353.880 1124.730 1354.140 1125.050 ;
        RECT 1353.420 1124.390 1353.680 1124.710 ;
        RECT 1353.480 1077.110 1353.620 1124.390 ;
        RECT 1353.420 1076.790 1353.680 1077.110 ;
        RECT 1353.420 1062.170 1353.680 1062.490 ;
        RECT 1353.480 1055.690 1353.620 1062.170 ;
        RECT 1353.420 1055.370 1353.680 1055.690 ;
        RECT 1353.420 1027.830 1353.680 1028.150 ;
        RECT 1353.480 1007.490 1353.620 1027.830 ;
        RECT 1353.480 1007.350 1354.080 1007.490 ;
        RECT 1353.940 980.550 1354.080 1007.350 ;
        RECT 1353.880 980.230 1354.140 980.550 ;
        RECT 1352.960 965.610 1353.220 965.930 ;
        RECT 1353.020 959.130 1353.160 965.610 ;
        RECT 1352.960 958.810 1353.220 959.130 ;
        RECT 1353.420 917.330 1353.680 917.650 ;
        RECT 1353.480 910.930 1353.620 917.330 ;
        RECT 1353.480 910.790 1354.080 910.930 ;
        RECT 1353.940 893.930 1354.080 910.790 ;
        RECT 1353.940 893.790 1354.540 893.930 ;
        RECT 1354.400 869.710 1354.540 893.790 ;
        RECT 1353.420 869.390 1353.680 869.710 ;
        RECT 1354.340 869.390 1354.600 869.710 ;
        RECT 1353.480 835.370 1353.620 869.390 ;
        RECT 1353.420 835.050 1353.680 835.370 ;
        RECT 1353.880 834.370 1354.140 834.690 ;
        RECT 1353.940 691.290 1354.080 834.370 ;
        RECT 1353.940 691.150 1354.540 691.290 ;
        RECT 1354.400 676.445 1354.540 691.150 ;
        RECT 1353.410 676.075 1353.690 676.445 ;
        RECT 1354.330 676.075 1354.610 676.445 ;
        RECT 1353.480 651.850 1353.620 676.075 ;
        RECT 1353.480 651.710 1354.080 651.850 ;
        RECT 1353.940 627.970 1354.080 651.710 ;
        RECT 1352.960 627.650 1353.220 627.970 ;
        RECT 1353.880 627.650 1354.140 627.970 ;
        RECT 1353.020 593.370 1353.160 627.650 ;
        RECT 1353.020 593.230 1353.620 593.370 ;
        RECT 1353.480 531.490 1353.620 593.230 ;
        RECT 1353.480 531.350 1354.080 531.490 ;
        RECT 1353.940 477.205 1354.080 531.350 ;
        RECT 1353.870 476.835 1354.150 477.205 ;
        RECT 1353.410 476.155 1353.690 476.525 ;
        RECT 1353.480 451.930 1353.620 476.155 ;
        RECT 1353.020 451.790 1353.620 451.930 ;
        RECT 1353.020 434.510 1353.160 451.790 ;
        RECT 1352.960 434.190 1353.220 434.510 ;
        RECT 1354.340 434.190 1354.600 434.510 ;
        RECT 1354.400 386.570 1354.540 434.190 ;
        RECT 1353.420 386.250 1353.680 386.570 ;
        RECT 1354.340 386.250 1354.600 386.570 ;
        RECT 1353.480 379.430 1353.620 386.250 ;
        RECT 1353.420 379.110 1353.680 379.430 ;
        RECT 1353.880 331.170 1354.140 331.490 ;
        RECT 1353.940 304.290 1354.080 331.170 ;
        RECT 1353.880 303.970 1354.140 304.290 ;
        RECT 1353.420 303.290 1353.680 303.610 ;
        RECT 1353.480 235.270 1353.620 303.290 ;
        RECT 1353.420 234.950 1353.680 235.270 ;
        RECT 1352.960 234.610 1353.220 234.930 ;
        RECT 1353.020 193.530 1353.160 234.610 ;
        RECT 1353.020 193.390 1353.620 193.530 ;
        RECT 1353.480 145.170 1353.620 193.390 ;
        RECT 1353.420 144.850 1353.680 145.170 ;
        RECT 1353.880 144.850 1354.140 145.170 ;
        RECT 1353.940 138.030 1354.080 144.850 ;
        RECT 1353.880 137.710 1354.140 138.030 ;
        RECT 1353.420 89.770 1353.680 90.090 ;
        RECT 1353.480 73.770 1353.620 89.770 ;
        RECT 413.640 73.450 413.900 73.770 ;
        RECT 1353.420 73.450 1353.680 73.770 ;
        RECT 413.700 16.310 413.840 73.450 ;
        RECT 407.200 15.990 407.460 16.310 ;
        RECT 413.640 15.990 413.900 16.310 ;
        RECT 407.260 2.400 407.400 15.990 ;
        RECT 407.050 -4.800 407.610 2.400 ;
      LAYER via2 ;
        RECT 1353.870 1303.760 1354.150 1304.040 ;
        RECT 1354.790 1303.760 1355.070 1304.040 ;
        RECT 1353.410 676.120 1353.690 676.400 ;
        RECT 1354.330 676.120 1354.610 676.400 ;
        RECT 1353.870 476.880 1354.150 477.160 ;
        RECT 1353.410 476.200 1353.690 476.480 ;
      LAYER met3 ;
        RECT 1353.845 1304.050 1354.175 1304.065 ;
        RECT 1354.765 1304.050 1355.095 1304.065 ;
        RECT 1353.845 1303.750 1355.095 1304.050 ;
        RECT 1353.845 1303.735 1354.175 1303.750 ;
        RECT 1354.765 1303.735 1355.095 1303.750 ;
        RECT 1353.385 676.410 1353.715 676.425 ;
        RECT 1354.305 676.410 1354.635 676.425 ;
        RECT 1353.385 676.110 1354.635 676.410 ;
        RECT 1353.385 676.095 1353.715 676.110 ;
        RECT 1354.305 676.095 1354.635 676.110 ;
        RECT 1353.845 477.170 1354.175 477.185 ;
        RECT 1352.710 476.870 1354.175 477.170 ;
        RECT 1352.710 476.490 1353.010 476.870 ;
        RECT 1353.845 476.855 1354.175 476.870 ;
        RECT 1353.385 476.490 1353.715 476.505 ;
        RECT 1352.710 476.190 1353.715 476.490 ;
        RECT 1353.385 476.175 1353.715 476.190 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 68.150 58.720 68.470 58.780 ;
        RECT 1180.890 58.720 1181.210 58.780 ;
        RECT 68.150 58.580 1181.210 58.720 ;
        RECT 68.150 58.520 68.470 58.580 ;
        RECT 1180.890 58.520 1181.210 58.580 ;
      LAYER via ;
        RECT 68.180 58.520 68.440 58.780 ;
        RECT 1180.920 58.520 1181.180 58.780 ;
      LAYER met2 ;
        RECT 1183.600 1700.410 1183.880 1704.000 ;
        RECT 1180.980 1700.270 1183.880 1700.410 ;
        RECT 1180.980 58.810 1181.120 1700.270 ;
        RECT 1183.600 1700.000 1183.880 1700.270 ;
        RECT 68.180 58.490 68.440 58.810 ;
        RECT 1180.920 58.490 1181.180 58.810 ;
        RECT 68.240 2.400 68.380 58.490 ;
        RECT 68.030 -4.800 68.590 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 427.410 74.020 427.730 74.080 ;
        RECT 1366.730 74.020 1367.050 74.080 ;
        RECT 427.410 73.880 1367.050 74.020 ;
        RECT 427.410 73.820 427.730 73.880 ;
        RECT 1366.730 73.820 1367.050 73.880 ;
        RECT 424.650 16.220 424.970 16.280 ;
        RECT 427.410 16.220 427.730 16.280 ;
        RECT 424.650 16.080 427.730 16.220 ;
        RECT 424.650 16.020 424.970 16.080 ;
        RECT 427.410 16.020 427.730 16.080 ;
      LAYER via ;
        RECT 427.440 73.820 427.700 74.080 ;
        RECT 1366.760 73.820 1367.020 74.080 ;
        RECT 424.680 16.020 424.940 16.280 ;
        RECT 427.440 16.020 427.700 16.280 ;
      LAYER met2 ;
        RECT 1367.140 1700.410 1367.420 1704.000 ;
        RECT 1366.820 1700.270 1367.420 1700.410 ;
        RECT 1366.820 74.110 1366.960 1700.270 ;
        RECT 1367.140 1700.000 1367.420 1700.270 ;
        RECT 427.440 73.790 427.700 74.110 ;
        RECT 1366.760 73.790 1367.020 74.110 ;
        RECT 427.500 16.310 427.640 73.790 ;
        RECT 424.680 15.990 424.940 16.310 ;
        RECT 427.440 15.990 427.700 16.310 ;
        RECT 424.740 2.400 424.880 15.990 ;
        RECT 424.530 -4.800 425.090 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 448.110 74.360 448.430 74.420 ;
        RECT 1373.630 74.360 1373.950 74.420 ;
        RECT 448.110 74.220 1373.950 74.360 ;
        RECT 448.110 74.160 448.430 74.220 ;
        RECT 1373.630 74.160 1373.950 74.220 ;
        RECT 442.590 16.220 442.910 16.280 ;
        RECT 448.110 16.220 448.430 16.280 ;
        RECT 442.590 16.080 448.430 16.220 ;
        RECT 442.590 16.020 442.910 16.080 ;
        RECT 448.110 16.020 448.430 16.080 ;
      LAYER via ;
        RECT 448.140 74.160 448.400 74.420 ;
        RECT 1373.660 74.160 1373.920 74.420 ;
        RECT 442.620 16.020 442.880 16.280 ;
        RECT 448.140 16.020 448.400 16.280 ;
      LAYER met2 ;
        RECT 1376.340 1700.410 1376.620 1704.000 ;
        RECT 1373.720 1700.270 1376.620 1700.410 ;
        RECT 1373.720 74.450 1373.860 1700.270 ;
        RECT 1376.340 1700.000 1376.620 1700.270 ;
        RECT 448.140 74.130 448.400 74.450 ;
        RECT 1373.660 74.130 1373.920 74.450 ;
        RECT 448.200 16.310 448.340 74.130 ;
        RECT 442.620 15.990 442.880 16.310 ;
        RECT 448.140 15.990 448.400 16.310 ;
        RECT 442.680 2.400 442.820 15.990 ;
        RECT 442.470 -4.800 443.030 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 461.910 74.700 462.230 74.760 ;
        RECT 1380.530 74.700 1380.850 74.760 ;
        RECT 461.910 74.560 1380.850 74.700 ;
        RECT 461.910 74.500 462.230 74.560 ;
        RECT 1380.530 74.500 1380.850 74.560 ;
      LAYER via ;
        RECT 461.940 74.500 462.200 74.760 ;
        RECT 1380.560 74.500 1380.820 74.760 ;
      LAYER met2 ;
        RECT 1385.540 1700.410 1385.820 1704.000 ;
        RECT 1382.920 1700.270 1385.820 1700.410 ;
        RECT 1382.920 1678.650 1383.060 1700.270 ;
        RECT 1385.540 1700.000 1385.820 1700.270 ;
        RECT 1380.620 1678.510 1383.060 1678.650 ;
        RECT 1380.620 74.790 1380.760 1678.510 ;
        RECT 461.940 74.470 462.200 74.790 ;
        RECT 1380.560 74.470 1380.820 74.790 ;
        RECT 462.000 17.410 462.140 74.470 ;
        RECT 460.620 17.270 462.140 17.410 ;
        RECT 460.620 2.400 460.760 17.270 ;
        RECT 460.410 -4.800 460.970 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 482.610 75.040 482.930 75.100 ;
        RECT 1394.330 75.040 1394.650 75.100 ;
        RECT 482.610 74.900 1394.650 75.040 ;
        RECT 482.610 74.840 482.930 74.900 ;
        RECT 1394.330 74.840 1394.650 74.900 ;
        RECT 478.470 15.540 478.790 15.600 ;
        RECT 482.610 15.540 482.930 15.600 ;
        RECT 478.470 15.400 482.930 15.540 ;
        RECT 478.470 15.340 478.790 15.400 ;
        RECT 482.610 15.340 482.930 15.400 ;
      LAYER via ;
        RECT 482.640 74.840 482.900 75.100 ;
        RECT 1394.360 74.840 1394.620 75.100 ;
        RECT 478.500 15.340 478.760 15.600 ;
        RECT 482.640 15.340 482.900 15.600 ;
      LAYER met2 ;
        RECT 1394.740 1700.410 1395.020 1704.000 ;
        RECT 1394.420 1700.270 1395.020 1700.410 ;
        RECT 1394.420 75.130 1394.560 1700.270 ;
        RECT 1394.740 1700.000 1395.020 1700.270 ;
        RECT 482.640 74.810 482.900 75.130 ;
        RECT 1394.360 74.810 1394.620 75.130 ;
        RECT 482.700 15.630 482.840 74.810 ;
        RECT 478.500 15.310 478.760 15.630 ;
        RECT 482.640 15.310 482.900 15.630 ;
        RECT 478.560 2.400 478.700 15.310 ;
        RECT 478.350 -4.800 478.910 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 496.410 75.380 496.730 75.440 ;
        RECT 1401.230 75.380 1401.550 75.440 ;
        RECT 496.410 75.240 1401.550 75.380 ;
        RECT 496.410 75.180 496.730 75.240 ;
        RECT 1401.230 75.180 1401.550 75.240 ;
      LAYER via ;
        RECT 496.440 75.180 496.700 75.440 ;
        RECT 1401.260 75.180 1401.520 75.440 ;
      LAYER met2 ;
        RECT 1403.940 1700.410 1404.220 1704.000 ;
        RECT 1401.320 1700.270 1404.220 1700.410 ;
        RECT 1401.320 75.470 1401.460 1700.270 ;
        RECT 1403.940 1700.000 1404.220 1700.270 ;
        RECT 496.440 75.150 496.700 75.470 ;
        RECT 1401.260 75.150 1401.520 75.470 ;
        RECT 496.500 2.400 496.640 75.150 ;
        RECT 496.290 -4.800 496.850 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1408.205 1538.925 1408.375 1587.035 ;
        RECT 1408.205 1449.165 1408.375 1497.275 ;
        RECT 1409.125 1297.185 1409.295 1345.295 ;
        RECT 1408.665 1062.245 1408.835 1145.375 ;
        RECT 1409.585 965.685 1409.755 1007.335 ;
        RECT 1408.205 506.685 1408.375 531.335 ;
        RECT 1408.665 379.525 1408.835 386.495 ;
        RECT 1408.665 307.105 1408.835 337.875 ;
        RECT 1408.205 234.685 1408.375 282.795 ;
        RECT 1408.665 96.645 1408.835 144.755 ;
      LAYER mcon ;
        RECT 1408.205 1586.865 1408.375 1587.035 ;
        RECT 1408.205 1497.105 1408.375 1497.275 ;
        RECT 1409.125 1345.125 1409.295 1345.295 ;
        RECT 1408.665 1145.205 1408.835 1145.375 ;
        RECT 1409.585 1007.165 1409.755 1007.335 ;
        RECT 1408.205 531.165 1408.375 531.335 ;
        RECT 1408.665 386.325 1408.835 386.495 ;
        RECT 1408.665 337.705 1408.835 337.875 ;
        RECT 1408.205 282.625 1408.375 282.795 ;
        RECT 1408.665 144.585 1408.835 144.755 ;
      LAYER met1 ;
        RECT 1408.130 1635.300 1408.450 1635.360 ;
        RECT 1409.970 1635.300 1410.290 1635.360 ;
        RECT 1408.130 1635.160 1410.290 1635.300 ;
        RECT 1408.130 1635.100 1408.450 1635.160 ;
        RECT 1409.970 1635.100 1410.290 1635.160 ;
        RECT 1408.130 1587.020 1408.450 1587.080 ;
        RECT 1407.935 1586.880 1408.450 1587.020 ;
        RECT 1408.130 1586.820 1408.450 1586.880 ;
        RECT 1408.130 1539.080 1408.450 1539.140 ;
        RECT 1407.935 1538.940 1408.450 1539.080 ;
        RECT 1408.130 1538.880 1408.450 1538.940 ;
        RECT 1408.130 1511.340 1408.450 1511.600 ;
        RECT 1408.220 1510.520 1408.360 1511.340 ;
        RECT 1409.050 1510.520 1409.370 1510.580 ;
        RECT 1408.220 1510.380 1409.370 1510.520 ;
        RECT 1409.050 1510.320 1409.370 1510.380 ;
        RECT 1408.145 1497.260 1408.435 1497.305 ;
        RECT 1409.050 1497.260 1409.370 1497.320 ;
        RECT 1408.145 1497.120 1409.370 1497.260 ;
        RECT 1408.145 1497.075 1408.435 1497.120 ;
        RECT 1409.050 1497.060 1409.370 1497.120 ;
        RECT 1408.130 1449.320 1408.450 1449.380 ;
        RECT 1407.935 1449.180 1408.450 1449.320 ;
        RECT 1408.130 1449.120 1408.450 1449.180 ;
        RECT 1408.590 1401.040 1408.910 1401.100 ;
        RECT 1409.510 1401.040 1409.830 1401.100 ;
        RECT 1408.590 1400.900 1409.830 1401.040 ;
        RECT 1408.590 1400.840 1408.910 1400.900 ;
        RECT 1409.510 1400.840 1409.830 1400.900 ;
        RECT 1409.050 1345.280 1409.370 1345.340 ;
        RECT 1408.855 1345.140 1409.370 1345.280 ;
        RECT 1409.050 1345.080 1409.370 1345.140 ;
        RECT 1409.065 1297.340 1409.355 1297.385 ;
        RECT 1409.970 1297.340 1410.290 1297.400 ;
        RECT 1409.065 1297.200 1410.290 1297.340 ;
        RECT 1409.065 1297.155 1409.355 1297.200 ;
        RECT 1409.970 1297.140 1410.290 1297.200 ;
        RECT 1409.970 1241.920 1410.290 1241.980 ;
        RECT 1410.890 1241.920 1411.210 1241.980 ;
        RECT 1409.970 1241.780 1411.210 1241.920 ;
        RECT 1409.970 1241.720 1410.290 1241.780 ;
        RECT 1410.890 1241.720 1411.210 1241.780 ;
        RECT 1409.510 1173.580 1409.830 1173.640 ;
        RECT 1409.140 1173.440 1409.830 1173.580 ;
        RECT 1409.140 1172.960 1409.280 1173.440 ;
        RECT 1409.510 1173.380 1409.830 1173.440 ;
        RECT 1409.050 1172.700 1409.370 1172.960 ;
        RECT 1408.605 1145.360 1408.895 1145.405 ;
        RECT 1409.050 1145.360 1409.370 1145.420 ;
        RECT 1408.605 1145.220 1409.370 1145.360 ;
        RECT 1408.605 1145.175 1408.895 1145.220 ;
        RECT 1409.050 1145.160 1409.370 1145.220 ;
        RECT 1408.605 1062.400 1408.895 1062.445 ;
        RECT 1409.050 1062.400 1409.370 1062.460 ;
        RECT 1408.605 1062.260 1409.370 1062.400 ;
        RECT 1408.605 1062.215 1408.895 1062.260 ;
        RECT 1409.050 1062.200 1409.370 1062.260 ;
        RECT 1408.590 1014.460 1408.910 1014.520 ;
        RECT 1409.510 1014.460 1409.830 1014.520 ;
        RECT 1408.590 1014.320 1409.830 1014.460 ;
        RECT 1408.590 1014.260 1408.910 1014.320 ;
        RECT 1409.510 1014.260 1409.830 1014.320 ;
        RECT 1409.510 1007.320 1409.830 1007.380 ;
        RECT 1409.315 1007.180 1409.830 1007.320 ;
        RECT 1409.510 1007.120 1409.830 1007.180 ;
        RECT 1409.510 965.840 1409.830 965.900 ;
        RECT 1409.315 965.700 1409.830 965.840 ;
        RECT 1409.510 965.640 1409.830 965.700 ;
        RECT 1408.590 765.920 1408.910 765.980 ;
        RECT 1409.050 765.920 1409.370 765.980 ;
        RECT 1408.590 765.780 1409.370 765.920 ;
        RECT 1408.590 765.720 1408.910 765.780 ;
        RECT 1409.050 765.720 1409.370 765.780 ;
        RECT 1408.130 531.320 1408.450 531.380 ;
        RECT 1407.935 531.180 1408.450 531.320 ;
        RECT 1408.130 531.120 1408.450 531.180 ;
        RECT 1408.130 506.840 1408.450 506.900 ;
        RECT 1407.935 506.700 1408.450 506.840 ;
        RECT 1408.130 506.640 1408.450 506.700 ;
        RECT 1408.590 386.480 1408.910 386.540 ;
        RECT 1408.395 386.340 1408.910 386.480 ;
        RECT 1408.590 386.280 1408.910 386.340 ;
        RECT 1408.590 379.680 1408.910 379.740 ;
        RECT 1408.395 379.540 1408.910 379.680 ;
        RECT 1408.590 379.480 1408.910 379.540 ;
        RECT 1408.590 337.860 1408.910 337.920 ;
        RECT 1408.395 337.720 1408.910 337.860 ;
        RECT 1408.590 337.660 1408.910 337.720 ;
        RECT 1408.590 307.260 1408.910 307.320 ;
        RECT 1408.395 307.120 1408.910 307.260 ;
        RECT 1408.590 307.060 1408.910 307.120 ;
        RECT 1408.145 282.780 1408.435 282.825 ;
        RECT 1408.590 282.780 1408.910 282.840 ;
        RECT 1408.145 282.640 1408.910 282.780 ;
        RECT 1408.145 282.595 1408.435 282.640 ;
        RECT 1408.590 282.580 1408.910 282.640 ;
        RECT 1408.130 234.840 1408.450 234.900 ;
        RECT 1407.935 234.700 1408.450 234.840 ;
        RECT 1408.130 234.640 1408.450 234.700 ;
        RECT 1408.590 144.740 1408.910 144.800 ;
        RECT 1408.395 144.600 1408.910 144.740 ;
        RECT 1408.590 144.540 1408.910 144.600 ;
        RECT 1408.590 96.800 1408.910 96.860 ;
        RECT 1408.395 96.660 1408.910 96.800 ;
        RECT 1408.590 96.600 1408.910 96.660 ;
        RECT 517.110 80.140 517.430 80.200 ;
        RECT 1408.590 80.140 1408.910 80.200 ;
        RECT 517.110 80.000 1408.910 80.140 ;
        RECT 517.110 79.940 517.430 80.000 ;
        RECT 1408.590 79.940 1408.910 80.000 ;
        RECT 513.890 15.540 514.210 15.600 ;
        RECT 517.110 15.540 517.430 15.600 ;
        RECT 513.890 15.400 517.430 15.540 ;
        RECT 513.890 15.340 514.210 15.400 ;
        RECT 517.110 15.340 517.430 15.400 ;
      LAYER via ;
        RECT 1408.160 1635.100 1408.420 1635.360 ;
        RECT 1410.000 1635.100 1410.260 1635.360 ;
        RECT 1408.160 1586.820 1408.420 1587.080 ;
        RECT 1408.160 1538.880 1408.420 1539.140 ;
        RECT 1408.160 1511.340 1408.420 1511.600 ;
        RECT 1409.080 1510.320 1409.340 1510.580 ;
        RECT 1409.080 1497.060 1409.340 1497.320 ;
        RECT 1408.160 1449.120 1408.420 1449.380 ;
        RECT 1408.620 1400.840 1408.880 1401.100 ;
        RECT 1409.540 1400.840 1409.800 1401.100 ;
        RECT 1409.080 1345.080 1409.340 1345.340 ;
        RECT 1410.000 1297.140 1410.260 1297.400 ;
        RECT 1410.000 1241.720 1410.260 1241.980 ;
        RECT 1410.920 1241.720 1411.180 1241.980 ;
        RECT 1409.540 1173.380 1409.800 1173.640 ;
        RECT 1409.080 1172.700 1409.340 1172.960 ;
        RECT 1409.080 1145.160 1409.340 1145.420 ;
        RECT 1409.080 1062.200 1409.340 1062.460 ;
        RECT 1408.620 1014.260 1408.880 1014.520 ;
        RECT 1409.540 1014.260 1409.800 1014.520 ;
        RECT 1409.540 1007.120 1409.800 1007.380 ;
        RECT 1409.540 965.640 1409.800 965.900 ;
        RECT 1408.620 765.720 1408.880 765.980 ;
        RECT 1409.080 765.720 1409.340 765.980 ;
        RECT 1408.160 531.120 1408.420 531.380 ;
        RECT 1408.160 506.640 1408.420 506.900 ;
        RECT 1408.620 386.280 1408.880 386.540 ;
        RECT 1408.620 379.480 1408.880 379.740 ;
        RECT 1408.620 337.660 1408.880 337.920 ;
        RECT 1408.620 307.060 1408.880 307.320 ;
        RECT 1408.620 282.580 1408.880 282.840 ;
        RECT 1408.160 234.640 1408.420 234.900 ;
        RECT 1408.620 144.540 1408.880 144.800 ;
        RECT 1408.620 96.600 1408.880 96.860 ;
        RECT 517.140 79.940 517.400 80.200 ;
        RECT 1408.620 79.940 1408.880 80.200 ;
        RECT 513.920 15.340 514.180 15.600 ;
        RECT 517.140 15.340 517.400 15.600 ;
      LAYER met2 ;
        RECT 1413.140 1700.410 1413.420 1704.000 ;
        RECT 1410.520 1700.270 1413.420 1700.410 ;
        RECT 1410.520 1659.610 1410.660 1700.270 ;
        RECT 1413.140 1700.000 1413.420 1700.270 ;
        RECT 1409.600 1659.470 1410.660 1659.610 ;
        RECT 1409.600 1651.450 1409.740 1659.470 ;
        RECT 1409.600 1651.310 1410.200 1651.450 ;
        RECT 1410.060 1635.390 1410.200 1651.310 ;
        RECT 1408.160 1635.070 1408.420 1635.390 ;
        RECT 1410.000 1635.070 1410.260 1635.390 ;
        RECT 1408.220 1587.110 1408.360 1635.070 ;
        RECT 1408.160 1586.790 1408.420 1587.110 ;
        RECT 1408.160 1538.850 1408.420 1539.170 ;
        RECT 1408.220 1511.630 1408.360 1538.850 ;
        RECT 1408.160 1511.310 1408.420 1511.630 ;
        RECT 1409.080 1510.290 1409.340 1510.610 ;
        RECT 1409.140 1497.350 1409.280 1510.290 ;
        RECT 1409.080 1497.030 1409.340 1497.350 ;
        RECT 1408.160 1449.090 1408.420 1449.410 ;
        RECT 1408.220 1448.925 1408.360 1449.090 ;
        RECT 1408.150 1448.555 1408.430 1448.925 ;
        RECT 1409.530 1448.555 1409.810 1448.925 ;
        RECT 1409.600 1401.130 1409.740 1448.555 ;
        RECT 1408.620 1400.810 1408.880 1401.130 ;
        RECT 1409.540 1400.810 1409.800 1401.130 ;
        RECT 1408.680 1400.530 1408.820 1400.810 ;
        RECT 1408.680 1400.390 1409.280 1400.530 ;
        RECT 1409.140 1345.370 1409.280 1400.390 ;
        RECT 1409.080 1345.050 1409.340 1345.370 ;
        RECT 1410.000 1297.110 1410.260 1297.430 ;
        RECT 1410.060 1242.010 1410.200 1297.110 ;
        RECT 1410.000 1241.690 1410.260 1242.010 ;
        RECT 1410.920 1241.690 1411.180 1242.010 ;
        RECT 1410.980 1193.925 1411.120 1241.690 ;
        RECT 1409.530 1193.555 1409.810 1193.925 ;
        RECT 1410.910 1193.555 1411.190 1193.925 ;
        RECT 1409.600 1173.670 1409.740 1193.555 ;
        RECT 1409.540 1173.350 1409.800 1173.670 ;
        RECT 1409.080 1172.670 1409.340 1172.990 ;
        RECT 1409.140 1145.450 1409.280 1172.670 ;
        RECT 1409.080 1145.130 1409.340 1145.450 ;
        RECT 1409.080 1062.170 1409.340 1062.490 ;
        RECT 1409.140 1055.770 1409.280 1062.170 ;
        RECT 1409.140 1055.630 1409.740 1055.770 ;
        RECT 1409.600 1014.550 1409.740 1055.630 ;
        RECT 1408.620 1014.405 1408.880 1014.550 ;
        RECT 1409.540 1014.405 1409.800 1014.550 ;
        RECT 1408.610 1014.035 1408.890 1014.405 ;
        RECT 1409.530 1014.035 1409.810 1014.405 ;
        RECT 1409.600 1007.410 1409.740 1014.035 ;
        RECT 1409.540 1007.090 1409.800 1007.410 ;
        RECT 1409.540 965.610 1409.800 965.930 ;
        RECT 1409.600 959.210 1409.740 965.610 ;
        RECT 1409.600 959.070 1410.200 959.210 ;
        RECT 1410.060 918.525 1410.200 959.070 ;
        RECT 1409.990 918.155 1410.270 918.525 ;
        RECT 1409.990 916.795 1410.270 917.165 ;
        RECT 1410.060 881.690 1410.200 916.795 ;
        RECT 1409.140 881.550 1410.200 881.690 ;
        RECT 1409.140 795.330 1409.280 881.550 ;
        RECT 1408.680 795.190 1409.280 795.330 ;
        RECT 1408.680 766.010 1408.820 795.190 ;
        RECT 1408.620 765.690 1408.880 766.010 ;
        RECT 1409.080 765.690 1409.340 766.010 ;
        RECT 1409.140 594.050 1409.280 765.690 ;
        RECT 1408.680 593.910 1409.280 594.050 ;
        RECT 1408.680 545.770 1408.820 593.910 ;
        RECT 1408.680 545.630 1409.280 545.770 ;
        RECT 1409.140 531.605 1409.280 545.630 ;
        RECT 1408.150 531.235 1408.430 531.605 ;
        RECT 1409.070 531.235 1409.350 531.605 ;
        RECT 1408.160 531.090 1408.420 531.235 ;
        RECT 1408.160 506.610 1408.420 506.930 ;
        RECT 1408.220 483.210 1408.360 506.610 ;
        RECT 1408.220 483.070 1408.820 483.210 ;
        RECT 1408.680 458.730 1408.820 483.070 ;
        RECT 1408.680 458.590 1409.280 458.730 ;
        RECT 1409.140 448.530 1409.280 458.590 ;
        RECT 1408.680 448.390 1409.280 448.530 ;
        RECT 1408.680 386.570 1408.820 448.390 ;
        RECT 1408.620 386.250 1408.880 386.570 ;
        RECT 1408.620 379.450 1408.880 379.770 ;
        RECT 1408.680 337.950 1408.820 379.450 ;
        RECT 1408.620 337.630 1408.880 337.950 ;
        RECT 1408.620 307.030 1408.880 307.350 ;
        RECT 1408.680 282.870 1408.820 307.030 ;
        RECT 1408.620 282.550 1408.880 282.870 ;
        RECT 1408.160 234.610 1408.420 234.930 ;
        RECT 1408.220 234.330 1408.360 234.610 ;
        RECT 1408.220 234.190 1408.820 234.330 ;
        RECT 1408.680 144.830 1408.820 234.190 ;
        RECT 1408.620 144.510 1408.880 144.830 ;
        RECT 1408.620 96.570 1408.880 96.890 ;
        RECT 1408.680 80.230 1408.820 96.570 ;
        RECT 517.140 79.910 517.400 80.230 ;
        RECT 1408.620 79.910 1408.880 80.230 ;
        RECT 517.200 15.630 517.340 79.910 ;
        RECT 513.920 15.310 514.180 15.630 ;
        RECT 517.140 15.310 517.400 15.630 ;
        RECT 513.980 2.400 514.120 15.310 ;
        RECT 513.770 -4.800 514.330 2.400 ;
      LAYER via2 ;
        RECT 1408.150 1448.600 1408.430 1448.880 ;
        RECT 1409.530 1448.600 1409.810 1448.880 ;
        RECT 1409.530 1193.600 1409.810 1193.880 ;
        RECT 1410.910 1193.600 1411.190 1193.880 ;
        RECT 1408.610 1014.080 1408.890 1014.360 ;
        RECT 1409.530 1014.080 1409.810 1014.360 ;
        RECT 1409.990 918.200 1410.270 918.480 ;
        RECT 1409.990 916.840 1410.270 917.120 ;
        RECT 1408.150 531.280 1408.430 531.560 ;
        RECT 1409.070 531.280 1409.350 531.560 ;
      LAYER met3 ;
        RECT 1408.125 1448.890 1408.455 1448.905 ;
        RECT 1409.505 1448.890 1409.835 1448.905 ;
        RECT 1408.125 1448.590 1409.835 1448.890 ;
        RECT 1408.125 1448.575 1408.455 1448.590 ;
        RECT 1409.505 1448.575 1409.835 1448.590 ;
        RECT 1409.505 1193.890 1409.835 1193.905 ;
        RECT 1410.885 1193.890 1411.215 1193.905 ;
        RECT 1409.505 1193.590 1411.215 1193.890 ;
        RECT 1409.505 1193.575 1409.835 1193.590 ;
        RECT 1410.885 1193.575 1411.215 1193.590 ;
        RECT 1408.585 1014.370 1408.915 1014.385 ;
        RECT 1409.505 1014.370 1409.835 1014.385 ;
        RECT 1408.585 1014.070 1409.835 1014.370 ;
        RECT 1408.585 1014.055 1408.915 1014.070 ;
        RECT 1409.505 1014.055 1409.835 1014.070 ;
        RECT 1409.965 918.490 1410.295 918.505 ;
        RECT 1409.750 918.175 1410.295 918.490 ;
        RECT 1409.750 917.145 1410.050 918.175 ;
        RECT 1409.750 916.830 1410.295 917.145 ;
        RECT 1409.965 916.815 1410.295 916.830 ;
        RECT 1408.125 531.570 1408.455 531.585 ;
        RECT 1409.045 531.570 1409.375 531.585 ;
        RECT 1408.125 531.270 1409.375 531.570 ;
        RECT 1408.125 531.255 1408.455 531.270 ;
        RECT 1409.045 531.255 1409.375 531.270 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 537.810 80.480 538.130 80.540 ;
        RECT 1421.930 80.480 1422.250 80.540 ;
        RECT 537.810 80.340 1422.250 80.480 ;
        RECT 537.810 80.280 538.130 80.340 ;
        RECT 1421.930 80.280 1422.250 80.340 ;
        RECT 531.830 15.540 532.150 15.600 ;
        RECT 537.810 15.540 538.130 15.600 ;
        RECT 531.830 15.400 538.130 15.540 ;
        RECT 531.830 15.340 532.150 15.400 ;
        RECT 537.810 15.340 538.130 15.400 ;
      LAYER via ;
        RECT 537.840 80.280 538.100 80.540 ;
        RECT 1421.960 80.280 1422.220 80.540 ;
        RECT 531.860 15.340 532.120 15.600 ;
        RECT 537.840 15.340 538.100 15.600 ;
      LAYER met2 ;
        RECT 1422.340 1700.410 1422.620 1704.000 ;
        RECT 1422.020 1700.270 1422.620 1700.410 ;
        RECT 1422.020 80.570 1422.160 1700.270 ;
        RECT 1422.340 1700.000 1422.620 1700.270 ;
        RECT 537.840 80.250 538.100 80.570 ;
        RECT 1421.960 80.250 1422.220 80.570 ;
        RECT 537.900 15.630 538.040 80.250 ;
        RECT 531.860 15.310 532.120 15.630 ;
        RECT 537.840 15.310 538.100 15.630 ;
        RECT 531.920 2.400 532.060 15.310 ;
        RECT 531.710 -4.800 532.270 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 551.610 80.820 551.930 80.880 ;
        RECT 1428.830 80.820 1429.150 80.880 ;
        RECT 551.610 80.680 1429.150 80.820 ;
        RECT 551.610 80.620 551.930 80.680 ;
        RECT 1428.830 80.620 1429.150 80.680 ;
      LAYER via ;
        RECT 551.640 80.620 551.900 80.880 ;
        RECT 1428.860 80.620 1429.120 80.880 ;
      LAYER met2 ;
        RECT 1431.540 1700.410 1431.820 1704.000 ;
        RECT 1428.920 1700.270 1431.820 1700.410 ;
        RECT 1428.920 80.910 1429.060 1700.270 ;
        RECT 1431.540 1700.000 1431.820 1700.270 ;
        RECT 551.640 80.590 551.900 80.910 ;
        RECT 1428.860 80.590 1429.120 80.910 ;
        RECT 551.700 16.730 551.840 80.590 ;
        RECT 549.860 16.590 551.840 16.730 ;
        RECT 549.860 2.400 550.000 16.590 ;
        RECT 549.650 -4.800 550.210 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1436.265 1490.645 1436.435 1538.755 ;
        RECT 1436.265 669.545 1436.435 717.655 ;
        RECT 1435.805 572.645 1435.975 620.755 ;
        RECT 1435.805 428.145 1435.975 475.915 ;
        RECT 1436.265 379.525 1436.435 427.635 ;
        RECT 1436.265 283.305 1436.435 331.075 ;
        RECT 1436.265 235.025 1436.435 282.795 ;
      LAYER mcon ;
        RECT 1436.265 1538.585 1436.435 1538.755 ;
        RECT 1436.265 717.485 1436.435 717.655 ;
        RECT 1435.805 620.585 1435.975 620.755 ;
        RECT 1435.805 475.745 1435.975 475.915 ;
        RECT 1436.265 427.465 1436.435 427.635 ;
        RECT 1436.265 330.905 1436.435 331.075 ;
        RECT 1436.265 282.625 1436.435 282.795 ;
      LAYER met1 ;
        RECT 1435.730 1539.420 1436.050 1539.480 ;
        RECT 1436.650 1539.420 1436.970 1539.480 ;
        RECT 1435.730 1539.280 1436.970 1539.420 ;
        RECT 1435.730 1539.220 1436.050 1539.280 ;
        RECT 1436.650 1539.220 1436.970 1539.280 ;
        RECT 1436.205 1538.740 1436.495 1538.785 ;
        RECT 1436.650 1538.740 1436.970 1538.800 ;
        RECT 1436.205 1538.600 1436.970 1538.740 ;
        RECT 1436.205 1538.555 1436.495 1538.600 ;
        RECT 1436.650 1538.540 1436.970 1538.600 ;
        RECT 1436.190 1490.800 1436.510 1490.860 ;
        RECT 1435.995 1490.660 1436.510 1490.800 ;
        RECT 1436.190 1490.600 1436.510 1490.660 ;
        RECT 1436.190 1345.620 1436.510 1345.680 ;
        RECT 1437.110 1345.620 1437.430 1345.680 ;
        RECT 1436.190 1345.480 1437.430 1345.620 ;
        RECT 1436.190 1345.420 1436.510 1345.480 ;
        RECT 1437.110 1345.420 1437.430 1345.480 ;
        RECT 1435.730 1249.400 1436.050 1249.460 ;
        RECT 1436.650 1249.400 1436.970 1249.460 ;
        RECT 1435.730 1249.260 1436.970 1249.400 ;
        RECT 1435.730 1249.200 1436.050 1249.260 ;
        RECT 1436.650 1249.200 1436.970 1249.260 ;
        RECT 1436.190 1200.780 1436.510 1200.840 ;
        RECT 1437.110 1200.780 1437.430 1200.840 ;
        RECT 1436.190 1200.640 1437.430 1200.780 ;
        RECT 1436.190 1200.580 1436.510 1200.640 ;
        RECT 1437.110 1200.580 1437.430 1200.640 ;
        RECT 1436.190 1103.540 1436.510 1103.600 ;
        RECT 1436.650 1103.540 1436.970 1103.600 ;
        RECT 1436.190 1103.400 1436.970 1103.540 ;
        RECT 1436.190 1103.340 1436.510 1103.400 ;
        RECT 1436.650 1103.340 1436.970 1103.400 ;
        RECT 1436.650 1007.320 1436.970 1007.380 ;
        RECT 1436.650 1007.180 1437.340 1007.320 ;
        RECT 1436.650 1007.120 1436.970 1007.180 ;
        RECT 1437.200 1007.040 1437.340 1007.180 ;
        RECT 1437.110 1006.780 1437.430 1007.040 ;
        RECT 1436.190 917.900 1436.510 917.960 ;
        RECT 1437.110 917.900 1437.430 917.960 ;
        RECT 1436.190 917.760 1437.430 917.900 ;
        RECT 1436.190 917.700 1436.510 917.760 ;
        RECT 1437.110 917.700 1437.430 917.760 ;
        RECT 1436.190 910.760 1436.510 910.820 ;
        RECT 1437.110 910.760 1437.430 910.820 ;
        RECT 1436.190 910.620 1437.430 910.760 ;
        RECT 1436.190 910.560 1436.510 910.620 ;
        RECT 1437.110 910.560 1437.430 910.620 ;
        RECT 1436.190 717.640 1436.510 717.700 ;
        RECT 1435.995 717.500 1436.510 717.640 ;
        RECT 1436.190 717.440 1436.510 717.500 ;
        RECT 1436.190 669.700 1436.510 669.760 ;
        RECT 1435.995 669.560 1436.510 669.700 ;
        RECT 1436.190 669.500 1436.510 669.560 ;
        RECT 1435.745 620.740 1436.035 620.785 ;
        RECT 1436.190 620.740 1436.510 620.800 ;
        RECT 1435.745 620.600 1436.510 620.740 ;
        RECT 1435.745 620.555 1436.035 620.600 ;
        RECT 1436.190 620.540 1436.510 620.600 ;
        RECT 1435.730 572.800 1436.050 572.860 ;
        RECT 1435.535 572.660 1436.050 572.800 ;
        RECT 1435.730 572.600 1436.050 572.660 ;
        RECT 1435.745 475.900 1436.035 475.945 ;
        RECT 1436.190 475.900 1436.510 475.960 ;
        RECT 1435.745 475.760 1436.510 475.900 ;
        RECT 1435.745 475.715 1436.035 475.760 ;
        RECT 1436.190 475.700 1436.510 475.760 ;
        RECT 1435.730 428.300 1436.050 428.360 ;
        RECT 1435.535 428.160 1436.050 428.300 ;
        RECT 1435.730 428.100 1436.050 428.160 ;
        RECT 1435.730 427.620 1436.050 427.680 ;
        RECT 1436.205 427.620 1436.495 427.665 ;
        RECT 1435.730 427.480 1436.495 427.620 ;
        RECT 1435.730 427.420 1436.050 427.480 ;
        RECT 1436.205 427.435 1436.495 427.480 ;
        RECT 1436.190 379.680 1436.510 379.740 ;
        RECT 1435.995 379.540 1436.510 379.680 ;
        RECT 1436.190 379.480 1436.510 379.540 ;
        RECT 1436.190 331.540 1436.510 331.800 ;
        RECT 1436.280 331.105 1436.420 331.540 ;
        RECT 1436.205 330.875 1436.495 331.105 ;
        RECT 1436.190 283.460 1436.510 283.520 ;
        RECT 1435.995 283.320 1436.510 283.460 ;
        RECT 1436.190 283.260 1436.510 283.320 ;
        RECT 1436.190 282.780 1436.510 282.840 ;
        RECT 1435.995 282.640 1436.510 282.780 ;
        RECT 1436.190 282.580 1436.510 282.640 ;
        RECT 1436.190 235.180 1436.510 235.240 ;
        RECT 1435.995 235.040 1436.510 235.180 ;
        RECT 1436.190 234.980 1436.510 235.040 ;
        RECT 1436.190 186.560 1436.510 186.620 ;
        RECT 1436.650 186.560 1436.970 186.620 ;
        RECT 1436.190 186.420 1436.970 186.560 ;
        RECT 1436.190 186.360 1436.510 186.420 ;
        RECT 1436.650 186.360 1436.970 186.420 ;
        RECT 572.310 81.160 572.630 81.220 ;
        RECT 1436.190 81.160 1436.510 81.220 ;
        RECT 572.310 81.020 1436.510 81.160 ;
        RECT 572.310 80.960 572.630 81.020 ;
        RECT 1436.190 80.960 1436.510 81.020 ;
        RECT 567.710 14.860 568.030 14.920 ;
        RECT 572.310 14.860 572.630 14.920 ;
        RECT 567.710 14.720 572.630 14.860 ;
        RECT 567.710 14.660 568.030 14.720 ;
        RECT 572.310 14.660 572.630 14.720 ;
      LAYER via ;
        RECT 1435.760 1539.220 1436.020 1539.480 ;
        RECT 1436.680 1539.220 1436.940 1539.480 ;
        RECT 1436.680 1538.540 1436.940 1538.800 ;
        RECT 1436.220 1490.600 1436.480 1490.860 ;
        RECT 1436.220 1345.420 1436.480 1345.680 ;
        RECT 1437.140 1345.420 1437.400 1345.680 ;
        RECT 1435.760 1249.200 1436.020 1249.460 ;
        RECT 1436.680 1249.200 1436.940 1249.460 ;
        RECT 1436.220 1200.580 1436.480 1200.840 ;
        RECT 1437.140 1200.580 1437.400 1200.840 ;
        RECT 1436.220 1103.340 1436.480 1103.600 ;
        RECT 1436.680 1103.340 1436.940 1103.600 ;
        RECT 1436.680 1007.120 1436.940 1007.380 ;
        RECT 1437.140 1006.780 1437.400 1007.040 ;
        RECT 1436.220 917.700 1436.480 917.960 ;
        RECT 1437.140 917.700 1437.400 917.960 ;
        RECT 1436.220 910.560 1436.480 910.820 ;
        RECT 1437.140 910.560 1437.400 910.820 ;
        RECT 1436.220 717.440 1436.480 717.700 ;
        RECT 1436.220 669.500 1436.480 669.760 ;
        RECT 1436.220 620.540 1436.480 620.800 ;
        RECT 1435.760 572.600 1436.020 572.860 ;
        RECT 1436.220 475.700 1436.480 475.960 ;
        RECT 1435.760 428.100 1436.020 428.360 ;
        RECT 1435.760 427.420 1436.020 427.680 ;
        RECT 1436.220 379.480 1436.480 379.740 ;
        RECT 1436.220 331.540 1436.480 331.800 ;
        RECT 1436.220 283.260 1436.480 283.520 ;
        RECT 1436.220 282.580 1436.480 282.840 ;
        RECT 1436.220 234.980 1436.480 235.240 ;
        RECT 1436.220 186.360 1436.480 186.620 ;
        RECT 1436.680 186.360 1436.940 186.620 ;
        RECT 572.340 80.960 572.600 81.220 ;
        RECT 1436.220 80.960 1436.480 81.220 ;
        RECT 567.740 14.660 568.000 14.920 ;
        RECT 572.340 14.660 572.600 14.920 ;
      LAYER met2 ;
        RECT 1440.740 1700.410 1441.020 1704.000 ;
        RECT 1438.580 1700.270 1441.020 1700.410 ;
        RECT 1438.580 1689.530 1438.720 1700.270 ;
        RECT 1440.740 1700.000 1441.020 1700.270 ;
        RECT 1436.280 1689.390 1438.720 1689.530 ;
        RECT 1436.280 1618.130 1436.420 1689.390 ;
        RECT 1435.820 1617.990 1436.420 1618.130 ;
        RECT 1435.820 1539.510 1435.960 1617.990 ;
        RECT 1435.760 1539.190 1436.020 1539.510 ;
        RECT 1436.680 1539.190 1436.940 1539.510 ;
        RECT 1436.740 1538.830 1436.880 1539.190 ;
        RECT 1436.680 1538.510 1436.940 1538.830 ;
        RECT 1436.220 1490.570 1436.480 1490.890 ;
        RECT 1436.280 1393.845 1436.420 1490.570 ;
        RECT 1436.210 1393.475 1436.490 1393.845 ;
        RECT 1437.130 1393.475 1437.410 1393.845 ;
        RECT 1437.200 1345.710 1437.340 1393.475 ;
        RECT 1436.220 1345.390 1436.480 1345.710 ;
        RECT 1437.140 1345.390 1437.400 1345.710 ;
        RECT 1436.280 1297.285 1436.420 1345.390 ;
        RECT 1436.210 1296.915 1436.490 1297.285 ;
        RECT 1436.670 1296.235 1436.950 1296.605 ;
        RECT 1436.740 1249.490 1436.880 1296.235 ;
        RECT 1435.760 1249.170 1436.020 1249.490 ;
        RECT 1436.680 1249.170 1436.940 1249.490 ;
        RECT 1435.820 1249.005 1435.960 1249.170 ;
        RECT 1435.750 1248.635 1436.030 1249.005 ;
        RECT 1437.130 1248.635 1437.410 1249.005 ;
        RECT 1437.200 1200.870 1437.340 1248.635 ;
        RECT 1436.220 1200.550 1436.480 1200.870 ;
        RECT 1437.140 1200.550 1437.400 1200.870 ;
        RECT 1436.280 1103.630 1436.420 1200.550 ;
        RECT 1436.220 1103.310 1436.480 1103.630 ;
        RECT 1436.680 1103.310 1436.940 1103.630 ;
        RECT 1436.740 1056.565 1436.880 1103.310 ;
        RECT 1436.670 1056.195 1436.950 1056.565 ;
        RECT 1436.210 1055.515 1436.490 1055.885 ;
        RECT 1436.280 1031.290 1436.420 1055.515 ;
        RECT 1435.820 1031.150 1436.420 1031.290 ;
        RECT 1435.820 1007.605 1435.960 1031.150 ;
        RECT 1435.750 1007.235 1436.030 1007.605 ;
        RECT 1436.670 1007.235 1436.950 1007.605 ;
        RECT 1436.680 1007.090 1436.940 1007.235 ;
        RECT 1437.140 1006.750 1437.400 1007.070 ;
        RECT 1437.200 917.990 1437.340 1006.750 ;
        RECT 1436.220 917.670 1436.480 917.990 ;
        RECT 1437.140 917.670 1437.400 917.990 ;
        RECT 1436.280 910.850 1436.420 917.670 ;
        RECT 1436.220 910.530 1436.480 910.850 ;
        RECT 1437.140 910.530 1437.400 910.850 ;
        RECT 1437.200 862.765 1437.340 910.530 ;
        RECT 1436.210 862.395 1436.490 862.765 ;
        RECT 1437.130 862.395 1437.410 862.765 ;
        RECT 1436.280 725.405 1436.420 862.395 ;
        RECT 1436.210 725.035 1436.490 725.405 ;
        RECT 1436.210 724.355 1436.490 724.725 ;
        RECT 1436.280 717.730 1436.420 724.355 ;
        RECT 1436.220 717.410 1436.480 717.730 ;
        RECT 1436.220 669.470 1436.480 669.790 ;
        RECT 1436.280 628.845 1436.420 669.470 ;
        RECT 1436.210 628.475 1436.490 628.845 ;
        RECT 1436.210 627.795 1436.490 628.165 ;
        RECT 1436.280 620.830 1436.420 627.795 ;
        RECT 1436.220 620.510 1436.480 620.830 ;
        RECT 1435.760 572.570 1436.020 572.890 ;
        RECT 1435.820 530.810 1435.960 572.570 ;
        RECT 1435.820 530.670 1436.420 530.810 ;
        RECT 1436.280 524.010 1436.420 530.670 ;
        RECT 1436.280 523.870 1436.880 524.010 ;
        RECT 1436.740 476.410 1436.880 523.870 ;
        RECT 1436.280 476.270 1436.880 476.410 ;
        RECT 1436.280 475.990 1436.420 476.270 ;
        RECT 1436.220 475.670 1436.480 475.990 ;
        RECT 1435.760 428.070 1436.020 428.390 ;
        RECT 1435.820 427.710 1435.960 428.070 ;
        RECT 1435.760 427.390 1436.020 427.710 ;
        RECT 1436.220 379.450 1436.480 379.770 ;
        RECT 1436.280 331.830 1436.420 379.450 ;
        RECT 1436.220 331.510 1436.480 331.830 ;
        RECT 1436.220 283.230 1436.480 283.550 ;
        RECT 1436.280 282.870 1436.420 283.230 ;
        RECT 1436.220 282.550 1436.480 282.870 ;
        RECT 1436.220 234.950 1436.480 235.270 ;
        RECT 1436.280 234.500 1436.420 234.950 ;
        RECT 1436.280 234.360 1436.880 234.500 ;
        RECT 1436.740 186.650 1436.880 234.360 ;
        RECT 1436.220 186.330 1436.480 186.650 ;
        RECT 1436.680 186.330 1436.940 186.650 ;
        RECT 1436.280 186.050 1436.420 186.330 ;
        RECT 1435.820 185.910 1436.420 186.050 ;
        RECT 1435.820 158.170 1435.960 185.910 ;
        RECT 1435.820 158.030 1436.420 158.170 ;
        RECT 1436.280 81.250 1436.420 158.030 ;
        RECT 572.340 80.930 572.600 81.250 ;
        RECT 1436.220 80.930 1436.480 81.250 ;
        RECT 572.400 14.950 572.540 80.930 ;
        RECT 567.740 14.630 568.000 14.950 ;
        RECT 572.340 14.630 572.600 14.950 ;
        RECT 567.800 2.400 567.940 14.630 ;
        RECT 567.590 -4.800 568.150 2.400 ;
      LAYER via2 ;
        RECT 1436.210 1393.520 1436.490 1393.800 ;
        RECT 1437.130 1393.520 1437.410 1393.800 ;
        RECT 1436.210 1296.960 1436.490 1297.240 ;
        RECT 1436.670 1296.280 1436.950 1296.560 ;
        RECT 1435.750 1248.680 1436.030 1248.960 ;
        RECT 1437.130 1248.680 1437.410 1248.960 ;
        RECT 1436.670 1056.240 1436.950 1056.520 ;
        RECT 1436.210 1055.560 1436.490 1055.840 ;
        RECT 1435.750 1007.280 1436.030 1007.560 ;
        RECT 1436.670 1007.280 1436.950 1007.560 ;
        RECT 1436.210 862.440 1436.490 862.720 ;
        RECT 1437.130 862.440 1437.410 862.720 ;
        RECT 1436.210 725.080 1436.490 725.360 ;
        RECT 1436.210 724.400 1436.490 724.680 ;
        RECT 1436.210 628.520 1436.490 628.800 ;
        RECT 1436.210 627.840 1436.490 628.120 ;
      LAYER met3 ;
        RECT 1436.185 1393.810 1436.515 1393.825 ;
        RECT 1437.105 1393.810 1437.435 1393.825 ;
        RECT 1436.185 1393.510 1437.435 1393.810 ;
        RECT 1436.185 1393.495 1436.515 1393.510 ;
        RECT 1437.105 1393.495 1437.435 1393.510 ;
        RECT 1436.185 1297.250 1436.515 1297.265 ;
        RECT 1436.185 1296.935 1436.730 1297.250 ;
        RECT 1436.430 1296.585 1436.730 1296.935 ;
        RECT 1436.430 1296.270 1436.975 1296.585 ;
        RECT 1436.645 1296.255 1436.975 1296.270 ;
        RECT 1435.725 1248.970 1436.055 1248.985 ;
        RECT 1437.105 1248.970 1437.435 1248.985 ;
        RECT 1435.725 1248.670 1437.435 1248.970 ;
        RECT 1435.725 1248.655 1436.055 1248.670 ;
        RECT 1437.105 1248.655 1437.435 1248.670 ;
        RECT 1436.645 1056.530 1436.975 1056.545 ;
        RECT 1436.430 1056.215 1436.975 1056.530 ;
        RECT 1436.430 1055.865 1436.730 1056.215 ;
        RECT 1436.185 1055.550 1436.730 1055.865 ;
        RECT 1436.185 1055.535 1436.515 1055.550 ;
        RECT 1435.725 1007.570 1436.055 1007.585 ;
        RECT 1436.645 1007.570 1436.975 1007.585 ;
        RECT 1435.725 1007.270 1436.975 1007.570 ;
        RECT 1435.725 1007.255 1436.055 1007.270 ;
        RECT 1436.645 1007.255 1436.975 1007.270 ;
        RECT 1436.185 862.730 1436.515 862.745 ;
        RECT 1437.105 862.730 1437.435 862.745 ;
        RECT 1436.185 862.430 1437.435 862.730 ;
        RECT 1436.185 862.415 1436.515 862.430 ;
        RECT 1437.105 862.415 1437.435 862.430 ;
        RECT 1436.185 725.370 1436.515 725.385 ;
        RECT 1435.510 725.070 1436.515 725.370 ;
        RECT 1435.510 724.690 1435.810 725.070 ;
        RECT 1436.185 725.055 1436.515 725.070 ;
        RECT 1436.185 724.690 1436.515 724.705 ;
        RECT 1435.510 724.390 1436.515 724.690 ;
        RECT 1436.185 724.375 1436.515 724.390 ;
        RECT 1436.185 628.810 1436.515 628.825 ;
        RECT 1436.185 628.495 1436.730 628.810 ;
        RECT 1436.430 628.145 1436.730 628.495 ;
        RECT 1436.185 627.830 1436.730 628.145 ;
        RECT 1436.185 627.815 1436.515 627.830 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1449.990 1688.000 1450.310 1688.060 ;
        RECT 1242.160 1687.860 1450.310 1688.000 ;
        RECT 1231.490 1687.660 1231.810 1687.720 ;
        RECT 1242.160 1687.660 1242.300 1687.860 ;
        RECT 1449.990 1687.800 1450.310 1687.860 ;
        RECT 1231.490 1687.520 1242.300 1687.660 ;
        RECT 1231.490 1687.460 1231.810 1687.520 ;
        RECT 586.110 70.620 586.430 70.680 ;
        RECT 1231.490 70.620 1231.810 70.680 ;
        RECT 586.110 70.480 1231.810 70.620 ;
        RECT 586.110 70.420 586.430 70.480 ;
        RECT 1231.490 70.420 1231.810 70.480 ;
      LAYER via ;
        RECT 1231.520 1687.460 1231.780 1687.720 ;
        RECT 1450.020 1687.800 1450.280 1688.060 ;
        RECT 586.140 70.420 586.400 70.680 ;
        RECT 1231.520 70.420 1231.780 70.680 ;
      LAYER met2 ;
        RECT 1449.940 1700.000 1450.220 1704.000 ;
        RECT 1450.080 1688.090 1450.220 1700.000 ;
        RECT 1450.020 1687.770 1450.280 1688.090 ;
        RECT 1231.520 1687.430 1231.780 1687.750 ;
        RECT 1231.580 70.710 1231.720 1687.430 ;
        RECT 586.140 70.390 586.400 70.710 ;
        RECT 1231.520 70.390 1231.780 70.710 ;
        RECT 586.200 17.410 586.340 70.390 ;
        RECT 585.740 17.270 586.340 17.410 ;
        RECT 585.740 2.400 585.880 17.270 ;
        RECT 585.530 -4.800 586.090 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 96.210 65.520 96.530 65.580 ;
        RECT 1194.230 65.520 1194.550 65.580 ;
        RECT 96.210 65.380 1194.550 65.520 ;
        RECT 96.210 65.320 96.530 65.380 ;
        RECT 1194.230 65.320 1194.550 65.380 ;
        RECT 91.610 17.920 91.930 17.980 ;
        RECT 96.210 17.920 96.530 17.980 ;
        RECT 91.610 17.780 96.530 17.920 ;
        RECT 91.610 17.720 91.930 17.780 ;
        RECT 96.210 17.720 96.530 17.780 ;
      LAYER via ;
        RECT 96.240 65.320 96.500 65.580 ;
        RECT 1194.260 65.320 1194.520 65.580 ;
        RECT 91.640 17.720 91.900 17.980 ;
        RECT 96.240 17.720 96.500 17.980 ;
      LAYER met2 ;
        RECT 1195.560 1700.410 1195.840 1704.000 ;
        RECT 1194.320 1700.270 1195.840 1700.410 ;
        RECT 1194.320 65.610 1194.460 1700.270 ;
        RECT 1195.560 1700.000 1195.840 1700.270 ;
        RECT 96.240 65.290 96.500 65.610 ;
        RECT 1194.260 65.290 1194.520 65.610 ;
        RECT 96.300 18.010 96.440 65.290 ;
        RECT 91.640 17.690 91.900 18.010 ;
        RECT 96.240 17.690 96.500 18.010 ;
        RECT 91.700 2.400 91.840 17.690 ;
        RECT 91.490 -4.800 92.050 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 606.810 81.500 607.130 81.560 ;
        RECT 1456.430 81.500 1456.750 81.560 ;
        RECT 606.810 81.360 1456.750 81.500 ;
        RECT 606.810 81.300 607.130 81.360 ;
        RECT 1456.430 81.300 1456.750 81.360 ;
        RECT 603.130 14.860 603.450 14.920 ;
        RECT 606.810 14.860 607.130 14.920 ;
        RECT 603.130 14.720 607.130 14.860 ;
        RECT 603.130 14.660 603.450 14.720 ;
        RECT 606.810 14.660 607.130 14.720 ;
      LAYER via ;
        RECT 606.840 81.300 607.100 81.560 ;
        RECT 1456.460 81.300 1456.720 81.560 ;
        RECT 603.160 14.660 603.420 14.920 ;
        RECT 606.840 14.660 607.100 14.920 ;
      LAYER met2 ;
        RECT 1459.140 1700.410 1459.420 1704.000 ;
        RECT 1456.520 1700.270 1459.420 1700.410 ;
        RECT 1456.520 81.590 1456.660 1700.270 ;
        RECT 1459.140 1700.000 1459.420 1700.270 ;
        RECT 606.840 81.270 607.100 81.590 ;
        RECT 1456.460 81.270 1456.720 81.590 ;
        RECT 606.900 14.950 607.040 81.270 ;
        RECT 603.160 14.630 603.420 14.950 ;
        RECT 606.840 14.630 607.100 14.950 ;
        RECT 603.220 2.400 603.360 14.630 ;
        RECT 603.010 -4.800 603.570 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1463.865 1587.205 1464.035 1635.315 ;
        RECT 1463.405 1442.025 1463.575 1490.475 ;
        RECT 1463.405 1303.645 1463.575 1345.295 ;
        RECT 1463.865 1200.625 1464.035 1255.875 ;
        RECT 1463.865 1152.345 1464.035 1200.115 ;
        RECT 1463.865 820.845 1464.035 862.495 ;
        RECT 1463.865 737.885 1464.035 779.535 ;
        RECT 1463.865 676.345 1464.035 724.455 ;
        RECT 1463.865 627.725 1464.035 669.375 ;
        RECT 1464.325 565.845 1464.495 620.755 ;
        RECT 1463.865 235.025 1464.035 331.075 ;
        RECT 1464.325 179.605 1464.495 227.715 ;
      LAYER mcon ;
        RECT 1463.865 1635.145 1464.035 1635.315 ;
        RECT 1463.405 1490.305 1463.575 1490.475 ;
        RECT 1463.405 1345.125 1463.575 1345.295 ;
        RECT 1463.865 1255.705 1464.035 1255.875 ;
        RECT 1463.865 1199.945 1464.035 1200.115 ;
        RECT 1463.865 862.325 1464.035 862.495 ;
        RECT 1463.865 779.365 1464.035 779.535 ;
        RECT 1463.865 724.285 1464.035 724.455 ;
        RECT 1463.865 669.205 1464.035 669.375 ;
        RECT 1464.325 620.585 1464.495 620.755 ;
        RECT 1463.865 330.905 1464.035 331.075 ;
        RECT 1464.325 227.545 1464.495 227.715 ;
      LAYER met1 ;
        RECT 1463.790 1635.300 1464.110 1635.360 ;
        RECT 1463.595 1635.160 1464.110 1635.300 ;
        RECT 1463.790 1635.100 1464.110 1635.160 ;
        RECT 1463.790 1587.360 1464.110 1587.420 ;
        RECT 1463.595 1587.220 1464.110 1587.360 ;
        RECT 1463.790 1587.160 1464.110 1587.220 ;
        RECT 1463.345 1490.460 1463.635 1490.505 ;
        RECT 1463.790 1490.460 1464.110 1490.520 ;
        RECT 1463.345 1490.320 1464.110 1490.460 ;
        RECT 1463.345 1490.275 1463.635 1490.320 ;
        RECT 1463.790 1490.260 1464.110 1490.320 ;
        RECT 1463.330 1442.180 1463.650 1442.240 ;
        RECT 1463.135 1442.040 1463.650 1442.180 ;
        RECT 1463.330 1441.980 1463.650 1442.040 ;
        RECT 1463.330 1401.040 1463.650 1401.100 ;
        RECT 1463.790 1401.040 1464.110 1401.100 ;
        RECT 1463.330 1400.900 1464.110 1401.040 ;
        RECT 1463.330 1400.840 1463.650 1400.900 ;
        RECT 1463.790 1400.840 1464.110 1400.900 ;
        RECT 1463.330 1345.280 1463.650 1345.340 ;
        RECT 1463.135 1345.140 1463.650 1345.280 ;
        RECT 1463.330 1345.080 1463.650 1345.140 ;
        RECT 1463.345 1303.800 1463.635 1303.845 ;
        RECT 1463.790 1303.800 1464.110 1303.860 ;
        RECT 1463.345 1303.660 1464.110 1303.800 ;
        RECT 1463.345 1303.615 1463.635 1303.660 ;
        RECT 1463.790 1303.600 1464.110 1303.660 ;
        RECT 1463.790 1255.860 1464.110 1255.920 ;
        RECT 1463.595 1255.720 1464.110 1255.860 ;
        RECT 1463.790 1255.660 1464.110 1255.720 ;
        RECT 1463.790 1200.780 1464.110 1200.840 ;
        RECT 1463.595 1200.640 1464.110 1200.780 ;
        RECT 1463.790 1200.580 1464.110 1200.640 ;
        RECT 1463.790 1200.100 1464.110 1200.160 ;
        RECT 1463.595 1199.960 1464.110 1200.100 ;
        RECT 1463.790 1199.900 1464.110 1199.960 ;
        RECT 1463.790 1152.500 1464.110 1152.560 ;
        RECT 1463.595 1152.360 1464.110 1152.500 ;
        RECT 1463.790 1152.300 1464.110 1152.360 ;
        RECT 1463.790 1104.560 1464.110 1104.620 ;
        RECT 1463.420 1104.420 1464.110 1104.560 ;
        RECT 1463.420 1104.280 1463.560 1104.420 ;
        RECT 1463.790 1104.360 1464.110 1104.420 ;
        RECT 1463.330 1104.020 1463.650 1104.280 ;
        RECT 1463.330 1055.940 1463.650 1056.000 ;
        RECT 1463.790 1055.940 1464.110 1056.000 ;
        RECT 1463.330 1055.800 1464.110 1055.940 ;
        RECT 1463.330 1055.740 1463.650 1055.800 ;
        RECT 1463.790 1055.740 1464.110 1055.800 ;
        RECT 1463.790 1028.200 1464.110 1028.460 ;
        RECT 1463.880 1027.720 1464.020 1028.200 ;
        RECT 1464.250 1027.720 1464.570 1027.780 ;
        RECT 1463.880 1027.580 1464.570 1027.720 ;
        RECT 1464.250 1027.520 1464.570 1027.580 ;
        RECT 1463.790 966.180 1464.110 966.240 ;
        RECT 1464.710 966.180 1465.030 966.240 ;
        RECT 1463.790 966.040 1465.030 966.180 ;
        RECT 1463.790 965.980 1464.110 966.040 ;
        RECT 1464.710 965.980 1465.030 966.040 ;
        RECT 1464.250 910.760 1464.570 910.820 ;
        RECT 1464.710 910.760 1465.030 910.820 ;
        RECT 1464.250 910.620 1465.030 910.760 ;
        RECT 1464.250 910.560 1464.570 910.620 ;
        RECT 1464.710 910.560 1465.030 910.620 ;
        RECT 1463.790 862.480 1464.110 862.540 ;
        RECT 1463.595 862.340 1464.110 862.480 ;
        RECT 1463.790 862.280 1464.110 862.340 ;
        RECT 1463.790 821.000 1464.110 821.060 ;
        RECT 1463.595 820.860 1464.110 821.000 ;
        RECT 1463.790 820.800 1464.110 820.860 ;
        RECT 1463.805 779.520 1464.095 779.565 ;
        RECT 1464.250 779.520 1464.570 779.580 ;
        RECT 1463.805 779.380 1464.570 779.520 ;
        RECT 1463.805 779.335 1464.095 779.380 ;
        RECT 1464.250 779.320 1464.570 779.380 ;
        RECT 1463.790 738.040 1464.110 738.100 ;
        RECT 1463.595 737.900 1464.110 738.040 ;
        RECT 1463.790 737.840 1464.110 737.900 ;
        RECT 1463.790 724.440 1464.110 724.500 ;
        RECT 1463.595 724.300 1464.110 724.440 ;
        RECT 1463.790 724.240 1464.110 724.300 ;
        RECT 1463.790 676.500 1464.110 676.560 ;
        RECT 1463.595 676.360 1464.110 676.500 ;
        RECT 1463.790 676.300 1464.110 676.360 ;
        RECT 1463.790 669.360 1464.110 669.420 ;
        RECT 1463.595 669.220 1464.110 669.360 ;
        RECT 1463.790 669.160 1464.110 669.220 ;
        RECT 1463.790 627.880 1464.110 627.940 ;
        RECT 1463.595 627.740 1464.110 627.880 ;
        RECT 1463.790 627.680 1464.110 627.740 ;
        RECT 1464.250 620.740 1464.570 620.800 ;
        RECT 1464.055 620.600 1464.570 620.740 ;
        RECT 1464.250 620.540 1464.570 620.600 ;
        RECT 1464.265 566.000 1464.555 566.045 ;
        RECT 1464.710 566.000 1465.030 566.060 ;
        RECT 1464.265 565.860 1465.030 566.000 ;
        RECT 1464.265 565.815 1464.555 565.860 ;
        RECT 1464.710 565.800 1465.030 565.860 ;
        RECT 1463.790 524.520 1464.110 524.580 ;
        RECT 1464.710 524.520 1465.030 524.580 ;
        RECT 1463.790 524.380 1465.030 524.520 ;
        RECT 1463.790 524.320 1464.110 524.380 ;
        RECT 1464.710 524.320 1465.030 524.380 ;
        RECT 1463.790 338.200 1464.110 338.260 ;
        RECT 1464.250 338.200 1464.570 338.260 ;
        RECT 1463.790 338.060 1464.570 338.200 ;
        RECT 1463.790 338.000 1464.110 338.060 ;
        RECT 1464.250 338.000 1464.570 338.060 ;
        RECT 1463.790 331.060 1464.110 331.120 ;
        RECT 1463.595 330.920 1464.110 331.060 ;
        RECT 1463.790 330.860 1464.110 330.920 ;
        RECT 1463.805 235.180 1464.095 235.225 ;
        RECT 1464.250 235.180 1464.570 235.240 ;
        RECT 1463.805 235.040 1464.570 235.180 ;
        RECT 1463.805 234.995 1464.095 235.040 ;
        RECT 1464.250 234.980 1464.570 235.040 ;
        RECT 1464.250 227.700 1464.570 227.760 ;
        RECT 1464.055 227.560 1464.570 227.700 ;
        RECT 1464.250 227.500 1464.570 227.560 ;
        RECT 1464.250 179.760 1464.570 179.820 ;
        RECT 1464.055 179.620 1464.570 179.760 ;
        RECT 1464.250 179.560 1464.570 179.620 ;
        RECT 627.050 81.840 627.370 81.900 ;
        RECT 1463.790 81.840 1464.110 81.900 ;
        RECT 627.050 81.700 1464.110 81.840 ;
        RECT 627.050 81.640 627.370 81.700 ;
        RECT 1463.790 81.640 1464.110 81.700 ;
        RECT 621.070 20.980 621.390 21.040 ;
        RECT 627.050 20.980 627.370 21.040 ;
        RECT 621.070 20.840 627.370 20.980 ;
        RECT 621.070 20.780 621.390 20.840 ;
        RECT 627.050 20.780 627.370 20.840 ;
      LAYER via ;
        RECT 1463.820 1635.100 1464.080 1635.360 ;
        RECT 1463.820 1587.160 1464.080 1587.420 ;
        RECT 1463.820 1490.260 1464.080 1490.520 ;
        RECT 1463.360 1441.980 1463.620 1442.240 ;
        RECT 1463.360 1400.840 1463.620 1401.100 ;
        RECT 1463.820 1400.840 1464.080 1401.100 ;
        RECT 1463.360 1345.080 1463.620 1345.340 ;
        RECT 1463.820 1303.600 1464.080 1303.860 ;
        RECT 1463.820 1255.660 1464.080 1255.920 ;
        RECT 1463.820 1200.580 1464.080 1200.840 ;
        RECT 1463.820 1199.900 1464.080 1200.160 ;
        RECT 1463.820 1152.300 1464.080 1152.560 ;
        RECT 1463.820 1104.360 1464.080 1104.620 ;
        RECT 1463.360 1104.020 1463.620 1104.280 ;
        RECT 1463.360 1055.740 1463.620 1056.000 ;
        RECT 1463.820 1055.740 1464.080 1056.000 ;
        RECT 1463.820 1028.200 1464.080 1028.460 ;
        RECT 1464.280 1027.520 1464.540 1027.780 ;
        RECT 1463.820 965.980 1464.080 966.240 ;
        RECT 1464.740 965.980 1465.000 966.240 ;
        RECT 1464.280 910.560 1464.540 910.820 ;
        RECT 1464.740 910.560 1465.000 910.820 ;
        RECT 1463.820 862.280 1464.080 862.540 ;
        RECT 1463.820 820.800 1464.080 821.060 ;
        RECT 1464.280 779.320 1464.540 779.580 ;
        RECT 1463.820 737.840 1464.080 738.100 ;
        RECT 1463.820 724.240 1464.080 724.500 ;
        RECT 1463.820 676.300 1464.080 676.560 ;
        RECT 1463.820 669.160 1464.080 669.420 ;
        RECT 1463.820 627.680 1464.080 627.940 ;
        RECT 1464.280 620.540 1464.540 620.800 ;
        RECT 1464.740 565.800 1465.000 566.060 ;
        RECT 1463.820 524.320 1464.080 524.580 ;
        RECT 1464.740 524.320 1465.000 524.580 ;
        RECT 1463.820 338.000 1464.080 338.260 ;
        RECT 1464.280 338.000 1464.540 338.260 ;
        RECT 1463.820 330.860 1464.080 331.120 ;
        RECT 1464.280 234.980 1464.540 235.240 ;
        RECT 1464.280 227.500 1464.540 227.760 ;
        RECT 1464.280 179.560 1464.540 179.820 ;
        RECT 627.080 81.640 627.340 81.900 ;
        RECT 1463.820 81.640 1464.080 81.900 ;
        RECT 621.100 20.780 621.360 21.040 ;
        RECT 627.080 20.780 627.340 21.040 ;
      LAYER met2 ;
        RECT 1468.340 1700.410 1468.620 1704.000 ;
        RECT 1466.180 1700.270 1468.620 1700.410 ;
        RECT 1466.180 1636.605 1466.320 1700.270 ;
        RECT 1468.340 1700.000 1468.620 1700.270 ;
        RECT 1466.110 1636.235 1466.390 1636.605 ;
        RECT 1463.810 1635.555 1464.090 1635.925 ;
        RECT 1463.880 1635.390 1464.020 1635.555 ;
        RECT 1463.820 1635.070 1464.080 1635.390 ;
        RECT 1463.820 1587.130 1464.080 1587.450 ;
        RECT 1463.880 1490.550 1464.020 1587.130 ;
        RECT 1463.820 1490.230 1464.080 1490.550 ;
        RECT 1463.360 1441.950 1463.620 1442.270 ;
        RECT 1463.420 1401.130 1463.560 1441.950 ;
        RECT 1463.360 1400.810 1463.620 1401.130 ;
        RECT 1463.820 1400.810 1464.080 1401.130 ;
        RECT 1463.880 1371.290 1464.020 1400.810 ;
        RECT 1463.880 1371.150 1464.940 1371.290 ;
        RECT 1464.800 1346.245 1464.940 1371.150 ;
        RECT 1463.350 1345.875 1463.630 1346.245 ;
        RECT 1464.730 1345.875 1465.010 1346.245 ;
        RECT 1463.420 1345.370 1463.560 1345.875 ;
        RECT 1463.360 1345.050 1463.620 1345.370 ;
        RECT 1463.820 1303.570 1464.080 1303.890 ;
        RECT 1463.880 1255.950 1464.020 1303.570 ;
        RECT 1463.820 1255.630 1464.080 1255.950 ;
        RECT 1463.820 1200.550 1464.080 1200.870 ;
        RECT 1463.880 1200.190 1464.020 1200.550 ;
        RECT 1463.820 1199.870 1464.080 1200.190 ;
        RECT 1463.820 1152.270 1464.080 1152.590 ;
        RECT 1463.880 1104.650 1464.020 1152.270 ;
        RECT 1463.820 1104.330 1464.080 1104.650 ;
        RECT 1463.360 1103.990 1463.620 1104.310 ;
        RECT 1463.420 1056.030 1463.560 1103.990 ;
        RECT 1463.360 1055.710 1463.620 1056.030 ;
        RECT 1463.820 1055.710 1464.080 1056.030 ;
        RECT 1463.880 1028.490 1464.020 1055.710 ;
        RECT 1463.820 1028.170 1464.080 1028.490 ;
        RECT 1464.280 1027.490 1464.540 1027.810 ;
        RECT 1464.340 990.490 1464.480 1027.490 ;
        RECT 1464.340 990.350 1464.940 990.490 ;
        RECT 1464.800 966.270 1464.940 990.350 ;
        RECT 1463.820 966.125 1464.080 966.270 ;
        RECT 1464.740 966.125 1465.000 966.270 ;
        RECT 1463.810 965.755 1464.090 966.125 ;
        RECT 1464.730 965.755 1465.010 966.125 ;
        RECT 1464.800 910.850 1464.940 965.755 ;
        RECT 1464.280 910.530 1464.540 910.850 ;
        RECT 1464.740 910.530 1465.000 910.850 ;
        RECT 1464.340 862.650 1464.480 910.530 ;
        RECT 1463.880 862.570 1464.480 862.650 ;
        RECT 1463.820 862.510 1464.480 862.570 ;
        RECT 1463.820 862.250 1464.080 862.510 ;
        RECT 1463.880 862.095 1464.020 862.250 ;
        RECT 1463.820 820.770 1464.080 821.090 ;
        RECT 1463.880 814.370 1464.020 820.770 ;
        RECT 1463.880 814.230 1464.480 814.370 ;
        RECT 1464.340 779.610 1464.480 814.230 ;
        RECT 1464.280 779.290 1464.540 779.610 ;
        RECT 1463.820 737.810 1464.080 738.130 ;
        RECT 1463.880 724.530 1464.020 737.810 ;
        RECT 1463.820 724.210 1464.080 724.530 ;
        RECT 1463.820 676.270 1464.080 676.590 ;
        RECT 1463.880 669.450 1464.020 676.270 ;
        RECT 1463.820 669.130 1464.080 669.450 ;
        RECT 1463.820 627.650 1464.080 627.970 ;
        RECT 1463.880 621.250 1464.020 627.650 ;
        RECT 1463.880 621.110 1464.480 621.250 ;
        RECT 1464.340 620.830 1464.480 621.110 ;
        RECT 1464.280 620.510 1464.540 620.830 ;
        RECT 1464.740 565.770 1465.000 566.090 ;
        RECT 1464.800 524.610 1464.940 565.770 ;
        RECT 1463.820 524.290 1464.080 524.610 ;
        RECT 1464.740 524.290 1465.000 524.610 ;
        RECT 1463.880 494.090 1464.020 524.290 ;
        RECT 1463.880 493.950 1464.480 494.090 ;
        RECT 1464.340 387.330 1464.480 493.950 ;
        RECT 1463.880 387.190 1464.480 387.330 ;
        RECT 1463.880 385.970 1464.020 387.190 ;
        RECT 1463.880 385.830 1464.480 385.970 ;
        RECT 1464.340 338.290 1464.480 385.830 ;
        RECT 1463.820 337.970 1464.080 338.290 ;
        RECT 1464.280 337.970 1464.540 338.290 ;
        RECT 1463.880 331.150 1464.020 337.970 ;
        RECT 1463.820 330.830 1464.080 331.150 ;
        RECT 1464.280 234.950 1464.540 235.270 ;
        RECT 1464.340 227.790 1464.480 234.950 ;
        RECT 1464.280 227.470 1464.540 227.790 ;
        RECT 1464.280 179.530 1464.540 179.850 ;
        RECT 1464.340 152.730 1464.480 179.530 ;
        RECT 1463.880 152.590 1464.480 152.730 ;
        RECT 1463.880 81.930 1464.020 152.590 ;
        RECT 627.080 81.610 627.340 81.930 ;
        RECT 1463.820 81.610 1464.080 81.930 ;
        RECT 627.140 21.070 627.280 81.610 ;
        RECT 621.100 20.750 621.360 21.070 ;
        RECT 627.080 20.750 627.340 21.070 ;
        RECT 621.160 2.400 621.300 20.750 ;
        RECT 620.950 -4.800 621.510 2.400 ;
      LAYER via2 ;
        RECT 1466.110 1636.280 1466.390 1636.560 ;
        RECT 1463.810 1635.600 1464.090 1635.880 ;
        RECT 1463.350 1345.920 1463.630 1346.200 ;
        RECT 1464.730 1345.920 1465.010 1346.200 ;
        RECT 1463.810 965.800 1464.090 966.080 ;
        RECT 1464.730 965.800 1465.010 966.080 ;
      LAYER met3 ;
        RECT 1466.085 1636.570 1466.415 1636.585 ;
        RECT 1463.110 1636.270 1466.415 1636.570 ;
        RECT 1463.110 1635.890 1463.410 1636.270 ;
        RECT 1466.085 1636.255 1466.415 1636.270 ;
        RECT 1463.785 1635.890 1464.115 1635.905 ;
        RECT 1463.110 1635.590 1464.115 1635.890 ;
        RECT 1463.785 1635.575 1464.115 1635.590 ;
        RECT 1463.325 1346.210 1463.655 1346.225 ;
        RECT 1464.705 1346.210 1465.035 1346.225 ;
        RECT 1463.325 1345.910 1465.035 1346.210 ;
        RECT 1463.325 1345.895 1463.655 1345.910 ;
        RECT 1464.705 1345.895 1465.035 1345.910 ;
        RECT 1463.785 966.090 1464.115 966.105 ;
        RECT 1464.705 966.090 1465.035 966.105 ;
        RECT 1463.785 965.790 1465.035 966.090 ;
        RECT 1463.785 965.775 1464.115 965.790 ;
        RECT 1464.705 965.775 1465.035 965.790 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 116.910 72.320 117.230 72.380 ;
        RECT 1208.490 72.320 1208.810 72.380 ;
        RECT 116.910 72.180 1208.810 72.320 ;
        RECT 116.910 72.120 117.230 72.180 ;
        RECT 1208.490 72.120 1208.810 72.180 ;
      LAYER via ;
        RECT 116.940 72.120 117.200 72.380 ;
        RECT 1208.520 72.120 1208.780 72.380 ;
      LAYER met2 ;
        RECT 1207.980 1700.410 1208.260 1704.000 ;
        RECT 1207.980 1700.270 1208.720 1700.410 ;
        RECT 1207.980 1700.000 1208.260 1700.270 ;
        RECT 1208.580 72.410 1208.720 1700.270 ;
        RECT 116.940 72.090 117.200 72.410 ;
        RECT 1208.520 72.090 1208.780 72.410 ;
        RECT 117.000 17.410 117.140 72.090 ;
        RECT 115.620 17.270 117.140 17.410 ;
        RECT 115.620 2.400 115.760 17.270 ;
        RECT 115.410 -4.800 115.970 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1215.005 1490.985 1215.175 1538.755 ;
        RECT 1215.005 1400.885 1215.175 1490.475 ;
        RECT 1215.465 1304.325 1215.635 1352.435 ;
        RECT 1215.465 1062.585 1215.635 1110.355 ;
        RECT 1215.925 1014.305 1216.095 1028.415 ;
        RECT 1215.465 966.025 1215.635 1013.795 ;
        RECT 1215.005 814.385 1215.175 835.635 ;
        RECT 1215.005 737.885 1215.175 772.735 ;
        RECT 1216.385 620.925 1216.555 669.375 ;
        RECT 1215.465 530.825 1215.635 548.675 ;
        RECT 1215.925 338.045 1216.095 403.835 ;
      LAYER mcon ;
        RECT 1215.005 1538.585 1215.175 1538.755 ;
        RECT 1215.005 1490.305 1215.175 1490.475 ;
        RECT 1215.465 1352.265 1215.635 1352.435 ;
        RECT 1215.465 1110.185 1215.635 1110.355 ;
        RECT 1215.925 1028.245 1216.095 1028.415 ;
        RECT 1215.465 1013.625 1215.635 1013.795 ;
        RECT 1215.005 835.465 1215.175 835.635 ;
        RECT 1215.005 772.565 1215.175 772.735 ;
        RECT 1216.385 669.205 1216.555 669.375 ;
        RECT 1215.465 548.505 1215.635 548.675 ;
        RECT 1215.925 403.665 1216.095 403.835 ;
      LAYER met1 ;
        RECT 1215.390 1678.140 1215.710 1678.200 ;
        RECT 1219.070 1678.140 1219.390 1678.200 ;
        RECT 1215.390 1678.000 1219.390 1678.140 ;
        RECT 1215.390 1677.940 1215.710 1678.000 ;
        RECT 1219.070 1677.940 1219.390 1678.000 ;
        RECT 1214.945 1538.740 1215.235 1538.785 ;
        RECT 1215.390 1538.740 1215.710 1538.800 ;
        RECT 1214.945 1538.600 1215.710 1538.740 ;
        RECT 1214.945 1538.555 1215.235 1538.600 ;
        RECT 1215.390 1538.540 1215.710 1538.600 ;
        RECT 1214.930 1491.140 1215.250 1491.200 ;
        RECT 1214.735 1491.000 1215.250 1491.140 ;
        RECT 1214.930 1490.940 1215.250 1491.000 ;
        RECT 1214.930 1490.460 1215.250 1490.520 ;
        RECT 1214.735 1490.320 1215.250 1490.460 ;
        RECT 1214.930 1490.260 1215.250 1490.320 ;
        RECT 1214.945 1401.040 1215.235 1401.085 ;
        RECT 1215.850 1401.040 1216.170 1401.100 ;
        RECT 1214.945 1400.900 1216.170 1401.040 ;
        RECT 1214.945 1400.855 1215.235 1400.900 ;
        RECT 1215.850 1400.840 1216.170 1400.900 ;
        RECT 1215.390 1352.420 1215.710 1352.480 ;
        RECT 1215.195 1352.280 1215.710 1352.420 ;
        RECT 1215.390 1352.220 1215.710 1352.280 ;
        RECT 1215.405 1304.480 1215.695 1304.525 ;
        RECT 1215.850 1304.480 1216.170 1304.540 ;
        RECT 1215.405 1304.340 1216.170 1304.480 ;
        RECT 1215.405 1304.295 1215.695 1304.340 ;
        RECT 1215.850 1304.280 1216.170 1304.340 ;
        RECT 1215.390 1221.320 1215.710 1221.580 ;
        RECT 1215.480 1220.840 1215.620 1221.320 ;
        RECT 1215.850 1220.840 1216.170 1220.900 ;
        RECT 1215.480 1220.700 1216.170 1220.840 ;
        RECT 1215.850 1220.640 1216.170 1220.700 ;
        RECT 1213.550 1152.500 1213.870 1152.560 ;
        RECT 1214.010 1152.500 1214.330 1152.560 ;
        RECT 1213.550 1152.360 1214.330 1152.500 ;
        RECT 1213.550 1152.300 1213.870 1152.360 ;
        RECT 1214.010 1152.300 1214.330 1152.360 ;
        RECT 1214.010 1111.020 1214.330 1111.080 ;
        RECT 1215.850 1111.020 1216.170 1111.080 ;
        RECT 1214.010 1110.880 1216.170 1111.020 ;
        RECT 1214.010 1110.820 1214.330 1110.880 ;
        RECT 1215.850 1110.820 1216.170 1110.880 ;
        RECT 1215.390 1110.340 1215.710 1110.400 ;
        RECT 1215.195 1110.200 1215.710 1110.340 ;
        RECT 1215.390 1110.140 1215.710 1110.200 ;
        RECT 1215.405 1062.740 1215.695 1062.785 ;
        RECT 1215.850 1062.740 1216.170 1062.800 ;
        RECT 1215.405 1062.600 1216.170 1062.740 ;
        RECT 1215.405 1062.555 1215.695 1062.600 ;
        RECT 1215.850 1062.540 1216.170 1062.600 ;
        RECT 1215.850 1028.400 1216.170 1028.460 ;
        RECT 1215.655 1028.260 1216.170 1028.400 ;
        RECT 1215.850 1028.200 1216.170 1028.260 ;
        RECT 1215.850 1014.460 1216.170 1014.520 ;
        RECT 1215.655 1014.320 1216.170 1014.460 ;
        RECT 1215.850 1014.260 1216.170 1014.320 ;
        RECT 1215.390 1013.780 1215.710 1013.840 ;
        RECT 1215.195 1013.640 1215.710 1013.780 ;
        RECT 1215.390 1013.580 1215.710 1013.640 ;
        RECT 1215.405 966.180 1215.695 966.225 ;
        RECT 1215.850 966.180 1216.170 966.240 ;
        RECT 1215.405 966.040 1216.170 966.180 ;
        RECT 1215.405 965.995 1215.695 966.040 ;
        RECT 1215.850 965.980 1216.170 966.040 ;
        RECT 1215.850 931.840 1216.170 931.900 ;
        RECT 1215.480 931.700 1216.170 931.840 ;
        RECT 1215.480 931.560 1215.620 931.700 ;
        RECT 1215.850 931.640 1216.170 931.700 ;
        RECT 1215.390 931.300 1215.710 931.560 ;
        RECT 1215.850 869.620 1216.170 869.680 ;
        RECT 1216.310 869.620 1216.630 869.680 ;
        RECT 1215.850 869.480 1216.630 869.620 ;
        RECT 1215.850 869.420 1216.170 869.480 ;
        RECT 1216.310 869.420 1216.630 869.480 ;
        RECT 1214.945 835.620 1215.235 835.665 ;
        RECT 1215.850 835.620 1216.170 835.680 ;
        RECT 1214.945 835.480 1216.170 835.620 ;
        RECT 1214.945 835.435 1215.235 835.480 ;
        RECT 1215.850 835.420 1216.170 835.480 ;
        RECT 1214.930 814.540 1215.250 814.600 ;
        RECT 1214.735 814.400 1215.250 814.540 ;
        RECT 1214.930 814.340 1215.250 814.400 ;
        RECT 1214.930 772.720 1215.250 772.780 ;
        RECT 1214.735 772.580 1215.250 772.720 ;
        RECT 1214.930 772.520 1215.250 772.580 ;
        RECT 1214.945 738.040 1215.235 738.085 ;
        RECT 1215.390 738.040 1215.710 738.100 ;
        RECT 1214.945 737.900 1215.710 738.040 ;
        RECT 1214.945 737.855 1215.235 737.900 ;
        RECT 1215.390 737.840 1215.710 737.900 ;
        RECT 1215.850 724.440 1216.170 724.500 ;
        RECT 1216.310 724.440 1216.630 724.500 ;
        RECT 1215.850 724.300 1216.630 724.440 ;
        RECT 1215.850 724.240 1216.170 724.300 ;
        RECT 1216.310 724.240 1216.630 724.300 ;
        RECT 1215.390 676.160 1215.710 676.220 ;
        RECT 1216.310 676.160 1216.630 676.220 ;
        RECT 1215.390 676.020 1216.630 676.160 ;
        RECT 1215.390 675.960 1215.710 676.020 ;
        RECT 1216.310 675.960 1216.630 676.020 ;
        RECT 1216.310 669.360 1216.630 669.420 ;
        RECT 1216.115 669.220 1216.630 669.360 ;
        RECT 1216.310 669.160 1216.630 669.220 ;
        RECT 1216.325 621.080 1216.615 621.125 ;
        RECT 1216.770 621.080 1217.090 621.140 ;
        RECT 1216.325 620.940 1217.090 621.080 ;
        RECT 1216.325 620.895 1216.615 620.940 ;
        RECT 1216.770 620.880 1217.090 620.940 ;
        RECT 1215.850 572.800 1216.170 572.860 ;
        RECT 1216.770 572.800 1217.090 572.860 ;
        RECT 1215.850 572.660 1217.090 572.800 ;
        RECT 1215.850 572.600 1216.170 572.660 ;
        RECT 1216.770 572.600 1217.090 572.660 ;
        RECT 1215.390 548.660 1215.710 548.720 ;
        RECT 1215.195 548.520 1215.710 548.660 ;
        RECT 1215.390 548.460 1215.710 548.520 ;
        RECT 1215.405 530.980 1215.695 531.025 ;
        RECT 1216.310 530.980 1216.630 531.040 ;
        RECT 1215.405 530.840 1216.630 530.980 ;
        RECT 1215.405 530.795 1215.695 530.840 ;
        RECT 1216.310 530.780 1216.630 530.840 ;
        RECT 1214.930 458.900 1215.250 458.960 ;
        RECT 1217.230 458.900 1217.550 458.960 ;
        RECT 1214.930 458.760 1217.550 458.900 ;
        RECT 1214.930 458.700 1215.250 458.760 ;
        RECT 1217.230 458.700 1217.550 458.760 ;
        RECT 1215.865 403.820 1216.155 403.865 ;
        RECT 1216.770 403.820 1217.090 403.880 ;
        RECT 1215.865 403.680 1217.090 403.820 ;
        RECT 1215.865 403.635 1216.155 403.680 ;
        RECT 1216.770 403.620 1217.090 403.680 ;
        RECT 1215.850 338.200 1216.170 338.260 ;
        RECT 1215.655 338.060 1216.170 338.200 ;
        RECT 1215.850 338.000 1216.170 338.060 ;
        RECT 1215.390 144.740 1215.710 144.800 ;
        RECT 1215.850 144.740 1216.170 144.800 ;
        RECT 1215.390 144.600 1216.170 144.740 ;
        RECT 1215.390 144.540 1215.710 144.600 ;
        RECT 1215.850 144.540 1216.170 144.600 ;
        RECT 144.510 79.460 144.830 79.520 ;
        RECT 1215.390 79.460 1215.710 79.520 ;
        RECT 144.510 79.320 1215.710 79.460 ;
        RECT 144.510 79.260 144.830 79.320 ;
        RECT 1215.390 79.260 1215.710 79.320 ;
        RECT 139.450 15.880 139.770 15.940 ;
        RECT 144.510 15.880 144.830 15.940 ;
        RECT 139.450 15.740 144.830 15.880 ;
        RECT 139.450 15.680 139.770 15.740 ;
        RECT 144.510 15.680 144.830 15.740 ;
      LAYER via ;
        RECT 1215.420 1677.940 1215.680 1678.200 ;
        RECT 1219.100 1677.940 1219.360 1678.200 ;
        RECT 1215.420 1538.540 1215.680 1538.800 ;
        RECT 1214.960 1490.940 1215.220 1491.200 ;
        RECT 1214.960 1490.260 1215.220 1490.520 ;
        RECT 1215.880 1400.840 1216.140 1401.100 ;
        RECT 1215.420 1352.220 1215.680 1352.480 ;
        RECT 1215.880 1304.280 1216.140 1304.540 ;
        RECT 1215.420 1221.320 1215.680 1221.580 ;
        RECT 1215.880 1220.640 1216.140 1220.900 ;
        RECT 1213.580 1152.300 1213.840 1152.560 ;
        RECT 1214.040 1152.300 1214.300 1152.560 ;
        RECT 1214.040 1110.820 1214.300 1111.080 ;
        RECT 1215.880 1110.820 1216.140 1111.080 ;
        RECT 1215.420 1110.140 1215.680 1110.400 ;
        RECT 1215.880 1062.540 1216.140 1062.800 ;
        RECT 1215.880 1028.200 1216.140 1028.460 ;
        RECT 1215.880 1014.260 1216.140 1014.520 ;
        RECT 1215.420 1013.580 1215.680 1013.840 ;
        RECT 1215.880 965.980 1216.140 966.240 ;
        RECT 1215.880 931.640 1216.140 931.900 ;
        RECT 1215.420 931.300 1215.680 931.560 ;
        RECT 1215.880 869.420 1216.140 869.680 ;
        RECT 1216.340 869.420 1216.600 869.680 ;
        RECT 1215.880 835.420 1216.140 835.680 ;
        RECT 1214.960 814.340 1215.220 814.600 ;
        RECT 1214.960 772.520 1215.220 772.780 ;
        RECT 1215.420 737.840 1215.680 738.100 ;
        RECT 1215.880 724.240 1216.140 724.500 ;
        RECT 1216.340 724.240 1216.600 724.500 ;
        RECT 1215.420 675.960 1215.680 676.220 ;
        RECT 1216.340 675.960 1216.600 676.220 ;
        RECT 1216.340 669.160 1216.600 669.420 ;
        RECT 1216.800 620.880 1217.060 621.140 ;
        RECT 1215.880 572.600 1216.140 572.860 ;
        RECT 1216.800 572.600 1217.060 572.860 ;
        RECT 1215.420 548.460 1215.680 548.720 ;
        RECT 1216.340 530.780 1216.600 531.040 ;
        RECT 1214.960 458.700 1215.220 458.960 ;
        RECT 1217.260 458.700 1217.520 458.960 ;
        RECT 1216.800 403.620 1217.060 403.880 ;
        RECT 1215.880 338.000 1216.140 338.260 ;
        RECT 1215.420 144.540 1215.680 144.800 ;
        RECT 1215.880 144.540 1216.140 144.800 ;
        RECT 144.540 79.260 144.800 79.520 ;
        RECT 1215.420 79.260 1215.680 79.520 ;
        RECT 139.480 15.680 139.740 15.940 ;
        RECT 144.540 15.680 144.800 15.940 ;
      LAYER met2 ;
        RECT 1220.400 1700.410 1220.680 1704.000 ;
        RECT 1219.160 1700.270 1220.680 1700.410 ;
        RECT 1219.160 1678.230 1219.300 1700.270 ;
        RECT 1220.400 1700.000 1220.680 1700.270 ;
        RECT 1215.420 1677.910 1215.680 1678.230 ;
        RECT 1219.100 1677.910 1219.360 1678.230 ;
        RECT 1215.480 1538.830 1215.620 1677.910 ;
        RECT 1215.420 1538.510 1215.680 1538.830 ;
        RECT 1214.960 1490.910 1215.220 1491.230 ;
        RECT 1215.020 1490.550 1215.160 1490.910 ;
        RECT 1214.960 1490.230 1215.220 1490.550 ;
        RECT 1215.880 1400.810 1216.140 1401.130 ;
        RECT 1215.940 1400.645 1216.080 1400.810 ;
        RECT 1215.870 1400.275 1216.150 1400.645 ;
        RECT 1216.790 1400.275 1217.070 1400.645 ;
        RECT 1216.860 1353.725 1217.000 1400.275 ;
        RECT 1216.790 1353.355 1217.070 1353.725 ;
        RECT 1215.410 1352.675 1215.690 1353.045 ;
        RECT 1215.480 1352.510 1215.620 1352.675 ;
        RECT 1215.420 1352.190 1215.680 1352.510 ;
        RECT 1215.880 1304.250 1216.140 1304.570 ;
        RECT 1215.940 1304.085 1216.080 1304.250 ;
        RECT 1215.870 1303.715 1216.150 1304.085 ;
        RECT 1216.790 1303.715 1217.070 1304.085 ;
        RECT 1216.860 1257.165 1217.000 1303.715 ;
        RECT 1216.790 1256.795 1217.070 1257.165 ;
        RECT 1215.410 1256.115 1215.690 1256.485 ;
        RECT 1215.480 1221.610 1215.620 1256.115 ;
        RECT 1215.420 1221.290 1215.680 1221.610 ;
        RECT 1215.880 1220.610 1216.140 1220.930 ;
        RECT 1215.940 1207.410 1216.080 1220.610 ;
        RECT 1215.020 1207.270 1216.080 1207.410 ;
        RECT 1215.020 1200.725 1215.160 1207.270 ;
        RECT 1213.570 1200.355 1213.850 1200.725 ;
        RECT 1214.950 1200.355 1215.230 1200.725 ;
        RECT 1213.640 1152.590 1213.780 1200.355 ;
        RECT 1213.580 1152.270 1213.840 1152.590 ;
        RECT 1214.040 1152.270 1214.300 1152.590 ;
        RECT 1214.100 1111.110 1214.240 1152.270 ;
        RECT 1215.940 1111.110 1216.080 1111.265 ;
        RECT 1214.040 1110.790 1214.300 1111.110 ;
        RECT 1215.880 1110.850 1216.140 1111.110 ;
        RECT 1215.480 1110.790 1216.140 1110.850 ;
        RECT 1215.480 1110.710 1216.080 1110.790 ;
        RECT 1215.480 1110.430 1215.620 1110.710 ;
        RECT 1215.420 1110.110 1215.680 1110.430 ;
        RECT 1215.880 1062.510 1216.140 1062.830 ;
        RECT 1215.940 1028.490 1216.080 1062.510 ;
        RECT 1215.880 1028.170 1216.140 1028.490 ;
        RECT 1215.940 1014.550 1216.080 1014.705 ;
        RECT 1215.880 1014.290 1216.140 1014.550 ;
        RECT 1215.480 1014.230 1216.140 1014.290 ;
        RECT 1215.480 1014.150 1216.080 1014.230 ;
        RECT 1215.480 1013.870 1215.620 1014.150 ;
        RECT 1215.420 1013.550 1215.680 1013.870 ;
        RECT 1215.880 965.950 1216.140 966.270 ;
        RECT 1215.940 931.930 1216.080 965.950 ;
        RECT 1215.880 931.610 1216.140 931.930 ;
        RECT 1215.420 931.270 1215.680 931.590 ;
        RECT 1215.480 918.525 1215.620 931.270 ;
        RECT 1215.410 918.155 1215.690 918.525 ;
        RECT 1216.330 917.475 1216.610 917.845 ;
        RECT 1216.400 869.710 1216.540 917.475 ;
        RECT 1215.880 869.390 1216.140 869.710 ;
        RECT 1216.340 869.390 1216.600 869.710 ;
        RECT 1215.940 835.710 1216.080 869.390 ;
        RECT 1215.880 835.390 1216.140 835.710 ;
        RECT 1214.960 814.310 1215.220 814.630 ;
        RECT 1215.020 772.810 1215.160 814.310 ;
        RECT 1214.960 772.490 1215.220 772.810 ;
        RECT 1215.420 737.810 1215.680 738.130 ;
        RECT 1215.480 724.610 1215.620 737.810 ;
        RECT 1215.480 724.530 1216.080 724.610 ;
        RECT 1215.480 724.470 1216.140 724.530 ;
        RECT 1215.880 724.210 1216.140 724.470 ;
        RECT 1216.340 724.210 1216.600 724.530 ;
        RECT 1216.400 676.445 1216.540 724.210 ;
        RECT 1215.410 676.075 1215.690 676.445 ;
        RECT 1216.330 676.075 1216.610 676.445 ;
        RECT 1215.420 675.930 1215.680 676.075 ;
        RECT 1216.340 675.930 1216.600 676.075 ;
        RECT 1216.400 669.450 1216.540 675.930 ;
        RECT 1216.340 669.130 1216.600 669.450 ;
        RECT 1216.800 620.850 1217.060 621.170 ;
        RECT 1216.860 572.890 1217.000 620.850 ;
        RECT 1215.880 572.800 1216.140 572.890 ;
        RECT 1215.480 572.660 1216.140 572.800 ;
        RECT 1215.480 548.750 1215.620 572.660 ;
        RECT 1215.880 572.570 1216.140 572.660 ;
        RECT 1216.800 572.570 1217.060 572.890 ;
        RECT 1215.420 548.430 1215.680 548.750 ;
        RECT 1216.340 530.750 1216.600 531.070 ;
        RECT 1216.400 496.810 1216.540 530.750 ;
        RECT 1215.020 496.670 1216.540 496.810 ;
        RECT 1215.020 458.990 1215.160 496.670 ;
        RECT 1214.960 458.670 1215.220 458.990 ;
        RECT 1217.260 458.670 1217.520 458.990 ;
        RECT 1217.320 434.930 1217.460 458.670 ;
        RECT 1216.860 434.790 1217.460 434.930 ;
        RECT 1216.860 403.910 1217.000 434.790 ;
        RECT 1216.800 403.590 1217.060 403.910 ;
        RECT 1215.880 337.970 1216.140 338.290 ;
        RECT 1215.940 207.130 1216.080 337.970 ;
        RECT 1215.480 206.990 1216.080 207.130 ;
        RECT 1215.480 169.050 1215.620 206.990 ;
        RECT 1215.020 168.910 1215.620 169.050 ;
        RECT 1215.020 158.170 1215.160 168.910 ;
        RECT 1215.020 158.030 1216.080 158.170 ;
        RECT 1215.940 144.830 1216.080 158.030 ;
        RECT 1215.420 144.510 1215.680 144.830 ;
        RECT 1215.880 144.510 1216.140 144.830 ;
        RECT 1215.480 79.550 1215.620 144.510 ;
        RECT 144.540 79.230 144.800 79.550 ;
        RECT 1215.420 79.230 1215.680 79.550 ;
        RECT 144.600 15.970 144.740 79.230 ;
        RECT 139.480 15.650 139.740 15.970 ;
        RECT 144.540 15.650 144.800 15.970 ;
        RECT 139.540 2.400 139.680 15.650 ;
        RECT 139.330 -4.800 139.890 2.400 ;
      LAYER via2 ;
        RECT 1215.870 1400.320 1216.150 1400.600 ;
        RECT 1216.790 1400.320 1217.070 1400.600 ;
        RECT 1216.790 1353.400 1217.070 1353.680 ;
        RECT 1215.410 1352.720 1215.690 1353.000 ;
        RECT 1215.870 1303.760 1216.150 1304.040 ;
        RECT 1216.790 1303.760 1217.070 1304.040 ;
        RECT 1216.790 1256.840 1217.070 1257.120 ;
        RECT 1215.410 1256.160 1215.690 1256.440 ;
        RECT 1213.570 1200.400 1213.850 1200.680 ;
        RECT 1214.950 1200.400 1215.230 1200.680 ;
        RECT 1215.410 918.200 1215.690 918.480 ;
        RECT 1216.330 917.520 1216.610 917.800 ;
        RECT 1215.410 676.120 1215.690 676.400 ;
        RECT 1216.330 676.120 1216.610 676.400 ;
      LAYER met3 ;
        RECT 1215.845 1400.610 1216.175 1400.625 ;
        RECT 1216.765 1400.610 1217.095 1400.625 ;
        RECT 1215.845 1400.310 1217.095 1400.610 ;
        RECT 1215.845 1400.295 1216.175 1400.310 ;
        RECT 1216.765 1400.295 1217.095 1400.310 ;
        RECT 1216.765 1353.690 1217.095 1353.705 ;
        RECT 1214.710 1353.390 1217.095 1353.690 ;
        RECT 1214.710 1353.010 1215.010 1353.390 ;
        RECT 1216.765 1353.375 1217.095 1353.390 ;
        RECT 1215.385 1353.010 1215.715 1353.025 ;
        RECT 1214.710 1352.710 1215.715 1353.010 ;
        RECT 1215.385 1352.695 1215.715 1352.710 ;
        RECT 1215.845 1304.050 1216.175 1304.065 ;
        RECT 1216.765 1304.050 1217.095 1304.065 ;
        RECT 1215.845 1303.750 1217.095 1304.050 ;
        RECT 1215.845 1303.735 1216.175 1303.750 ;
        RECT 1216.765 1303.735 1217.095 1303.750 ;
        RECT 1216.765 1257.130 1217.095 1257.145 ;
        RECT 1214.710 1256.830 1217.095 1257.130 ;
        RECT 1214.710 1256.450 1215.010 1256.830 ;
        RECT 1216.765 1256.815 1217.095 1256.830 ;
        RECT 1215.385 1256.450 1215.715 1256.465 ;
        RECT 1214.710 1256.150 1215.715 1256.450 ;
        RECT 1215.385 1256.135 1215.715 1256.150 ;
        RECT 1213.545 1200.690 1213.875 1200.705 ;
        RECT 1214.925 1200.690 1215.255 1200.705 ;
        RECT 1213.545 1200.390 1215.255 1200.690 ;
        RECT 1213.545 1200.375 1213.875 1200.390 ;
        RECT 1214.925 1200.375 1215.255 1200.390 ;
        RECT 1215.385 918.490 1215.715 918.505 ;
        RECT 1215.385 918.175 1215.930 918.490 ;
        RECT 1215.630 917.810 1215.930 918.175 ;
        RECT 1216.305 917.810 1216.635 917.825 ;
        RECT 1215.630 917.510 1216.635 917.810 ;
        RECT 1216.305 917.495 1216.635 917.510 ;
        RECT 1215.385 676.410 1215.715 676.425 ;
        RECT 1216.305 676.410 1216.635 676.425 ;
        RECT 1215.385 676.110 1216.635 676.410 ;
        RECT 1215.385 676.095 1215.715 676.110 ;
        RECT 1216.305 676.095 1216.635 676.110 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 158.310 79.800 158.630 79.860 ;
        RECT 1228.730 79.800 1229.050 79.860 ;
        RECT 158.310 79.660 1229.050 79.800 ;
        RECT 158.310 79.600 158.630 79.660 ;
        RECT 1228.730 79.600 1229.050 79.660 ;
      LAYER via ;
        RECT 158.340 79.600 158.600 79.860 ;
        RECT 1228.760 79.600 1229.020 79.860 ;
      LAYER met2 ;
        RECT 1229.600 1700.410 1229.880 1704.000 ;
        RECT 1228.820 1700.270 1229.880 1700.410 ;
        RECT 1228.820 79.890 1228.960 1700.270 ;
        RECT 1229.600 1700.000 1229.880 1700.270 ;
        RECT 158.340 79.570 158.600 79.890 ;
        RECT 1228.760 79.570 1229.020 79.890 ;
        RECT 158.400 3.130 158.540 79.570 ;
        RECT 157.480 2.990 158.540 3.130 ;
        RECT 157.480 2.400 157.620 2.990 ;
        RECT 157.270 -4.800 157.830 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 230.990 1689.020 231.310 1689.080 ;
        RECT 1238.390 1689.020 1238.710 1689.080 ;
        RECT 230.990 1688.880 1238.710 1689.020 ;
        RECT 230.990 1688.820 231.310 1688.880 ;
        RECT 1238.390 1688.820 1238.710 1688.880 ;
        RECT 174.870 19.960 175.190 20.020 ;
        RECT 230.990 19.960 231.310 20.020 ;
        RECT 174.870 19.820 231.310 19.960 ;
        RECT 174.870 19.760 175.190 19.820 ;
        RECT 230.990 19.760 231.310 19.820 ;
      LAYER via ;
        RECT 231.020 1688.820 231.280 1689.080 ;
        RECT 1238.420 1688.820 1238.680 1689.080 ;
        RECT 174.900 19.760 175.160 20.020 ;
        RECT 231.020 19.760 231.280 20.020 ;
      LAYER met2 ;
        RECT 1238.340 1700.000 1238.620 1704.000 ;
        RECT 1238.480 1689.110 1238.620 1700.000 ;
        RECT 231.020 1688.790 231.280 1689.110 ;
        RECT 1238.420 1688.790 1238.680 1689.110 ;
        RECT 231.080 20.050 231.220 1688.790 ;
        RECT 174.900 19.730 175.160 20.050 ;
        RECT 231.020 19.730 231.280 20.050 ;
        RECT 174.960 2.400 175.100 19.730 ;
        RECT 174.750 -4.800 175.310 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1242.070 1678.140 1242.390 1678.200 ;
        RECT 1245.750 1678.140 1246.070 1678.200 ;
        RECT 1242.070 1678.000 1246.070 1678.140 ;
        RECT 1242.070 1677.940 1242.390 1678.000 ;
        RECT 1245.750 1677.940 1246.070 1678.000 ;
        RECT 192.810 19.280 193.130 19.340 ;
        RECT 1242.070 19.280 1242.390 19.340 ;
        RECT 192.810 19.140 1242.390 19.280 ;
        RECT 192.810 19.080 193.130 19.140 ;
        RECT 1242.070 19.080 1242.390 19.140 ;
      LAYER via ;
        RECT 1242.100 1677.940 1242.360 1678.200 ;
        RECT 1245.780 1677.940 1246.040 1678.200 ;
        RECT 192.840 19.080 193.100 19.340 ;
        RECT 1242.100 19.080 1242.360 19.340 ;
      LAYER met2 ;
        RECT 1247.540 1700.410 1247.820 1704.000 ;
        RECT 1245.840 1700.270 1247.820 1700.410 ;
        RECT 1245.840 1678.230 1245.980 1700.270 ;
        RECT 1247.540 1700.000 1247.820 1700.270 ;
        RECT 1242.100 1677.910 1242.360 1678.230 ;
        RECT 1245.780 1677.910 1246.040 1678.230 ;
        RECT 1242.160 19.370 1242.300 1677.910 ;
        RECT 192.840 19.050 193.100 19.370 ;
        RECT 1242.100 19.050 1242.360 19.370 ;
        RECT 192.900 2.400 193.040 19.050 ;
        RECT 192.690 -4.800 193.250 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 251.690 1689.360 252.010 1689.420 ;
        RECT 1256.790 1689.360 1257.110 1689.420 ;
        RECT 251.690 1689.220 1257.110 1689.360 ;
        RECT 251.690 1689.160 252.010 1689.220 ;
        RECT 1256.790 1689.160 1257.110 1689.220 ;
        RECT 210.750 20.640 211.070 20.700 ;
        RECT 251.690 20.640 252.010 20.700 ;
        RECT 210.750 20.500 252.010 20.640 ;
        RECT 210.750 20.440 211.070 20.500 ;
        RECT 251.690 20.440 252.010 20.500 ;
      LAYER via ;
        RECT 251.720 1689.160 251.980 1689.420 ;
        RECT 1256.820 1689.160 1257.080 1689.420 ;
        RECT 210.780 20.440 211.040 20.700 ;
        RECT 251.720 20.440 251.980 20.700 ;
      LAYER met2 ;
        RECT 1256.740 1700.000 1257.020 1704.000 ;
        RECT 1256.880 1689.450 1257.020 1700.000 ;
        RECT 251.720 1689.130 251.980 1689.450 ;
        RECT 1256.820 1689.130 1257.080 1689.450 ;
        RECT 251.780 20.730 251.920 1689.130 ;
        RECT 210.780 20.410 211.040 20.730 ;
        RECT 251.720 20.410 251.980 20.730 ;
        RECT 210.840 2.400 210.980 20.410 ;
        RECT 210.630 -4.800 211.190 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1259.090 1686.640 1259.410 1686.700 ;
        RECT 1265.990 1686.640 1266.310 1686.700 ;
        RECT 1259.090 1686.500 1266.310 1686.640 ;
        RECT 1259.090 1686.440 1259.410 1686.500 ;
        RECT 1265.990 1686.440 1266.310 1686.500 ;
        RECT 228.690 19.620 229.010 19.680 ;
        RECT 1259.090 19.620 1259.410 19.680 ;
        RECT 228.690 19.480 1259.410 19.620 ;
        RECT 228.690 19.420 229.010 19.480 ;
        RECT 1259.090 19.420 1259.410 19.480 ;
      LAYER via ;
        RECT 1259.120 1686.440 1259.380 1686.700 ;
        RECT 1266.020 1686.440 1266.280 1686.700 ;
        RECT 228.720 19.420 228.980 19.680 ;
        RECT 1259.120 19.420 1259.380 19.680 ;
      LAYER met2 ;
        RECT 1265.940 1700.000 1266.220 1704.000 ;
        RECT 1266.080 1686.730 1266.220 1700.000 ;
        RECT 1259.120 1686.410 1259.380 1686.730 ;
        RECT 1266.020 1686.410 1266.280 1686.730 ;
        RECT 1259.180 19.710 1259.320 1686.410 ;
        RECT 228.720 19.390 228.980 19.710 ;
        RECT 1259.120 19.390 1259.380 19.710 ;
        RECT 228.780 2.400 228.920 19.390 ;
        RECT 228.570 -4.800 229.130 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1140.870 1687.660 1141.190 1687.720 ;
        RECT 1174.450 1687.660 1174.770 1687.720 ;
        RECT 1140.870 1687.520 1174.770 1687.660 ;
        RECT 1140.870 1687.460 1141.190 1687.520 ;
        RECT 1174.450 1687.460 1174.770 1687.520 ;
        RECT 79.190 1686.980 79.510 1687.040 ;
        RECT 1140.870 1686.980 1141.190 1687.040 ;
        RECT 79.190 1686.840 1141.190 1686.980 ;
        RECT 79.190 1686.780 79.510 1686.840 ;
        RECT 1140.870 1686.780 1141.190 1686.840 ;
        RECT 50.210 15.200 50.530 15.260 ;
        RECT 79.190 15.200 79.510 15.260 ;
        RECT 50.210 15.060 79.510 15.200 ;
        RECT 50.210 15.000 50.530 15.060 ;
        RECT 79.190 15.000 79.510 15.060 ;
      LAYER via ;
        RECT 1140.900 1687.460 1141.160 1687.720 ;
        RECT 1174.480 1687.460 1174.740 1687.720 ;
        RECT 79.220 1686.780 79.480 1687.040 ;
        RECT 1140.900 1686.780 1141.160 1687.040 ;
        RECT 50.240 15.000 50.500 15.260 ;
        RECT 79.220 15.000 79.480 15.260 ;
      LAYER met2 ;
        RECT 1174.400 1700.000 1174.680 1704.000 ;
        RECT 1174.540 1687.750 1174.680 1700.000 ;
        RECT 1140.900 1687.430 1141.160 1687.750 ;
        RECT 1174.480 1687.430 1174.740 1687.750 ;
        RECT 1140.960 1687.070 1141.100 1687.430 ;
        RECT 79.220 1686.750 79.480 1687.070 ;
        RECT 1140.900 1686.750 1141.160 1687.070 ;
        RECT 79.280 15.290 79.420 1686.750 ;
        RECT 50.240 14.970 50.500 15.290 ;
        RECT 79.220 14.970 79.480 15.290 ;
        RECT 50.300 2.400 50.440 14.970 ;
        RECT 50.090 -4.800 50.650 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1266.910 1688.340 1267.230 1688.400 ;
        RECT 1278.410 1688.340 1278.730 1688.400 ;
        RECT 1266.910 1688.200 1278.730 1688.340 ;
        RECT 1266.910 1688.140 1267.230 1688.200 ;
        RECT 1278.410 1688.140 1278.730 1688.200 ;
        RECT 252.610 20.300 252.930 20.360 ;
        RECT 1265.990 20.300 1266.310 20.360 ;
        RECT 252.610 20.160 1266.310 20.300 ;
        RECT 252.610 20.100 252.930 20.160 ;
        RECT 1265.990 20.100 1266.310 20.160 ;
      LAYER via ;
        RECT 1266.940 1688.140 1267.200 1688.400 ;
        RECT 1278.440 1688.140 1278.700 1688.400 ;
        RECT 252.640 20.100 252.900 20.360 ;
        RECT 1266.020 20.100 1266.280 20.360 ;
      LAYER met2 ;
        RECT 1278.360 1700.000 1278.640 1704.000 ;
        RECT 1278.500 1688.430 1278.640 1700.000 ;
        RECT 1266.940 1688.110 1267.200 1688.430 ;
        RECT 1278.440 1688.110 1278.700 1688.430 ;
        RECT 1267.000 1672.530 1267.140 1688.110 ;
        RECT 1266.080 1672.390 1267.140 1672.530 ;
        RECT 1266.080 20.390 1266.220 1672.390 ;
        RECT 252.640 20.070 252.900 20.390 ;
        RECT 1266.020 20.070 1266.280 20.390 ;
        RECT 252.700 2.400 252.840 20.070 ;
        RECT 252.490 -4.800 253.050 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 286.190 1689.700 286.510 1689.760 ;
        RECT 1287.610 1689.700 1287.930 1689.760 ;
        RECT 286.190 1689.560 1287.930 1689.700 ;
        RECT 286.190 1689.500 286.510 1689.560 ;
        RECT 1287.610 1689.500 1287.930 1689.560 ;
        RECT 270.090 16.560 270.410 16.620 ;
        RECT 286.190 16.560 286.510 16.620 ;
        RECT 270.090 16.420 286.510 16.560 ;
        RECT 270.090 16.360 270.410 16.420 ;
        RECT 286.190 16.360 286.510 16.420 ;
      LAYER via ;
        RECT 286.220 1689.500 286.480 1689.760 ;
        RECT 1287.640 1689.500 1287.900 1689.760 ;
        RECT 270.120 16.360 270.380 16.620 ;
        RECT 286.220 16.360 286.480 16.620 ;
      LAYER met2 ;
        RECT 1287.560 1700.000 1287.840 1704.000 ;
        RECT 1287.700 1689.790 1287.840 1700.000 ;
        RECT 286.220 1689.470 286.480 1689.790 ;
        RECT 1287.640 1689.470 1287.900 1689.790 ;
        RECT 286.280 16.650 286.420 1689.470 ;
        RECT 270.120 16.330 270.380 16.650 ;
        RECT 286.220 16.330 286.480 16.650 ;
        RECT 270.180 2.400 270.320 16.330 ;
        RECT 269.970 -4.800 270.530 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1279.790 1686.640 1280.110 1686.700 ;
        RECT 1296.810 1686.640 1297.130 1686.700 ;
        RECT 1279.790 1686.500 1297.130 1686.640 ;
        RECT 1279.790 1686.440 1280.110 1686.500 ;
        RECT 1296.810 1686.440 1297.130 1686.500 ;
        RECT 288.030 20.640 288.350 20.700 ;
        RECT 1279.790 20.640 1280.110 20.700 ;
        RECT 288.030 20.500 1280.110 20.640 ;
        RECT 288.030 20.440 288.350 20.500 ;
        RECT 1279.790 20.440 1280.110 20.500 ;
      LAYER via ;
        RECT 1279.820 1686.440 1280.080 1686.700 ;
        RECT 1296.840 1686.440 1297.100 1686.700 ;
        RECT 288.060 20.440 288.320 20.700 ;
        RECT 1279.820 20.440 1280.080 20.700 ;
      LAYER met2 ;
        RECT 1296.760 1700.000 1297.040 1704.000 ;
        RECT 1296.900 1686.730 1297.040 1700.000 ;
        RECT 1279.820 1686.410 1280.080 1686.730 ;
        RECT 1296.840 1686.410 1297.100 1686.730 ;
        RECT 1279.880 20.730 1280.020 1686.410 ;
        RECT 288.060 20.410 288.320 20.730 ;
        RECT 1279.820 20.410 1280.080 20.730 ;
        RECT 288.120 2.400 288.260 20.410 ;
        RECT 287.910 -4.800 288.470 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 334.490 1690.040 334.810 1690.100 ;
        RECT 1306.010 1690.040 1306.330 1690.100 ;
        RECT 334.490 1689.900 1306.330 1690.040 ;
        RECT 334.490 1689.840 334.810 1689.900 ;
        RECT 1306.010 1689.840 1306.330 1689.900 ;
        RECT 305.970 15.880 306.290 15.940 ;
        RECT 334.490 15.880 334.810 15.940 ;
        RECT 305.970 15.740 334.810 15.880 ;
        RECT 305.970 15.680 306.290 15.740 ;
        RECT 334.490 15.680 334.810 15.740 ;
      LAYER via ;
        RECT 334.520 1689.840 334.780 1690.100 ;
        RECT 1306.040 1689.840 1306.300 1690.100 ;
        RECT 306.000 15.680 306.260 15.940 ;
        RECT 334.520 15.680 334.780 15.940 ;
      LAYER met2 ;
        RECT 1305.960 1700.000 1306.240 1704.000 ;
        RECT 1306.100 1690.130 1306.240 1700.000 ;
        RECT 334.520 1689.810 334.780 1690.130 ;
        RECT 1306.040 1689.810 1306.300 1690.130 ;
        RECT 334.580 15.970 334.720 1689.810 ;
        RECT 306.000 15.650 306.260 15.970 ;
        RECT 334.520 15.650 334.780 15.970 ;
        RECT 306.060 2.400 306.200 15.650 ;
        RECT 305.850 -4.800 306.410 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1286.690 1686.980 1287.010 1687.040 ;
        RECT 1315.210 1686.980 1315.530 1687.040 ;
        RECT 1286.690 1686.840 1315.530 1686.980 ;
        RECT 1286.690 1686.780 1287.010 1686.840 ;
        RECT 1315.210 1686.780 1315.530 1686.840 ;
        RECT 1286.690 16.900 1287.010 16.960 ;
        RECT 358.960 16.760 1287.010 16.900 ;
        RECT 323.910 16.220 324.230 16.280 ;
        RECT 358.960 16.220 359.100 16.760 ;
        RECT 1286.690 16.700 1287.010 16.760 ;
        RECT 323.910 16.080 359.100 16.220 ;
        RECT 323.910 16.020 324.230 16.080 ;
      LAYER via ;
        RECT 1286.720 1686.780 1286.980 1687.040 ;
        RECT 1315.240 1686.780 1315.500 1687.040 ;
        RECT 323.940 16.020 324.200 16.280 ;
        RECT 1286.720 16.700 1286.980 16.960 ;
      LAYER met2 ;
        RECT 1315.160 1700.000 1315.440 1704.000 ;
        RECT 1315.300 1687.070 1315.440 1700.000 ;
        RECT 1286.720 1686.750 1286.980 1687.070 ;
        RECT 1315.240 1686.750 1315.500 1687.070 ;
        RECT 1286.780 16.990 1286.920 1686.750 ;
        RECT 1286.720 16.670 1286.980 16.990 ;
        RECT 323.940 15.990 324.200 16.310 ;
        RECT 324.000 2.400 324.140 15.990 ;
        RECT 323.790 -4.800 324.350 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 355.190 1690.380 355.510 1690.440 ;
        RECT 1324.410 1690.380 1324.730 1690.440 ;
        RECT 355.190 1690.240 1324.730 1690.380 ;
        RECT 355.190 1690.180 355.510 1690.240 ;
        RECT 1324.410 1690.180 1324.730 1690.240 ;
        RECT 341.390 15.200 341.710 15.260 ;
        RECT 355.190 15.200 355.510 15.260 ;
        RECT 341.390 15.060 355.510 15.200 ;
        RECT 341.390 15.000 341.710 15.060 ;
        RECT 355.190 15.000 355.510 15.060 ;
      LAYER via ;
        RECT 355.220 1690.180 355.480 1690.440 ;
        RECT 1324.440 1690.180 1324.700 1690.440 ;
        RECT 341.420 15.000 341.680 15.260 ;
        RECT 355.220 15.000 355.480 15.260 ;
      LAYER met2 ;
        RECT 1324.360 1700.000 1324.640 1704.000 ;
        RECT 1324.500 1690.470 1324.640 1700.000 ;
        RECT 355.220 1690.150 355.480 1690.470 ;
        RECT 1324.440 1690.150 1324.700 1690.470 ;
        RECT 355.280 15.290 355.420 1690.150 ;
        RECT 341.420 14.970 341.680 15.290 ;
        RECT 355.220 14.970 355.480 15.290 ;
        RECT 341.480 2.400 341.620 14.970 ;
        RECT 341.270 -4.800 341.830 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1293.590 1688.680 1293.910 1688.740 ;
        RECT 1333.610 1688.680 1333.930 1688.740 ;
        RECT 1293.590 1688.540 1333.930 1688.680 ;
        RECT 1293.590 1688.480 1293.910 1688.540 ;
        RECT 1333.610 1688.480 1333.930 1688.540 ;
        RECT 359.330 16.560 359.650 16.620 ;
        RECT 1293.590 16.560 1293.910 16.620 ;
        RECT 359.330 16.420 1293.910 16.560 ;
        RECT 359.330 16.360 359.650 16.420 ;
        RECT 1293.590 16.360 1293.910 16.420 ;
      LAYER via ;
        RECT 1293.620 1688.480 1293.880 1688.740 ;
        RECT 1333.640 1688.480 1333.900 1688.740 ;
        RECT 359.360 16.360 359.620 16.620 ;
        RECT 1293.620 16.360 1293.880 16.620 ;
      LAYER met2 ;
        RECT 1333.560 1700.000 1333.840 1704.000 ;
        RECT 1333.700 1688.770 1333.840 1700.000 ;
        RECT 1293.620 1688.450 1293.880 1688.770 ;
        RECT 1333.640 1688.450 1333.900 1688.770 ;
        RECT 1293.680 16.650 1293.820 1688.450 ;
        RECT 359.360 16.330 359.620 16.650 ;
        RECT 1293.620 16.330 1293.880 16.650 ;
        RECT 359.420 2.400 359.560 16.330 ;
        RECT 359.210 -4.800 359.770 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 534.590 1683.920 534.910 1683.980 ;
        RECT 1342.810 1683.920 1343.130 1683.980 ;
        RECT 534.590 1683.780 1335.220 1683.920 ;
        RECT 534.590 1683.720 534.910 1683.780 ;
        RECT 1335.080 1683.580 1335.220 1683.780 ;
        RECT 1338.300 1683.780 1343.130 1683.920 ;
        RECT 1338.300 1683.580 1338.440 1683.780 ;
        RECT 1342.810 1683.720 1343.130 1683.780 ;
        RECT 1335.080 1683.440 1338.440 1683.580 ;
        RECT 534.590 14.860 534.910 14.920 ;
        RECT 502.020 14.720 534.910 14.860 ;
        RECT 377.270 14.520 377.590 14.580 ;
        RECT 502.020 14.520 502.160 14.720 ;
        RECT 534.590 14.660 534.910 14.720 ;
        RECT 377.270 14.380 502.160 14.520 ;
        RECT 377.270 14.320 377.590 14.380 ;
      LAYER via ;
        RECT 534.620 1683.720 534.880 1683.980 ;
        RECT 1342.840 1683.720 1343.100 1683.980 ;
        RECT 377.300 14.320 377.560 14.580 ;
        RECT 534.620 14.660 534.880 14.920 ;
      LAYER met2 ;
        RECT 1342.760 1700.000 1343.040 1704.000 ;
        RECT 1342.900 1684.010 1343.040 1700.000 ;
        RECT 534.620 1683.690 534.880 1684.010 ;
        RECT 1342.840 1683.690 1343.100 1684.010 ;
        RECT 534.680 14.950 534.820 1683.690 ;
        RECT 534.620 14.630 534.880 14.950 ;
        RECT 377.300 14.290 377.560 14.610 ;
        RECT 377.360 2.400 377.500 14.290 ;
        RECT 377.150 -4.800 377.710 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 414.605 14.705 414.775 15.895 ;
      LAYER mcon ;
        RECT 414.605 15.725 414.775 15.895 ;
      LAYER met1 ;
        RECT 1307.390 1687.320 1307.710 1687.380 ;
        RECT 1307.390 1687.180 1320.960 1687.320 ;
        RECT 1307.390 1687.120 1307.710 1687.180 ;
        RECT 1320.820 1686.640 1320.960 1687.180 ;
        RECT 1352.010 1686.640 1352.330 1686.700 ;
        RECT 1320.820 1686.500 1352.330 1686.640 ;
        RECT 1352.010 1686.440 1352.330 1686.500 ;
        RECT 1307.390 16.220 1307.710 16.280 ;
        RECT 448.660 16.080 1307.710 16.220 ;
        RECT 414.545 15.880 414.835 15.925 ;
        RECT 448.660 15.880 448.800 16.080 ;
        RECT 1307.390 16.020 1307.710 16.080 ;
        RECT 414.545 15.740 448.800 15.880 ;
        RECT 414.545 15.695 414.835 15.740 ;
        RECT 395.210 14.860 395.530 14.920 ;
        RECT 414.545 14.860 414.835 14.905 ;
        RECT 395.210 14.720 414.835 14.860 ;
        RECT 395.210 14.660 395.530 14.720 ;
        RECT 414.545 14.675 414.835 14.720 ;
      LAYER via ;
        RECT 1307.420 1687.120 1307.680 1687.380 ;
        RECT 1352.040 1686.440 1352.300 1686.700 ;
        RECT 1307.420 16.020 1307.680 16.280 ;
        RECT 395.240 14.660 395.500 14.920 ;
      LAYER met2 ;
        RECT 1351.960 1700.000 1352.240 1704.000 ;
        RECT 1307.420 1687.090 1307.680 1687.410 ;
        RECT 1307.480 16.310 1307.620 1687.090 ;
        RECT 1352.100 1686.730 1352.240 1700.000 ;
        RECT 1352.040 1686.410 1352.300 1686.730 ;
        RECT 1307.420 15.990 1307.680 16.310 ;
        RECT 395.240 14.630 395.500 14.950 ;
        RECT 395.300 2.400 395.440 14.630 ;
        RECT 395.090 -4.800 395.650 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 424.190 1686.300 424.510 1686.360 ;
        RECT 1361.210 1686.300 1361.530 1686.360 ;
        RECT 424.190 1686.160 1361.530 1686.300 ;
        RECT 424.190 1686.100 424.510 1686.160 ;
        RECT 1361.210 1686.100 1361.530 1686.160 ;
        RECT 424.190 16.220 424.510 16.280 ;
        RECT 414.160 16.080 424.510 16.220 ;
        RECT 413.150 15.880 413.470 15.940 ;
        RECT 414.160 15.880 414.300 16.080 ;
        RECT 424.190 16.020 424.510 16.080 ;
        RECT 413.150 15.740 414.300 15.880 ;
        RECT 413.150 15.680 413.470 15.740 ;
      LAYER via ;
        RECT 424.220 1686.100 424.480 1686.360 ;
        RECT 1361.240 1686.100 1361.500 1686.360 ;
        RECT 413.180 15.680 413.440 15.940 ;
        RECT 424.220 16.020 424.480 16.280 ;
      LAYER met2 ;
        RECT 1361.160 1700.000 1361.440 1704.000 ;
        RECT 1361.300 1686.390 1361.440 1700.000 ;
        RECT 424.220 1686.070 424.480 1686.390 ;
        RECT 1361.240 1686.070 1361.500 1686.390 ;
        RECT 424.280 16.310 424.420 1686.070 ;
        RECT 424.220 15.990 424.480 16.310 ;
        RECT 413.180 15.650 413.440 15.970 ;
        RECT 413.240 2.400 413.380 15.650 ;
        RECT 413.030 -4.800 413.590 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1182.345 1421.625 1182.515 1462.595 ;
        RECT 1180.965 1318.265 1181.135 1365.695 ;
        RECT 1181.425 1221.705 1181.595 1269.475 ;
        RECT 1181.425 1173.085 1181.595 1221.195 ;
        RECT 1181.425 1076.525 1181.595 1124.295 ;
        RECT 1181.425 890.205 1181.595 937.975 ;
        RECT 1181.885 717.145 1182.055 758.795 ;
        RECT 1181.425 517.565 1181.595 565.675 ;
        RECT 1181.425 427.805 1181.595 475.915 ;
        RECT 1181.425 379.525 1181.595 427.295 ;
        RECT 1181.425 186.405 1181.595 234.515 ;
        RECT 1181.885 83.045 1182.055 131.155 ;
      LAYER mcon ;
        RECT 1182.345 1462.425 1182.515 1462.595 ;
        RECT 1180.965 1365.525 1181.135 1365.695 ;
        RECT 1181.425 1269.305 1181.595 1269.475 ;
        RECT 1181.425 1221.025 1181.595 1221.195 ;
        RECT 1181.425 1124.125 1181.595 1124.295 ;
        RECT 1181.425 937.805 1181.595 937.975 ;
        RECT 1181.885 758.625 1182.055 758.795 ;
        RECT 1181.425 565.505 1181.595 565.675 ;
        RECT 1181.425 475.745 1181.595 475.915 ;
        RECT 1181.425 427.125 1181.595 427.295 ;
        RECT 1181.425 234.345 1181.595 234.515 ;
        RECT 1181.885 130.985 1182.055 131.155 ;
      LAYER met1 ;
        RECT 1181.350 1642.440 1181.670 1642.500 ;
        RECT 1184.570 1642.440 1184.890 1642.500 ;
        RECT 1181.350 1642.300 1184.890 1642.440 ;
        RECT 1181.350 1642.240 1181.670 1642.300 ;
        RECT 1184.570 1642.240 1184.890 1642.300 ;
        RECT 1181.350 1594.160 1181.670 1594.220 ;
        RECT 1181.810 1594.160 1182.130 1594.220 ;
        RECT 1181.350 1594.020 1182.130 1594.160 ;
        RECT 1181.350 1593.960 1181.670 1594.020 ;
        RECT 1181.810 1593.960 1182.130 1594.020 ;
        RECT 1181.810 1524.800 1182.130 1524.860 ;
        RECT 1182.730 1524.800 1183.050 1524.860 ;
        RECT 1181.810 1524.660 1183.050 1524.800 ;
        RECT 1181.810 1524.600 1182.130 1524.660 ;
        RECT 1182.730 1524.600 1183.050 1524.660 ;
        RECT 1181.350 1476.520 1181.670 1476.580 ;
        RECT 1182.270 1476.520 1182.590 1476.580 ;
        RECT 1181.350 1476.380 1182.590 1476.520 ;
        RECT 1181.350 1476.320 1181.670 1476.380 ;
        RECT 1182.270 1476.320 1182.590 1476.380 ;
        RECT 1182.270 1462.580 1182.590 1462.640 ;
        RECT 1182.075 1462.440 1182.590 1462.580 ;
        RECT 1182.270 1462.380 1182.590 1462.440 ;
        RECT 1182.270 1421.780 1182.590 1421.840 ;
        RECT 1182.075 1421.640 1182.590 1421.780 ;
        RECT 1182.270 1421.580 1182.590 1421.640 ;
        RECT 1181.350 1366.160 1181.670 1366.420 ;
        RECT 1180.905 1365.680 1181.195 1365.725 ;
        RECT 1181.440 1365.680 1181.580 1366.160 ;
        RECT 1180.905 1365.540 1181.580 1365.680 ;
        RECT 1180.905 1365.495 1181.195 1365.540 ;
        RECT 1180.905 1318.420 1181.195 1318.465 ;
        RECT 1180.905 1318.280 1181.580 1318.420 ;
        RECT 1180.905 1318.235 1181.195 1318.280 ;
        RECT 1179.970 1317.740 1180.290 1317.800 ;
        RECT 1181.440 1317.740 1181.580 1318.280 ;
        RECT 1179.970 1317.600 1181.580 1317.740 ;
        RECT 1179.970 1317.540 1180.290 1317.600 ;
        RECT 1181.350 1269.460 1181.670 1269.520 ;
        RECT 1181.155 1269.320 1181.670 1269.460 ;
        RECT 1181.350 1269.260 1181.670 1269.320 ;
        RECT 1181.365 1221.675 1181.655 1221.905 ;
        RECT 1181.440 1221.225 1181.580 1221.675 ;
        RECT 1181.365 1220.995 1181.655 1221.225 ;
        RECT 1181.350 1173.240 1181.670 1173.300 ;
        RECT 1181.155 1173.100 1181.670 1173.240 ;
        RECT 1181.350 1173.040 1181.670 1173.100 ;
        RECT 1181.350 1125.440 1181.670 1125.700 ;
        RECT 1181.440 1125.020 1181.580 1125.440 ;
        RECT 1181.350 1124.760 1181.670 1125.020 ;
        RECT 1181.350 1124.280 1181.670 1124.340 ;
        RECT 1181.155 1124.140 1181.670 1124.280 ;
        RECT 1181.350 1124.080 1181.670 1124.140 ;
        RECT 1181.350 1076.680 1181.670 1076.740 ;
        RECT 1181.155 1076.540 1181.670 1076.680 ;
        RECT 1181.350 1076.480 1181.670 1076.540 ;
        RECT 1181.810 1035.200 1182.130 1035.260 ;
        RECT 1181.810 1035.060 1183.420 1035.200 ;
        RECT 1181.810 1035.000 1182.130 1035.060 ;
        RECT 1183.280 1034.580 1183.420 1035.060 ;
        RECT 1183.190 1034.320 1183.510 1034.580 ;
        RECT 1182.270 993.040 1182.590 993.100 ;
        RECT 1183.190 993.040 1183.510 993.100 ;
        RECT 1182.270 992.900 1183.510 993.040 ;
        RECT 1182.270 992.840 1182.590 992.900 ;
        RECT 1183.190 992.840 1183.510 992.900 ;
        RECT 1181.350 938.640 1181.670 938.700 ;
        RECT 1182.270 938.640 1182.590 938.700 ;
        RECT 1181.350 938.500 1182.590 938.640 ;
        RECT 1181.350 938.440 1181.670 938.500 ;
        RECT 1182.270 938.440 1182.590 938.500 ;
        RECT 1181.350 937.960 1181.670 938.020 ;
        RECT 1181.155 937.820 1181.670 937.960 ;
        RECT 1181.350 937.760 1181.670 937.820 ;
        RECT 1181.365 890.360 1181.655 890.405 ;
        RECT 1182.270 890.360 1182.590 890.420 ;
        RECT 1181.365 890.220 1182.590 890.360 ;
        RECT 1181.365 890.175 1181.655 890.220 ;
        RECT 1182.270 890.160 1182.590 890.220 ;
        RECT 1181.810 758.780 1182.130 758.840 ;
        RECT 1181.615 758.640 1182.130 758.780 ;
        RECT 1181.810 758.580 1182.130 758.640 ;
        RECT 1181.810 717.300 1182.130 717.360 ;
        RECT 1181.615 717.160 1182.130 717.300 ;
        RECT 1181.810 717.100 1182.130 717.160 ;
        RECT 1181.350 628.700 1181.670 628.960 ;
        RECT 1181.440 628.280 1181.580 628.700 ;
        RECT 1181.350 628.020 1181.670 628.280 ;
        RECT 1181.350 590.140 1181.670 590.200 ;
        RECT 1182.270 590.140 1182.590 590.200 ;
        RECT 1181.350 590.000 1182.590 590.140 ;
        RECT 1181.350 589.940 1181.670 590.000 ;
        RECT 1182.270 589.940 1182.590 590.000 ;
        RECT 1181.365 565.660 1181.655 565.705 ;
        RECT 1181.810 565.660 1182.130 565.720 ;
        RECT 1181.365 565.520 1182.130 565.660 ;
        RECT 1181.365 565.475 1181.655 565.520 ;
        RECT 1181.810 565.460 1182.130 565.520 ;
        RECT 1181.350 517.720 1181.670 517.780 ;
        RECT 1181.155 517.580 1181.670 517.720 ;
        RECT 1181.350 517.520 1181.670 517.580 ;
        RECT 1181.350 515.680 1181.670 515.740 ;
        RECT 1182.270 515.680 1182.590 515.740 ;
        RECT 1181.350 515.540 1182.590 515.680 ;
        RECT 1181.350 515.480 1181.670 515.540 ;
        RECT 1182.270 515.480 1182.590 515.540 ;
        RECT 1181.365 475.900 1181.655 475.945 ;
        RECT 1181.810 475.900 1182.130 475.960 ;
        RECT 1181.365 475.760 1182.130 475.900 ;
        RECT 1181.365 475.715 1181.655 475.760 ;
        RECT 1181.810 475.700 1182.130 475.760 ;
        RECT 1181.350 427.960 1181.670 428.020 ;
        RECT 1181.155 427.820 1181.670 427.960 ;
        RECT 1181.350 427.760 1181.670 427.820 ;
        RECT 1181.350 427.280 1181.670 427.340 ;
        RECT 1181.155 427.140 1181.670 427.280 ;
        RECT 1181.350 427.080 1181.670 427.140 ;
        RECT 1181.365 379.680 1181.655 379.725 ;
        RECT 1181.810 379.680 1182.130 379.740 ;
        RECT 1181.365 379.540 1182.130 379.680 ;
        RECT 1181.365 379.495 1181.655 379.540 ;
        RECT 1181.810 379.480 1182.130 379.540 ;
        RECT 1181.810 339.220 1182.130 339.280 ;
        RECT 1181.440 339.080 1182.130 339.220 ;
        RECT 1181.440 337.920 1181.580 339.080 ;
        RECT 1181.810 339.020 1182.130 339.080 ;
        RECT 1181.350 337.660 1181.670 337.920 ;
        RECT 1181.810 241.980 1182.130 242.040 ;
        RECT 1181.440 241.840 1182.130 241.980 ;
        RECT 1181.440 241.700 1181.580 241.840 ;
        RECT 1181.810 241.780 1182.130 241.840 ;
        RECT 1181.350 241.440 1181.670 241.700 ;
        RECT 1181.350 234.500 1181.670 234.560 ;
        RECT 1181.155 234.360 1181.670 234.500 ;
        RECT 1181.350 234.300 1181.670 234.360 ;
        RECT 1181.365 186.560 1181.655 186.605 ;
        RECT 1181.810 186.560 1182.130 186.620 ;
        RECT 1181.365 186.420 1182.130 186.560 ;
        RECT 1181.365 186.375 1181.655 186.420 ;
        RECT 1181.810 186.360 1182.130 186.420 ;
        RECT 1181.810 131.140 1182.130 131.200 ;
        RECT 1181.615 131.000 1182.130 131.140 ;
        RECT 1181.810 130.940 1182.130 131.000 ;
        RECT 1181.810 83.200 1182.130 83.260 ;
        RECT 1181.615 83.060 1182.130 83.200 ;
        RECT 1181.810 83.000 1182.130 83.060 ;
        RECT 74.130 17.240 74.450 17.300 ;
        RECT 1181.810 17.240 1182.130 17.300 ;
        RECT 74.130 17.100 1182.130 17.240 ;
        RECT 74.130 17.040 74.450 17.100 ;
        RECT 1181.810 17.040 1182.130 17.100 ;
      LAYER via ;
        RECT 1181.380 1642.240 1181.640 1642.500 ;
        RECT 1184.600 1642.240 1184.860 1642.500 ;
        RECT 1181.380 1593.960 1181.640 1594.220 ;
        RECT 1181.840 1593.960 1182.100 1594.220 ;
        RECT 1181.840 1524.600 1182.100 1524.860 ;
        RECT 1182.760 1524.600 1183.020 1524.860 ;
        RECT 1181.380 1476.320 1181.640 1476.580 ;
        RECT 1182.300 1476.320 1182.560 1476.580 ;
        RECT 1182.300 1462.380 1182.560 1462.640 ;
        RECT 1182.300 1421.580 1182.560 1421.840 ;
        RECT 1181.380 1366.160 1181.640 1366.420 ;
        RECT 1180.000 1317.540 1180.260 1317.800 ;
        RECT 1181.380 1269.260 1181.640 1269.520 ;
        RECT 1181.380 1173.040 1181.640 1173.300 ;
        RECT 1181.380 1125.440 1181.640 1125.700 ;
        RECT 1181.380 1124.760 1181.640 1125.020 ;
        RECT 1181.380 1124.080 1181.640 1124.340 ;
        RECT 1181.380 1076.480 1181.640 1076.740 ;
        RECT 1181.840 1035.000 1182.100 1035.260 ;
        RECT 1183.220 1034.320 1183.480 1034.580 ;
        RECT 1182.300 992.840 1182.560 993.100 ;
        RECT 1183.220 992.840 1183.480 993.100 ;
        RECT 1181.380 938.440 1181.640 938.700 ;
        RECT 1182.300 938.440 1182.560 938.700 ;
        RECT 1181.380 937.760 1181.640 938.020 ;
        RECT 1182.300 890.160 1182.560 890.420 ;
        RECT 1181.840 758.580 1182.100 758.840 ;
        RECT 1181.840 717.100 1182.100 717.360 ;
        RECT 1181.380 628.700 1181.640 628.960 ;
        RECT 1181.380 628.020 1181.640 628.280 ;
        RECT 1181.380 589.940 1181.640 590.200 ;
        RECT 1182.300 589.940 1182.560 590.200 ;
        RECT 1181.840 565.460 1182.100 565.720 ;
        RECT 1181.380 517.520 1181.640 517.780 ;
        RECT 1181.380 515.480 1181.640 515.740 ;
        RECT 1182.300 515.480 1182.560 515.740 ;
        RECT 1181.840 475.700 1182.100 475.960 ;
        RECT 1181.380 427.760 1181.640 428.020 ;
        RECT 1181.380 427.080 1181.640 427.340 ;
        RECT 1181.840 379.480 1182.100 379.740 ;
        RECT 1181.840 339.020 1182.100 339.280 ;
        RECT 1181.380 337.660 1181.640 337.920 ;
        RECT 1181.840 241.780 1182.100 242.040 ;
        RECT 1181.380 241.440 1181.640 241.700 ;
        RECT 1181.380 234.300 1181.640 234.560 ;
        RECT 1181.840 186.360 1182.100 186.620 ;
        RECT 1181.840 130.940 1182.100 131.200 ;
        RECT 1181.840 83.000 1182.100 83.260 ;
        RECT 74.160 17.040 74.420 17.300 ;
        RECT 1181.840 17.040 1182.100 17.300 ;
      LAYER met2 ;
        RECT 1186.360 1700.410 1186.640 1704.000 ;
        RECT 1184.660 1700.270 1186.640 1700.410 ;
        RECT 1184.660 1642.530 1184.800 1700.270 ;
        RECT 1186.360 1700.000 1186.640 1700.270 ;
        RECT 1181.380 1642.210 1181.640 1642.530 ;
        RECT 1184.600 1642.210 1184.860 1642.530 ;
        RECT 1181.440 1594.250 1181.580 1642.210 ;
        RECT 1181.380 1593.930 1181.640 1594.250 ;
        RECT 1181.840 1593.930 1182.100 1594.250 ;
        RECT 1181.900 1524.890 1182.040 1593.930 ;
        RECT 1181.840 1524.570 1182.100 1524.890 ;
        RECT 1182.760 1524.570 1183.020 1524.890 ;
        RECT 1182.820 1476.805 1182.960 1524.570 ;
        RECT 1181.370 1476.435 1181.650 1476.805 ;
        RECT 1181.380 1476.290 1181.640 1476.435 ;
        RECT 1182.300 1476.290 1182.560 1476.610 ;
        RECT 1182.750 1476.435 1183.030 1476.805 ;
        RECT 1182.360 1462.670 1182.500 1476.290 ;
        RECT 1182.300 1462.350 1182.560 1462.670 ;
        RECT 1182.300 1421.550 1182.560 1421.870 ;
        RECT 1182.360 1380.925 1182.500 1421.550 ;
        RECT 1182.290 1380.555 1182.570 1380.925 ;
        RECT 1181.370 1379.875 1181.650 1380.245 ;
        RECT 1181.440 1366.450 1181.580 1379.875 ;
        RECT 1181.380 1366.130 1181.640 1366.450 ;
        RECT 1180.000 1317.510 1180.260 1317.830 ;
        RECT 1180.060 1270.085 1180.200 1317.510 ;
        RECT 1179.990 1269.715 1180.270 1270.085 ;
        RECT 1181.370 1269.715 1181.650 1270.085 ;
        RECT 1181.440 1269.550 1181.580 1269.715 ;
        RECT 1181.380 1269.230 1181.640 1269.550 ;
        RECT 1181.380 1173.010 1181.640 1173.330 ;
        RECT 1181.440 1125.730 1181.580 1173.010 ;
        RECT 1181.380 1125.410 1181.640 1125.730 ;
        RECT 1181.380 1124.730 1181.640 1125.050 ;
        RECT 1181.440 1124.370 1181.580 1124.730 ;
        RECT 1181.380 1124.050 1181.640 1124.370 ;
        RECT 1181.380 1076.450 1181.640 1076.770 ;
        RECT 1181.440 1076.170 1181.580 1076.450 ;
        RECT 1181.440 1076.030 1182.040 1076.170 ;
        RECT 1181.900 1035.290 1182.040 1076.030 ;
        RECT 1181.840 1034.970 1182.100 1035.290 ;
        RECT 1183.220 1034.290 1183.480 1034.610 ;
        RECT 1183.280 993.130 1183.420 1034.290 ;
        RECT 1182.300 992.810 1182.560 993.130 ;
        RECT 1183.220 992.810 1183.480 993.130 ;
        RECT 1182.360 938.730 1182.500 992.810 ;
        RECT 1181.380 938.410 1181.640 938.730 ;
        RECT 1182.300 938.410 1182.560 938.730 ;
        RECT 1181.440 938.050 1181.580 938.410 ;
        RECT 1181.380 937.730 1181.640 938.050 ;
        RECT 1182.300 890.130 1182.560 890.450 ;
        RECT 1182.360 815.165 1182.500 890.130 ;
        RECT 1182.290 814.795 1182.570 815.165 ;
        RECT 1181.370 814.370 1181.650 814.485 ;
        RECT 1181.370 814.230 1182.040 814.370 ;
        RECT 1181.370 814.115 1181.650 814.230 ;
        RECT 1181.900 758.870 1182.040 814.230 ;
        RECT 1181.840 758.550 1182.100 758.870 ;
        RECT 1181.840 717.070 1182.100 717.390 ;
        RECT 1181.900 670.325 1182.040 717.070 ;
        RECT 1181.830 669.955 1182.110 670.325 ;
        RECT 1181.370 669.275 1181.650 669.645 ;
        RECT 1181.440 628.990 1181.580 669.275 ;
        RECT 1181.380 628.670 1181.640 628.990 ;
        RECT 1181.380 627.990 1181.640 628.310 ;
        RECT 1181.440 590.230 1181.580 627.990 ;
        RECT 1181.380 589.910 1181.640 590.230 ;
        RECT 1182.300 589.910 1182.560 590.230 ;
        RECT 1182.360 566.170 1182.500 589.910 ;
        RECT 1181.900 566.030 1182.500 566.170 ;
        RECT 1181.900 565.750 1182.040 566.030 ;
        RECT 1181.840 565.430 1182.100 565.750 ;
        RECT 1181.380 517.490 1181.640 517.810 ;
        RECT 1181.440 515.770 1181.580 517.490 ;
        RECT 1181.380 515.450 1181.640 515.770 ;
        RECT 1182.300 515.450 1182.560 515.770 ;
        RECT 1182.360 483.210 1182.500 515.450 ;
        RECT 1181.900 483.070 1182.500 483.210 ;
        RECT 1181.900 475.990 1182.040 483.070 ;
        RECT 1181.840 475.670 1182.100 475.990 ;
        RECT 1181.380 427.730 1181.640 428.050 ;
        RECT 1181.440 427.370 1181.580 427.730 ;
        RECT 1181.380 427.050 1181.640 427.370 ;
        RECT 1181.840 379.450 1182.100 379.770 ;
        RECT 1181.900 339.310 1182.040 379.450 ;
        RECT 1181.840 338.990 1182.100 339.310 ;
        RECT 1181.380 337.630 1181.640 337.950 ;
        RECT 1181.440 330.890 1181.580 337.630 ;
        RECT 1181.440 330.750 1182.040 330.890 ;
        RECT 1181.900 242.070 1182.040 330.750 ;
        RECT 1181.840 241.750 1182.100 242.070 ;
        RECT 1181.380 241.410 1181.640 241.730 ;
        RECT 1181.440 234.590 1181.580 241.410 ;
        RECT 1181.380 234.270 1181.640 234.590 ;
        RECT 1181.840 186.330 1182.100 186.650 ;
        RECT 1181.900 131.230 1182.040 186.330 ;
        RECT 1181.840 130.910 1182.100 131.230 ;
        RECT 1181.840 82.970 1182.100 83.290 ;
        RECT 1181.900 17.330 1182.040 82.970 ;
        RECT 74.160 17.010 74.420 17.330 ;
        RECT 1181.840 17.010 1182.100 17.330 ;
        RECT 74.220 2.400 74.360 17.010 ;
        RECT 74.010 -4.800 74.570 2.400 ;
      LAYER via2 ;
        RECT 1181.370 1476.480 1181.650 1476.760 ;
        RECT 1182.750 1476.480 1183.030 1476.760 ;
        RECT 1182.290 1380.600 1182.570 1380.880 ;
        RECT 1181.370 1379.920 1181.650 1380.200 ;
        RECT 1179.990 1269.760 1180.270 1270.040 ;
        RECT 1181.370 1269.760 1181.650 1270.040 ;
        RECT 1182.290 814.840 1182.570 815.120 ;
        RECT 1181.370 814.160 1181.650 814.440 ;
        RECT 1181.830 670.000 1182.110 670.280 ;
        RECT 1181.370 669.320 1181.650 669.600 ;
      LAYER met3 ;
        RECT 1181.345 1476.770 1181.675 1476.785 ;
        RECT 1182.725 1476.770 1183.055 1476.785 ;
        RECT 1181.345 1476.470 1183.055 1476.770 ;
        RECT 1181.345 1476.455 1181.675 1476.470 ;
        RECT 1182.725 1476.455 1183.055 1476.470 ;
        RECT 1182.265 1380.890 1182.595 1380.905 ;
        RECT 1180.670 1380.590 1182.595 1380.890 ;
        RECT 1180.670 1380.210 1180.970 1380.590 ;
        RECT 1182.265 1380.575 1182.595 1380.590 ;
        RECT 1181.345 1380.210 1181.675 1380.225 ;
        RECT 1180.670 1379.910 1181.675 1380.210 ;
        RECT 1181.345 1379.895 1181.675 1379.910 ;
        RECT 1179.965 1270.050 1180.295 1270.065 ;
        RECT 1181.345 1270.050 1181.675 1270.065 ;
        RECT 1179.965 1269.750 1181.675 1270.050 ;
        RECT 1179.965 1269.735 1180.295 1269.750 ;
        RECT 1181.345 1269.735 1181.675 1269.750 ;
        RECT 1182.265 815.130 1182.595 815.145 ;
        RECT 1181.360 814.830 1182.595 815.130 ;
        RECT 1181.360 814.465 1181.660 814.830 ;
        RECT 1182.265 814.815 1182.595 814.830 ;
        RECT 1181.345 814.135 1181.675 814.465 ;
        RECT 1181.805 670.290 1182.135 670.305 ;
        RECT 1181.590 669.975 1182.135 670.290 ;
        RECT 1181.590 669.625 1181.890 669.975 ;
        RECT 1181.345 669.310 1181.890 669.625 ;
        RECT 1181.345 669.295 1181.675 669.310 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 493.265 14.025 493.435 14.875 ;
      LAYER mcon ;
        RECT 493.265 14.705 493.435 14.875 ;
      LAYER met1 ;
        RECT 527.690 1684.260 528.010 1684.320 ;
        RECT 1370.410 1684.260 1370.730 1684.320 ;
        RECT 527.690 1684.120 1370.730 1684.260 ;
        RECT 527.690 1684.060 528.010 1684.120 ;
        RECT 1370.410 1684.060 1370.730 1684.120 ;
        RECT 430.630 14.860 430.950 14.920 ;
        RECT 493.205 14.860 493.495 14.905 ;
        RECT 430.630 14.720 493.495 14.860 ;
        RECT 430.630 14.660 430.950 14.720 ;
        RECT 493.205 14.675 493.495 14.720 ;
        RECT 493.205 14.180 493.495 14.225 ;
        RECT 527.690 14.180 528.010 14.240 ;
        RECT 493.205 14.040 528.010 14.180 ;
        RECT 493.205 13.995 493.495 14.040 ;
        RECT 527.690 13.980 528.010 14.040 ;
      LAYER via ;
        RECT 527.720 1684.060 527.980 1684.320 ;
        RECT 1370.440 1684.060 1370.700 1684.320 ;
        RECT 430.660 14.660 430.920 14.920 ;
        RECT 527.720 13.980 527.980 14.240 ;
      LAYER met2 ;
        RECT 1370.360 1700.000 1370.640 1704.000 ;
        RECT 1370.500 1684.350 1370.640 1700.000 ;
        RECT 527.720 1684.030 527.980 1684.350 ;
        RECT 1370.440 1684.030 1370.700 1684.350 ;
        RECT 430.660 14.630 430.920 14.950 ;
        RECT 430.720 2.400 430.860 14.630 ;
        RECT 527.780 14.270 527.920 1684.030 ;
        RECT 527.720 13.950 527.980 14.270 ;
        RECT 430.510 -4.800 431.070 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1337.365 1686.825 1337.535 1687.675 ;
      LAYER mcon ;
        RECT 1337.365 1687.505 1337.535 1687.675 ;
      LAYER met1 ;
        RECT 1314.290 1687.660 1314.610 1687.720 ;
        RECT 1337.305 1687.660 1337.595 1687.705 ;
        RECT 1314.290 1687.520 1337.595 1687.660 ;
        RECT 1314.290 1687.460 1314.610 1687.520 ;
        RECT 1337.305 1687.475 1337.595 1687.520 ;
        RECT 1337.305 1686.980 1337.595 1687.025 ;
        RECT 1379.610 1686.980 1379.930 1687.040 ;
        RECT 1337.305 1686.840 1379.930 1686.980 ;
        RECT 1337.305 1686.795 1337.595 1686.840 ;
        RECT 1379.610 1686.780 1379.930 1686.840 ;
        RECT 449.030 15.880 449.350 15.940 ;
        RECT 1314.290 15.880 1314.610 15.940 ;
        RECT 449.030 15.740 1314.610 15.880 ;
        RECT 449.030 15.680 449.350 15.740 ;
        RECT 1314.290 15.680 1314.610 15.740 ;
      LAYER via ;
        RECT 1314.320 1687.460 1314.580 1687.720 ;
        RECT 1379.640 1686.780 1379.900 1687.040 ;
        RECT 449.060 15.680 449.320 15.940 ;
        RECT 1314.320 15.680 1314.580 15.940 ;
      LAYER met2 ;
        RECT 1379.560 1700.000 1379.840 1704.000 ;
        RECT 1314.320 1687.430 1314.580 1687.750 ;
        RECT 1314.380 15.970 1314.520 1687.430 ;
        RECT 1379.700 1687.070 1379.840 1700.000 ;
        RECT 1379.640 1686.750 1379.900 1687.070 ;
        RECT 449.060 15.650 449.320 15.970 ;
        RECT 1314.320 15.650 1314.580 15.970 ;
        RECT 449.120 7.890 449.260 15.650 ;
        RECT 448.660 7.750 449.260 7.890 ;
        RECT 448.660 2.400 448.800 7.750 ;
        RECT 448.450 -4.800 449.010 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 486.290 1685.960 486.610 1686.020 ;
        RECT 1388.810 1685.960 1389.130 1686.020 ;
        RECT 486.290 1685.820 1389.130 1685.960 ;
        RECT 486.290 1685.760 486.610 1685.820 ;
        RECT 1388.810 1685.760 1389.130 1685.820 ;
        RECT 486.290 15.540 486.610 15.600 ;
        RECT 483.160 15.400 486.610 15.540 ;
        RECT 466.510 15.200 466.830 15.260 ;
        RECT 483.160 15.200 483.300 15.400 ;
        RECT 486.290 15.340 486.610 15.400 ;
        RECT 466.510 15.060 483.300 15.200 ;
        RECT 466.510 15.000 466.830 15.060 ;
      LAYER via ;
        RECT 486.320 1685.760 486.580 1686.020 ;
        RECT 1388.840 1685.760 1389.100 1686.020 ;
        RECT 466.540 15.000 466.800 15.260 ;
        RECT 486.320 15.340 486.580 15.600 ;
      LAYER met2 ;
        RECT 1388.760 1700.000 1389.040 1704.000 ;
        RECT 1388.900 1686.050 1389.040 1700.000 ;
        RECT 486.320 1685.730 486.580 1686.050 ;
        RECT 1388.840 1685.730 1389.100 1686.050 ;
        RECT 486.380 15.630 486.520 1685.730 ;
        RECT 486.320 15.310 486.580 15.630 ;
        RECT 466.540 14.970 466.800 15.290 ;
        RECT 466.600 2.400 466.740 14.970 ;
        RECT 466.390 -4.800 466.950 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1321.190 1687.320 1321.510 1687.380 ;
        RECT 1398.010 1687.320 1398.330 1687.380 ;
        RECT 1321.190 1687.180 1398.330 1687.320 ;
        RECT 1321.190 1687.120 1321.510 1687.180 ;
        RECT 1398.010 1687.120 1398.330 1687.180 ;
        RECT 1321.190 15.540 1321.510 15.600 ;
        RECT 559.060 15.400 1321.510 15.540 ;
        RECT 484.450 15.200 484.770 15.260 ;
        RECT 559.060 15.200 559.200 15.400 ;
        RECT 1321.190 15.340 1321.510 15.400 ;
        RECT 484.450 15.060 493.880 15.200 ;
        RECT 484.450 15.000 484.770 15.060 ;
        RECT 493.740 14.860 493.880 15.060 ;
        RECT 496.960 15.060 559.200 15.200 ;
        RECT 496.960 14.860 497.100 15.060 ;
        RECT 493.740 14.720 497.100 14.860 ;
      LAYER via ;
        RECT 1321.220 1687.120 1321.480 1687.380 ;
        RECT 1398.040 1687.120 1398.300 1687.380 ;
        RECT 484.480 15.000 484.740 15.260 ;
        RECT 1321.220 15.340 1321.480 15.600 ;
      LAYER met2 ;
        RECT 1397.960 1700.000 1398.240 1704.000 ;
        RECT 1398.100 1687.410 1398.240 1700.000 ;
        RECT 1321.220 1687.090 1321.480 1687.410 ;
        RECT 1398.040 1687.090 1398.300 1687.410 ;
        RECT 1321.280 15.630 1321.420 1687.090 ;
        RECT 1321.220 15.310 1321.480 15.630 ;
        RECT 484.480 14.970 484.740 15.290 ;
        RECT 484.540 2.400 484.680 14.970 ;
        RECT 484.330 -4.800 484.890 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1321.650 1688.340 1321.970 1688.400 ;
        RECT 1407.210 1688.340 1407.530 1688.400 ;
        RECT 1321.650 1688.200 1407.530 1688.340 ;
        RECT 1321.650 1688.140 1321.970 1688.200 ;
        RECT 1407.210 1688.140 1407.530 1688.200 ;
        RECT 1321.650 15.200 1321.970 15.260 ;
        RECT 559.520 15.060 1321.970 15.200 ;
        RECT 502.390 14.520 502.710 14.580 ;
        RECT 559.520 14.520 559.660 15.060 ;
        RECT 1321.650 15.000 1321.970 15.060 ;
        RECT 502.390 14.380 559.660 14.520 ;
        RECT 502.390 14.320 502.710 14.380 ;
      LAYER via ;
        RECT 1321.680 1688.140 1321.940 1688.400 ;
        RECT 1407.240 1688.140 1407.500 1688.400 ;
        RECT 502.420 14.320 502.680 14.580 ;
        RECT 1321.680 15.000 1321.940 15.260 ;
      LAYER met2 ;
        RECT 1407.160 1700.000 1407.440 1704.000 ;
        RECT 1407.300 1688.430 1407.440 1700.000 ;
        RECT 1321.680 1688.110 1321.940 1688.430 ;
        RECT 1407.240 1688.110 1407.500 1688.430 ;
        RECT 1321.740 15.290 1321.880 1688.110 ;
        RECT 1321.680 14.970 1321.940 15.290 ;
        RECT 502.420 14.290 502.680 14.610 ;
        RECT 502.480 2.400 502.620 14.290 ;
        RECT 502.270 -4.800 502.830 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 524.010 1685.620 524.330 1685.680 ;
        RECT 1415.950 1685.620 1416.270 1685.680 ;
        RECT 524.010 1685.480 1416.270 1685.620 ;
        RECT 524.010 1685.420 524.330 1685.480 ;
        RECT 1415.950 1685.420 1416.270 1685.480 ;
        RECT 519.870 15.540 520.190 15.600 ;
        RECT 524.010 15.540 524.330 15.600 ;
        RECT 519.870 15.400 524.330 15.540 ;
        RECT 519.870 15.340 520.190 15.400 ;
        RECT 524.010 15.340 524.330 15.400 ;
      LAYER via ;
        RECT 524.040 1685.420 524.300 1685.680 ;
        RECT 1415.980 1685.420 1416.240 1685.680 ;
        RECT 519.900 15.340 520.160 15.600 ;
        RECT 524.040 15.340 524.300 15.600 ;
      LAYER met2 ;
        RECT 1415.900 1700.000 1416.180 1704.000 ;
        RECT 1416.040 1685.710 1416.180 1700.000 ;
        RECT 524.040 1685.390 524.300 1685.710 ;
        RECT 1415.980 1685.390 1416.240 1685.710 ;
        RECT 524.100 15.630 524.240 1685.390 ;
        RECT 519.900 15.310 520.160 15.630 ;
        RECT 524.040 15.310 524.300 15.630 ;
        RECT 519.960 2.400 520.100 15.310 ;
        RECT 519.750 -4.800 520.310 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1337.825 1642.285 1337.995 1687.675 ;
        RECT 1335.525 1538.925 1335.695 1545.895 ;
        RECT 1335.065 1400.885 1335.235 1490.475 ;
        RECT 1335.525 1304.325 1335.695 1352.435 ;
        RECT 1335.985 866.405 1336.155 910.775 ;
        RECT 1335.985 614.125 1336.155 662.235 ;
        RECT 1335.065 227.885 1335.235 275.655 ;
        RECT 1335.525 144.925 1335.695 210.375 ;
      LAYER mcon ;
        RECT 1337.825 1687.505 1337.995 1687.675 ;
        RECT 1335.525 1545.725 1335.695 1545.895 ;
        RECT 1335.065 1490.305 1335.235 1490.475 ;
        RECT 1335.525 1352.265 1335.695 1352.435 ;
        RECT 1335.985 910.605 1336.155 910.775 ;
        RECT 1335.985 662.065 1336.155 662.235 ;
        RECT 1335.065 275.485 1335.235 275.655 ;
        RECT 1335.525 210.205 1335.695 210.375 ;
      LAYER met1 ;
        RECT 1337.765 1687.660 1338.055 1687.705 ;
        RECT 1425.150 1687.660 1425.470 1687.720 ;
        RECT 1337.765 1687.520 1425.470 1687.660 ;
        RECT 1337.765 1687.475 1338.055 1687.520 ;
        RECT 1425.150 1687.460 1425.470 1687.520 ;
        RECT 1335.450 1642.440 1335.770 1642.500 ;
        RECT 1337.765 1642.440 1338.055 1642.485 ;
        RECT 1335.450 1642.300 1338.055 1642.440 ;
        RECT 1335.450 1642.240 1335.770 1642.300 ;
        RECT 1337.765 1642.255 1338.055 1642.300 ;
        RECT 1335.450 1545.880 1335.770 1545.940 ;
        RECT 1335.255 1545.740 1335.770 1545.880 ;
        RECT 1335.450 1545.680 1335.770 1545.740 ;
        RECT 1335.450 1539.080 1335.770 1539.140 ;
        RECT 1335.255 1538.940 1335.770 1539.080 ;
        RECT 1335.450 1538.880 1335.770 1538.940 ;
        RECT 1335.005 1490.460 1335.295 1490.505 ;
        RECT 1335.450 1490.460 1335.770 1490.520 ;
        RECT 1335.005 1490.320 1335.770 1490.460 ;
        RECT 1335.005 1490.275 1335.295 1490.320 ;
        RECT 1335.450 1490.260 1335.770 1490.320 ;
        RECT 1334.990 1401.040 1335.310 1401.100 ;
        RECT 1334.795 1400.900 1335.310 1401.040 ;
        RECT 1334.990 1400.840 1335.310 1400.900 ;
        RECT 1335.450 1352.420 1335.770 1352.480 ;
        RECT 1335.255 1352.280 1335.770 1352.420 ;
        RECT 1335.450 1352.220 1335.770 1352.280 ;
        RECT 1335.450 1304.480 1335.770 1304.540 ;
        RECT 1335.255 1304.340 1335.770 1304.480 ;
        RECT 1335.450 1304.280 1335.770 1304.340 ;
        RECT 1335.450 1268.580 1335.770 1268.840 ;
        RECT 1335.540 1268.440 1335.680 1268.580 ;
        RECT 1335.910 1268.440 1336.230 1268.500 ;
        RECT 1335.540 1268.300 1336.230 1268.440 ;
        RECT 1335.910 1268.240 1336.230 1268.300 ;
        RECT 1334.070 1207.580 1334.390 1207.640 ;
        RECT 1334.530 1207.580 1334.850 1207.640 ;
        RECT 1334.070 1207.440 1334.850 1207.580 ;
        RECT 1334.070 1207.380 1334.390 1207.440 ;
        RECT 1334.530 1207.380 1334.850 1207.440 ;
        RECT 1333.610 1104.220 1333.930 1104.280 ;
        RECT 1334.530 1104.220 1334.850 1104.280 ;
        RECT 1333.610 1104.080 1334.850 1104.220 ;
        RECT 1333.610 1104.020 1333.930 1104.080 ;
        RECT 1334.530 1104.020 1334.850 1104.080 ;
        RECT 1334.990 966.180 1335.310 966.240 ;
        RECT 1335.450 966.180 1335.770 966.240 ;
        RECT 1334.990 966.040 1335.770 966.180 ;
        RECT 1334.990 965.980 1335.310 966.040 ;
        RECT 1335.450 965.980 1335.770 966.040 ;
        RECT 1335.910 910.760 1336.230 910.820 ;
        RECT 1335.715 910.620 1336.230 910.760 ;
        RECT 1335.910 910.560 1336.230 910.620 ;
        RECT 1335.910 866.560 1336.230 866.620 ;
        RECT 1335.715 866.420 1336.230 866.560 ;
        RECT 1335.910 866.360 1336.230 866.420 ;
        RECT 1334.530 821.000 1334.850 821.060 ;
        RECT 1334.990 821.000 1335.310 821.060 ;
        RECT 1334.530 820.860 1335.310 821.000 ;
        RECT 1334.530 820.800 1334.850 820.860 ;
        RECT 1334.990 820.800 1335.310 820.860 ;
        RECT 1335.925 662.220 1336.215 662.265 ;
        RECT 1336.370 662.220 1336.690 662.280 ;
        RECT 1335.925 662.080 1336.690 662.220 ;
        RECT 1335.925 662.035 1336.215 662.080 ;
        RECT 1336.370 662.020 1336.690 662.080 ;
        RECT 1335.910 614.280 1336.230 614.340 ;
        RECT 1335.715 614.140 1336.230 614.280 ;
        RECT 1335.910 614.080 1336.230 614.140 ;
        RECT 1334.530 589.120 1334.850 589.180 ;
        RECT 1335.910 589.120 1336.230 589.180 ;
        RECT 1334.530 588.980 1336.230 589.120 ;
        RECT 1334.530 588.920 1334.850 588.980 ;
        RECT 1335.910 588.920 1336.230 588.980 ;
        RECT 1334.530 476.240 1334.850 476.300 ;
        RECT 1335.450 476.240 1335.770 476.300 ;
        RECT 1334.530 476.100 1335.770 476.240 ;
        RECT 1334.530 476.040 1334.850 476.100 ;
        RECT 1335.450 476.040 1335.770 476.100 ;
        RECT 1335.450 435.100 1335.770 435.160 ;
        RECT 1335.080 434.960 1335.770 435.100 ;
        RECT 1335.080 434.820 1335.220 434.960 ;
        RECT 1335.450 434.900 1335.770 434.960 ;
        RECT 1334.990 434.560 1335.310 434.820 ;
        RECT 1334.990 373.220 1335.310 373.280 ;
        RECT 1334.990 373.080 1336.140 373.220 ;
        RECT 1334.990 373.020 1335.310 373.080 ;
        RECT 1334.070 372.540 1334.390 372.600 ;
        RECT 1336.000 372.540 1336.140 373.080 ;
        RECT 1334.070 372.400 1336.140 372.540 ;
        RECT 1334.070 372.340 1334.390 372.400 ;
        RECT 1334.070 276.320 1334.390 276.380 ;
        RECT 1334.990 276.320 1335.310 276.380 ;
        RECT 1334.070 276.180 1335.310 276.320 ;
        RECT 1334.070 276.120 1334.390 276.180 ;
        RECT 1334.990 276.120 1335.310 276.180 ;
        RECT 1334.990 275.640 1335.310 275.700 ;
        RECT 1334.795 275.500 1335.310 275.640 ;
        RECT 1334.990 275.440 1335.310 275.500 ;
        RECT 1335.005 228.040 1335.295 228.085 ;
        RECT 1335.450 228.040 1335.770 228.100 ;
        RECT 1335.005 227.900 1335.770 228.040 ;
        RECT 1335.005 227.855 1335.295 227.900 ;
        RECT 1335.450 227.840 1335.770 227.900 ;
        RECT 1335.450 210.360 1335.770 210.420 ;
        RECT 1335.255 210.220 1335.770 210.360 ;
        RECT 1335.450 210.160 1335.770 210.220 ;
        RECT 1335.450 145.080 1335.770 145.140 ;
        RECT 1335.255 144.940 1335.770 145.080 ;
        RECT 1335.450 144.880 1335.770 144.940 ;
        RECT 1334.530 14.860 1334.850 14.920 ;
        RECT 607.820 14.720 1334.850 14.860 ;
        RECT 537.810 14.180 538.130 14.240 ;
        RECT 607.820 14.180 607.960 14.720 ;
        RECT 1334.530 14.660 1334.850 14.720 ;
        RECT 537.810 14.040 607.960 14.180 ;
        RECT 537.810 13.980 538.130 14.040 ;
      LAYER via ;
        RECT 1425.180 1687.460 1425.440 1687.720 ;
        RECT 1335.480 1642.240 1335.740 1642.500 ;
        RECT 1335.480 1545.680 1335.740 1545.940 ;
        RECT 1335.480 1538.880 1335.740 1539.140 ;
        RECT 1335.480 1490.260 1335.740 1490.520 ;
        RECT 1335.020 1400.840 1335.280 1401.100 ;
        RECT 1335.480 1352.220 1335.740 1352.480 ;
        RECT 1335.480 1304.280 1335.740 1304.540 ;
        RECT 1335.480 1268.580 1335.740 1268.840 ;
        RECT 1335.940 1268.240 1336.200 1268.500 ;
        RECT 1334.100 1207.380 1334.360 1207.640 ;
        RECT 1334.560 1207.380 1334.820 1207.640 ;
        RECT 1333.640 1104.020 1333.900 1104.280 ;
        RECT 1334.560 1104.020 1334.820 1104.280 ;
        RECT 1335.020 965.980 1335.280 966.240 ;
        RECT 1335.480 965.980 1335.740 966.240 ;
        RECT 1335.940 910.560 1336.200 910.820 ;
        RECT 1335.940 866.360 1336.200 866.620 ;
        RECT 1334.560 820.800 1334.820 821.060 ;
        RECT 1335.020 820.800 1335.280 821.060 ;
        RECT 1336.400 662.020 1336.660 662.280 ;
        RECT 1335.940 614.080 1336.200 614.340 ;
        RECT 1334.560 588.920 1334.820 589.180 ;
        RECT 1335.940 588.920 1336.200 589.180 ;
        RECT 1334.560 476.040 1334.820 476.300 ;
        RECT 1335.480 476.040 1335.740 476.300 ;
        RECT 1335.480 434.900 1335.740 435.160 ;
        RECT 1335.020 434.560 1335.280 434.820 ;
        RECT 1335.020 373.020 1335.280 373.280 ;
        RECT 1334.100 372.340 1334.360 372.600 ;
        RECT 1334.100 276.120 1334.360 276.380 ;
        RECT 1335.020 276.120 1335.280 276.380 ;
        RECT 1335.020 275.440 1335.280 275.700 ;
        RECT 1335.480 227.840 1335.740 228.100 ;
        RECT 1335.480 210.160 1335.740 210.420 ;
        RECT 1335.480 144.880 1335.740 145.140 ;
        RECT 537.840 13.980 538.100 14.240 ;
        RECT 1334.560 14.660 1334.820 14.920 ;
      LAYER met2 ;
        RECT 1425.100 1700.000 1425.380 1704.000 ;
        RECT 1425.240 1687.750 1425.380 1700.000 ;
        RECT 1425.180 1687.430 1425.440 1687.750 ;
        RECT 1335.480 1642.210 1335.740 1642.530 ;
        RECT 1335.540 1545.970 1335.680 1642.210 ;
        RECT 1335.480 1545.650 1335.740 1545.970 ;
        RECT 1335.480 1538.850 1335.740 1539.170 ;
        RECT 1335.540 1490.550 1335.680 1538.850 ;
        RECT 1335.480 1490.230 1335.740 1490.550 ;
        RECT 1335.020 1400.810 1335.280 1401.130 ;
        RECT 1335.080 1376.050 1335.220 1400.810 ;
        RECT 1335.080 1375.910 1335.680 1376.050 ;
        RECT 1335.540 1352.510 1335.680 1375.910 ;
        RECT 1335.480 1352.190 1335.740 1352.510 ;
        RECT 1335.480 1304.250 1335.740 1304.570 ;
        RECT 1335.540 1268.870 1335.680 1304.250 ;
        RECT 1335.480 1268.550 1335.740 1268.870 ;
        RECT 1335.940 1268.210 1336.200 1268.530 ;
        RECT 1336.000 1256.200 1336.140 1268.210 ;
        RECT 1335.540 1256.060 1336.140 1256.200 ;
        RECT 1335.540 1255.690 1335.680 1256.060 ;
        RECT 1334.620 1255.550 1335.680 1255.690 ;
        RECT 1334.620 1207.670 1334.760 1255.550 ;
        RECT 1334.100 1207.350 1334.360 1207.670 ;
        RECT 1334.560 1207.350 1334.820 1207.670 ;
        RECT 1334.160 1200.725 1334.300 1207.350 ;
        RECT 1334.090 1200.355 1334.370 1200.725 ;
        RECT 1335.470 1200.355 1335.750 1200.725 ;
        RECT 1335.540 1152.445 1335.680 1200.355 ;
        RECT 1333.630 1152.075 1333.910 1152.445 ;
        RECT 1335.470 1152.075 1335.750 1152.445 ;
        RECT 1333.700 1104.310 1333.840 1152.075 ;
        RECT 1333.640 1103.990 1333.900 1104.310 ;
        RECT 1334.560 1103.990 1334.820 1104.310 ;
        RECT 1334.620 1055.770 1334.760 1103.990 ;
        RECT 1334.620 1055.630 1335.220 1055.770 ;
        RECT 1335.080 966.270 1335.220 1055.630 ;
        RECT 1335.020 965.950 1335.280 966.270 ;
        RECT 1335.480 965.950 1335.740 966.270 ;
        RECT 1335.540 942.210 1335.680 965.950 ;
        RECT 1335.080 942.070 1335.680 942.210 ;
        RECT 1335.080 917.845 1335.220 942.070 ;
        RECT 1335.010 917.475 1335.290 917.845 ;
        RECT 1335.930 917.475 1336.210 917.845 ;
        RECT 1336.000 910.850 1336.140 917.475 ;
        RECT 1335.940 910.530 1336.200 910.850 ;
        RECT 1335.940 866.330 1336.200 866.650 ;
        RECT 1336.000 821.285 1336.140 866.330 ;
        RECT 1334.560 820.770 1334.820 821.090 ;
        RECT 1335.010 820.915 1335.290 821.285 ;
        RECT 1335.930 820.915 1336.210 821.285 ;
        RECT 1335.020 820.770 1335.280 820.915 ;
        RECT 1334.620 773.005 1334.760 820.770 ;
        RECT 1334.550 772.635 1334.830 773.005 ;
        RECT 1335.470 772.635 1335.750 773.005 ;
        RECT 1335.540 665.450 1335.680 772.635 ;
        RECT 1335.540 665.310 1336.600 665.450 ;
        RECT 1336.460 662.310 1336.600 665.310 ;
        RECT 1336.400 661.990 1336.660 662.310 ;
        RECT 1335.940 614.050 1336.200 614.370 ;
        RECT 1336.000 589.210 1336.140 614.050 ;
        RECT 1334.560 588.890 1334.820 589.210 ;
        RECT 1335.940 588.890 1336.200 589.210 ;
        RECT 1334.620 476.330 1334.760 588.890 ;
        RECT 1334.560 476.010 1334.820 476.330 ;
        RECT 1335.480 476.010 1335.740 476.330 ;
        RECT 1335.540 435.190 1335.680 476.010 ;
        RECT 1335.480 434.870 1335.740 435.190 ;
        RECT 1335.020 434.530 1335.280 434.850 ;
        RECT 1335.080 373.310 1335.220 434.530 ;
        RECT 1335.020 372.990 1335.280 373.310 ;
        RECT 1334.100 372.310 1334.360 372.630 ;
        RECT 1334.160 276.410 1334.300 372.310 ;
        RECT 1334.100 276.090 1334.360 276.410 ;
        RECT 1335.020 276.090 1335.280 276.410 ;
        RECT 1335.080 275.730 1335.220 276.090 ;
        RECT 1335.020 275.410 1335.280 275.730 ;
        RECT 1335.480 227.810 1335.740 228.130 ;
        RECT 1335.540 210.450 1335.680 227.810 ;
        RECT 1335.480 210.130 1335.740 210.450 ;
        RECT 1335.480 144.850 1335.740 145.170 ;
        RECT 1335.540 48.010 1335.680 144.850 ;
        RECT 1334.620 47.870 1335.680 48.010 ;
        RECT 1334.620 14.950 1334.760 47.870 ;
        RECT 1334.560 14.630 1334.820 14.950 ;
        RECT 537.840 13.950 538.100 14.270 ;
        RECT 537.900 2.400 538.040 13.950 ;
        RECT 537.690 -4.800 538.250 2.400 ;
      LAYER via2 ;
        RECT 1334.090 1200.400 1334.370 1200.680 ;
        RECT 1335.470 1200.400 1335.750 1200.680 ;
        RECT 1333.630 1152.120 1333.910 1152.400 ;
        RECT 1335.470 1152.120 1335.750 1152.400 ;
        RECT 1335.010 917.520 1335.290 917.800 ;
        RECT 1335.930 917.520 1336.210 917.800 ;
        RECT 1335.010 820.960 1335.290 821.240 ;
        RECT 1335.930 820.960 1336.210 821.240 ;
        RECT 1334.550 772.680 1334.830 772.960 ;
        RECT 1335.470 772.680 1335.750 772.960 ;
      LAYER met3 ;
        RECT 1334.065 1200.690 1334.395 1200.705 ;
        RECT 1335.445 1200.690 1335.775 1200.705 ;
        RECT 1334.065 1200.390 1335.775 1200.690 ;
        RECT 1334.065 1200.375 1334.395 1200.390 ;
        RECT 1335.445 1200.375 1335.775 1200.390 ;
        RECT 1333.605 1152.410 1333.935 1152.425 ;
        RECT 1335.445 1152.410 1335.775 1152.425 ;
        RECT 1333.605 1152.110 1335.775 1152.410 ;
        RECT 1333.605 1152.095 1333.935 1152.110 ;
        RECT 1335.445 1152.095 1335.775 1152.110 ;
        RECT 1334.985 917.810 1335.315 917.825 ;
        RECT 1335.905 917.810 1336.235 917.825 ;
        RECT 1334.985 917.510 1336.235 917.810 ;
        RECT 1334.985 917.495 1335.315 917.510 ;
        RECT 1335.905 917.495 1336.235 917.510 ;
        RECT 1334.985 821.250 1335.315 821.265 ;
        RECT 1335.905 821.250 1336.235 821.265 ;
        RECT 1334.985 820.950 1336.235 821.250 ;
        RECT 1334.985 820.935 1335.315 820.950 ;
        RECT 1335.905 820.935 1336.235 820.950 ;
        RECT 1334.525 772.970 1334.855 772.985 ;
        RECT 1335.445 772.970 1335.775 772.985 ;
        RECT 1334.525 772.670 1335.775 772.970 ;
        RECT 1334.525 772.655 1334.855 772.670 ;
        RECT 1335.445 772.655 1335.775 772.670 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 558.510 1685.280 558.830 1685.340 ;
        RECT 1434.350 1685.280 1434.670 1685.340 ;
        RECT 558.510 1685.140 1434.670 1685.280 ;
        RECT 558.510 1685.080 558.830 1685.140 ;
        RECT 1434.350 1685.080 1434.670 1685.140 ;
        RECT 555.750 15.540 556.070 15.600 ;
        RECT 558.510 15.540 558.830 15.600 ;
        RECT 555.750 15.400 558.830 15.540 ;
        RECT 555.750 15.340 556.070 15.400 ;
        RECT 558.510 15.340 558.830 15.400 ;
      LAYER via ;
        RECT 558.540 1685.080 558.800 1685.340 ;
        RECT 1434.380 1685.080 1434.640 1685.340 ;
        RECT 555.780 15.340 556.040 15.600 ;
        RECT 558.540 15.340 558.800 15.600 ;
      LAYER met2 ;
        RECT 1434.300 1700.000 1434.580 1704.000 ;
        RECT 1434.440 1685.370 1434.580 1700.000 ;
        RECT 558.540 1685.050 558.800 1685.370 ;
        RECT 1434.380 1685.050 1434.640 1685.370 ;
        RECT 558.600 15.630 558.740 1685.050 ;
        RECT 555.780 15.310 556.040 15.630 ;
        RECT 558.540 15.310 558.800 15.630 ;
        RECT 555.840 2.400 555.980 15.310 ;
        RECT 555.630 -4.800 556.190 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 607.345 14.365 608.435 14.535 ;
      LAYER mcon ;
        RECT 608.265 14.365 608.435 14.535 ;
      LAYER met1 ;
        RECT 1341.890 1689.360 1342.210 1689.420 ;
        RECT 1443.550 1689.360 1443.870 1689.420 ;
        RECT 1341.890 1689.220 1443.870 1689.360 ;
        RECT 1341.890 1689.160 1342.210 1689.220 ;
        RECT 1443.550 1689.160 1443.870 1689.220 ;
        RECT 573.690 14.520 574.010 14.580 ;
        RECT 607.285 14.520 607.575 14.565 ;
        RECT 573.690 14.380 607.575 14.520 ;
        RECT 573.690 14.320 574.010 14.380 ;
        RECT 607.285 14.335 607.575 14.380 ;
        RECT 608.205 14.520 608.495 14.565 ;
        RECT 1341.890 14.520 1342.210 14.580 ;
        RECT 608.205 14.380 1342.210 14.520 ;
        RECT 608.205 14.335 608.495 14.380 ;
        RECT 1341.890 14.320 1342.210 14.380 ;
      LAYER via ;
        RECT 1341.920 1689.160 1342.180 1689.420 ;
        RECT 1443.580 1689.160 1443.840 1689.420 ;
        RECT 573.720 14.320 573.980 14.580 ;
        RECT 1341.920 14.320 1342.180 14.580 ;
      LAYER met2 ;
        RECT 1443.500 1700.000 1443.780 1704.000 ;
        RECT 1443.640 1689.450 1443.780 1700.000 ;
        RECT 1341.920 1689.130 1342.180 1689.450 ;
        RECT 1443.580 1689.130 1443.840 1689.450 ;
        RECT 1341.980 14.610 1342.120 1689.130 ;
        RECT 573.720 14.290 573.980 14.610 ;
        RECT 1341.920 14.290 1342.180 14.610 ;
        RECT 573.780 2.400 573.920 14.290 ;
        RECT 573.570 -4.800 574.130 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 593.010 1684.940 593.330 1685.000 ;
        RECT 1452.750 1684.940 1453.070 1685.000 ;
        RECT 593.010 1684.800 1453.070 1684.940 ;
        RECT 593.010 1684.740 593.330 1684.800 ;
        RECT 1452.750 1684.740 1453.070 1684.800 ;
      LAYER via ;
        RECT 593.040 1684.740 593.300 1685.000 ;
        RECT 1452.780 1684.740 1453.040 1685.000 ;
      LAYER met2 ;
        RECT 1452.700 1700.000 1452.980 1704.000 ;
        RECT 1452.840 1685.030 1452.980 1700.000 ;
        RECT 593.040 1684.710 593.300 1685.030 ;
        RECT 1452.780 1684.710 1453.040 1685.030 ;
        RECT 593.100 16.730 593.240 1684.710 ;
        RECT 591.260 16.590 593.240 16.730 ;
        RECT 591.260 2.400 591.400 16.590 ;
        RECT 591.050 -4.800 591.610 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 120.590 1687.320 120.910 1687.380 ;
        RECT 120.590 1687.180 1186.180 1687.320 ;
        RECT 120.590 1687.120 120.910 1687.180 ;
        RECT 1186.040 1686.980 1186.180 1687.180 ;
        RECT 1198.830 1686.980 1199.150 1687.040 ;
        RECT 1186.040 1686.840 1199.150 1686.980 ;
        RECT 1198.830 1686.780 1199.150 1686.840 ;
        RECT 97.590 17.920 97.910 17.980 ;
        RECT 120.590 17.920 120.910 17.980 ;
        RECT 97.590 17.780 120.910 17.920 ;
        RECT 97.590 17.720 97.910 17.780 ;
        RECT 120.590 17.720 120.910 17.780 ;
      LAYER via ;
        RECT 120.620 1687.120 120.880 1687.380 ;
        RECT 1198.860 1686.780 1199.120 1687.040 ;
        RECT 97.620 17.720 97.880 17.980 ;
        RECT 120.620 17.720 120.880 17.980 ;
      LAYER met2 ;
        RECT 1198.780 1700.000 1199.060 1704.000 ;
        RECT 120.620 1687.090 120.880 1687.410 ;
        RECT 120.680 18.010 120.820 1687.090 ;
        RECT 1198.920 1687.070 1199.060 1700.000 ;
        RECT 1198.860 1686.750 1199.120 1687.070 ;
        RECT 97.620 17.690 97.880 18.010 ;
        RECT 120.620 17.690 120.880 18.010 ;
        RECT 97.680 2.400 97.820 17.690 ;
        RECT 97.470 -4.800 98.030 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1348.790 1689.020 1349.110 1689.080 ;
        RECT 1461.950 1689.020 1462.270 1689.080 ;
        RECT 1348.790 1688.880 1462.270 1689.020 ;
        RECT 1348.790 1688.820 1349.110 1688.880 ;
        RECT 1461.950 1688.820 1462.270 1688.880 ;
        RECT 609.110 14.180 609.430 14.240 ;
        RECT 1348.790 14.180 1349.110 14.240 ;
        RECT 609.110 14.040 1349.110 14.180 ;
        RECT 609.110 13.980 609.430 14.040 ;
        RECT 1348.790 13.980 1349.110 14.040 ;
      LAYER via ;
        RECT 1348.820 1688.820 1349.080 1689.080 ;
        RECT 1461.980 1688.820 1462.240 1689.080 ;
        RECT 609.140 13.980 609.400 14.240 ;
        RECT 1348.820 13.980 1349.080 14.240 ;
      LAYER met2 ;
        RECT 1461.900 1700.000 1462.180 1704.000 ;
        RECT 1462.040 1689.110 1462.180 1700.000 ;
        RECT 1348.820 1688.790 1349.080 1689.110 ;
        RECT 1461.980 1688.790 1462.240 1689.110 ;
        RECT 1348.880 14.270 1349.020 1688.790 ;
        RECT 609.140 13.950 609.400 14.270 ;
        RECT 1348.820 13.950 1349.080 14.270 ;
        RECT 609.200 2.400 609.340 13.950 ;
        RECT 608.990 -4.800 609.550 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 627.510 1684.600 627.830 1684.660 ;
        RECT 1471.150 1684.600 1471.470 1684.660 ;
        RECT 627.510 1684.460 1471.470 1684.600 ;
        RECT 627.510 1684.400 627.830 1684.460 ;
        RECT 1471.150 1684.400 1471.470 1684.460 ;
      LAYER via ;
        RECT 627.540 1684.400 627.800 1684.660 ;
        RECT 1471.180 1684.400 1471.440 1684.660 ;
      LAYER met2 ;
        RECT 1471.100 1700.000 1471.380 1704.000 ;
        RECT 1471.240 1684.690 1471.380 1700.000 ;
        RECT 627.540 1684.370 627.800 1684.690 ;
        RECT 1471.180 1684.370 1471.440 1684.690 ;
        RECT 627.600 17.410 627.740 1684.370 ;
        RECT 627.140 17.270 627.740 17.410 ;
        RECT 627.140 2.400 627.280 17.270 ;
        RECT 626.930 -4.800 627.490 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1207.570 1678.140 1207.890 1678.200 ;
        RECT 1209.870 1678.140 1210.190 1678.200 ;
        RECT 1207.570 1678.000 1210.190 1678.140 ;
        RECT 1207.570 1677.940 1207.890 1678.000 ;
        RECT 1209.870 1677.940 1210.190 1678.000 ;
        RECT 121.510 17.920 121.830 17.980 ;
        RECT 1207.570 17.920 1207.890 17.980 ;
        RECT 121.510 17.780 1207.890 17.920 ;
        RECT 121.510 17.720 121.830 17.780 ;
        RECT 1207.570 17.720 1207.890 17.780 ;
      LAYER via ;
        RECT 1207.600 1677.940 1207.860 1678.200 ;
        RECT 1209.900 1677.940 1210.160 1678.200 ;
        RECT 121.540 17.720 121.800 17.980 ;
        RECT 1207.600 17.720 1207.860 17.980 ;
      LAYER met2 ;
        RECT 1211.200 1700.410 1211.480 1704.000 ;
        RECT 1209.960 1700.270 1211.480 1700.410 ;
        RECT 1209.960 1678.230 1210.100 1700.270 ;
        RECT 1211.200 1700.000 1211.480 1700.270 ;
        RECT 1207.600 1677.910 1207.860 1678.230 ;
        RECT 1209.900 1677.910 1210.160 1678.230 ;
        RECT 1207.660 18.010 1207.800 1677.910 ;
        RECT 121.540 17.690 121.800 18.010 ;
        RECT 1207.600 17.690 1207.860 18.010 ;
        RECT 121.600 2.400 121.740 17.690 ;
        RECT 121.390 -4.800 121.950 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1197.065 1687.505 1197.235 1688.355 ;
      LAYER mcon ;
        RECT 1197.065 1688.185 1197.235 1688.355 ;
      LAYER met1 ;
        RECT 161.990 1688.340 162.310 1688.400 ;
        RECT 1197.005 1688.340 1197.295 1688.385 ;
        RECT 161.990 1688.200 1197.295 1688.340 ;
        RECT 161.990 1688.140 162.310 1688.200 ;
        RECT 1197.005 1688.155 1197.295 1688.200 ;
        RECT 1197.005 1687.660 1197.295 1687.705 ;
        RECT 1223.210 1687.660 1223.530 1687.720 ;
        RECT 1197.005 1687.520 1223.530 1687.660 ;
        RECT 1197.005 1687.475 1197.295 1687.520 ;
        RECT 1223.210 1687.460 1223.530 1687.520 ;
        RECT 145.430 15.880 145.750 15.940 ;
        RECT 161.990 15.880 162.310 15.940 ;
        RECT 145.430 15.740 162.310 15.880 ;
        RECT 145.430 15.680 145.750 15.740 ;
        RECT 161.990 15.680 162.310 15.740 ;
      LAYER via ;
        RECT 162.020 1688.140 162.280 1688.400 ;
        RECT 1223.240 1687.460 1223.500 1687.720 ;
        RECT 145.460 15.680 145.720 15.940 ;
        RECT 162.020 15.680 162.280 15.940 ;
      LAYER met2 ;
        RECT 1223.160 1700.000 1223.440 1704.000 ;
        RECT 162.020 1688.110 162.280 1688.430 ;
        RECT 162.080 15.970 162.220 1688.110 ;
        RECT 1223.300 1687.750 1223.440 1700.000 ;
        RECT 1223.240 1687.430 1223.500 1687.750 ;
        RECT 145.460 15.650 145.720 15.970 ;
        RECT 162.020 15.650 162.280 15.970 ;
        RECT 145.520 2.400 145.660 15.650 ;
        RECT 145.310 -4.800 145.870 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1228.270 1678.140 1228.590 1678.200 ;
        RECT 1231.030 1678.140 1231.350 1678.200 ;
        RECT 1228.270 1678.000 1231.350 1678.140 ;
        RECT 1228.270 1677.940 1228.590 1678.000 ;
        RECT 1231.030 1677.940 1231.350 1678.000 ;
        RECT 163.370 18.600 163.690 18.660 ;
        RECT 1228.270 18.600 1228.590 18.660 ;
        RECT 163.370 18.460 1228.590 18.600 ;
        RECT 163.370 18.400 163.690 18.460 ;
        RECT 1228.270 18.400 1228.590 18.460 ;
      LAYER via ;
        RECT 1228.300 1677.940 1228.560 1678.200 ;
        RECT 1231.060 1677.940 1231.320 1678.200 ;
        RECT 163.400 18.400 163.660 18.660 ;
        RECT 1228.300 18.400 1228.560 18.660 ;
      LAYER met2 ;
        RECT 1232.360 1700.410 1232.640 1704.000 ;
        RECT 1231.120 1700.270 1232.640 1700.410 ;
        RECT 1231.120 1678.230 1231.260 1700.270 ;
        RECT 1232.360 1700.000 1232.640 1700.270 ;
        RECT 1228.300 1677.910 1228.560 1678.230 ;
        RECT 1231.060 1677.910 1231.320 1678.230 ;
        RECT 1228.360 18.690 1228.500 1677.910 ;
        RECT 163.400 18.370 163.660 18.690 ;
        RECT 1228.300 18.370 1228.560 18.690 ;
        RECT 163.460 2.400 163.600 18.370 ;
        RECT 163.250 -4.800 163.810 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1173.145 1688.525 1175.155 1688.695 ;
        RECT 1174.985 1687.505 1175.155 1688.525 ;
      LAYER met1 ;
        RECT 196.490 1688.680 196.810 1688.740 ;
        RECT 1173.085 1688.680 1173.375 1688.725 ;
        RECT 196.490 1688.540 1173.375 1688.680 ;
        RECT 196.490 1688.480 196.810 1688.540 ;
        RECT 1173.085 1688.495 1173.375 1688.540 ;
        RECT 1241.610 1688.000 1241.930 1688.060 ;
        RECT 1187.880 1687.860 1241.930 1688.000 ;
        RECT 1174.925 1687.660 1175.215 1687.705 ;
        RECT 1187.880 1687.660 1188.020 1687.860 ;
        RECT 1241.610 1687.800 1241.930 1687.860 ;
        RECT 1174.925 1687.520 1188.020 1687.660 ;
        RECT 1174.925 1687.475 1175.215 1687.520 ;
        RECT 180.850 16.900 181.170 16.960 ;
        RECT 196.490 16.900 196.810 16.960 ;
        RECT 180.850 16.760 196.810 16.900 ;
        RECT 180.850 16.700 181.170 16.760 ;
        RECT 196.490 16.700 196.810 16.760 ;
      LAYER via ;
        RECT 196.520 1688.480 196.780 1688.740 ;
        RECT 1241.640 1687.800 1241.900 1688.060 ;
        RECT 180.880 16.700 181.140 16.960 ;
        RECT 196.520 16.700 196.780 16.960 ;
      LAYER met2 ;
        RECT 1241.560 1700.000 1241.840 1704.000 ;
        RECT 196.520 1688.450 196.780 1688.770 ;
        RECT 196.580 16.990 196.720 1688.450 ;
        RECT 1241.700 1688.090 1241.840 1700.000 ;
        RECT 1241.640 1687.770 1241.900 1688.090 ;
        RECT 180.880 16.670 181.140 16.990 ;
        RECT 196.520 16.670 196.780 16.990 ;
        RECT 180.940 2.400 181.080 16.670 ;
        RECT 180.730 -4.800 181.290 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 198.790 18.940 199.110 19.000 ;
        RECT 1248.970 18.940 1249.290 19.000 ;
        RECT 198.790 18.800 1249.290 18.940 ;
        RECT 198.790 18.740 199.110 18.800 ;
        RECT 1248.970 18.740 1249.290 18.800 ;
      LAYER via ;
        RECT 198.820 18.740 199.080 19.000 ;
        RECT 1249.000 18.740 1249.260 19.000 ;
      LAYER met2 ;
        RECT 1250.760 1700.410 1251.040 1704.000 ;
        RECT 1249.060 1700.270 1251.040 1700.410 ;
        RECT 1249.060 19.030 1249.200 1700.270 ;
        RECT 1250.760 1700.000 1251.040 1700.270 ;
        RECT 198.820 18.710 199.080 19.030 ;
        RECT 1249.000 18.710 1249.260 19.030 ;
        RECT 198.880 2.400 199.020 18.710 ;
        RECT 198.670 -4.800 199.230 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 306.890 1686.640 307.210 1686.700 ;
        RECT 1258.630 1686.640 1258.950 1686.700 ;
        RECT 306.890 1686.500 1258.950 1686.640 ;
        RECT 306.890 1686.440 307.210 1686.500 ;
        RECT 1258.630 1686.440 1258.950 1686.500 ;
        RECT 251.780 16.760 291.480 16.900 ;
        RECT 216.730 16.220 217.050 16.280 ;
        RECT 251.780 16.220 251.920 16.760 ;
        RECT 291.340 16.560 291.480 16.760 ;
        RECT 306.890 16.560 307.210 16.620 ;
        RECT 291.340 16.420 307.210 16.560 ;
        RECT 306.890 16.360 307.210 16.420 ;
        RECT 216.730 16.080 251.920 16.220 ;
        RECT 216.730 16.020 217.050 16.080 ;
      LAYER via ;
        RECT 306.920 1686.440 307.180 1686.700 ;
        RECT 1258.660 1686.440 1258.920 1686.700 ;
        RECT 216.760 16.020 217.020 16.280 ;
        RECT 306.920 16.360 307.180 16.620 ;
      LAYER met2 ;
        RECT 1259.960 1700.410 1260.240 1704.000 ;
        RECT 1258.720 1700.270 1260.240 1700.410 ;
        RECT 1258.720 1686.730 1258.860 1700.270 ;
        RECT 1259.960 1700.000 1260.240 1700.270 ;
        RECT 306.920 1686.410 307.180 1686.730 ;
        RECT 1258.660 1686.410 1258.920 1686.730 ;
        RECT 306.980 16.650 307.120 1686.410 ;
        RECT 306.920 16.330 307.180 16.650 ;
        RECT 216.760 15.990 217.020 16.310 ;
        RECT 216.820 2.400 216.960 15.990 ;
        RECT 216.610 -4.800 217.170 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1263.765 1400.885 1263.935 1448.995 ;
        RECT 1263.765 1304.325 1263.935 1352.435 ;
        RECT 1263.765 869.465 1263.935 894.115 ;
        RECT 1263.765 531.505 1263.935 596.955 ;
        RECT 1263.765 158.185 1263.935 200.855 ;
        RECT 1264.225 96.645 1264.395 144.755 ;
        RECT 1263.765 58.565 1263.935 62.815 ;
      LAYER mcon ;
        RECT 1263.765 1448.825 1263.935 1448.995 ;
        RECT 1263.765 1352.265 1263.935 1352.435 ;
        RECT 1263.765 893.945 1263.935 894.115 ;
        RECT 1263.765 596.785 1263.935 596.955 ;
        RECT 1263.765 200.685 1263.935 200.855 ;
        RECT 1264.225 144.585 1264.395 144.755 ;
        RECT 1263.765 62.645 1263.935 62.815 ;
      LAYER met1 ;
        RECT 1263.690 1673.040 1264.010 1673.100 ;
        RECT 1266.450 1673.040 1266.770 1673.100 ;
        RECT 1263.690 1672.900 1266.770 1673.040 ;
        RECT 1263.690 1672.840 1264.010 1672.900 ;
        RECT 1266.450 1672.840 1266.770 1672.900 ;
        RECT 1263.690 1594.500 1264.010 1594.560 ;
        RECT 1262.860 1594.360 1264.010 1594.500 ;
        RECT 1262.860 1594.220 1263.000 1594.360 ;
        RECT 1263.690 1594.300 1264.010 1594.360 ;
        RECT 1262.770 1593.960 1263.090 1594.220 ;
        RECT 1262.770 1545.880 1263.090 1545.940 ;
        RECT 1263.690 1545.880 1264.010 1545.940 ;
        RECT 1262.770 1545.740 1264.010 1545.880 ;
        RECT 1262.770 1545.680 1263.090 1545.740 ;
        RECT 1263.690 1545.680 1264.010 1545.740 ;
        RECT 1263.690 1448.980 1264.010 1449.040 ;
        RECT 1263.495 1448.840 1264.010 1448.980 ;
        RECT 1263.690 1448.780 1264.010 1448.840 ;
        RECT 1263.690 1401.040 1264.010 1401.100 ;
        RECT 1263.495 1400.900 1264.010 1401.040 ;
        RECT 1263.690 1400.840 1264.010 1400.900 ;
        RECT 1263.690 1352.420 1264.010 1352.480 ;
        RECT 1263.495 1352.280 1264.010 1352.420 ;
        RECT 1263.690 1352.220 1264.010 1352.280 ;
        RECT 1263.690 1304.480 1264.010 1304.540 ;
        RECT 1263.495 1304.340 1264.010 1304.480 ;
        RECT 1263.690 1304.280 1264.010 1304.340 ;
        RECT 1263.690 1111.020 1264.010 1111.080 ;
        RECT 1264.610 1111.020 1264.930 1111.080 ;
        RECT 1263.690 1110.880 1264.930 1111.020 ;
        RECT 1263.690 1110.820 1264.010 1110.880 ;
        RECT 1264.610 1110.820 1264.930 1110.880 ;
        RECT 1263.690 1062.740 1264.010 1062.800 ;
        RECT 1264.150 1062.740 1264.470 1062.800 ;
        RECT 1263.690 1062.600 1264.470 1062.740 ;
        RECT 1263.690 1062.540 1264.010 1062.600 ;
        RECT 1264.150 1062.540 1264.470 1062.600 ;
        RECT 1264.150 966.180 1264.470 966.240 ;
        RECT 1265.070 966.180 1265.390 966.240 ;
        RECT 1264.150 966.040 1265.390 966.180 ;
        RECT 1264.150 965.980 1264.470 966.040 ;
        RECT 1265.070 965.980 1265.390 966.040 ;
        RECT 1264.150 917.900 1264.470 917.960 ;
        RECT 1265.070 917.900 1265.390 917.960 ;
        RECT 1264.150 917.760 1265.390 917.900 ;
        RECT 1264.150 917.700 1264.470 917.760 ;
        RECT 1265.070 917.700 1265.390 917.760 ;
        RECT 1263.705 894.100 1263.995 894.145 ;
        RECT 1264.150 894.100 1264.470 894.160 ;
        RECT 1263.705 893.960 1264.470 894.100 ;
        RECT 1263.705 893.915 1263.995 893.960 ;
        RECT 1264.150 893.900 1264.470 893.960 ;
        RECT 1263.690 869.620 1264.010 869.680 ;
        RECT 1263.495 869.480 1264.010 869.620 ;
        RECT 1263.690 869.420 1264.010 869.480 ;
        RECT 1262.770 790.060 1263.090 790.120 ;
        RECT 1263.690 790.060 1264.010 790.120 ;
        RECT 1262.770 789.920 1264.010 790.060 ;
        RECT 1262.770 789.860 1263.090 789.920 ;
        RECT 1263.690 789.860 1264.010 789.920 ;
        RECT 1263.690 724.780 1264.010 724.840 ;
        RECT 1264.150 724.780 1264.470 724.840 ;
        RECT 1263.690 724.640 1264.470 724.780 ;
        RECT 1263.690 724.580 1264.010 724.640 ;
        RECT 1264.150 724.580 1264.470 724.640 ;
        RECT 1263.690 717.640 1264.010 717.700 ;
        RECT 1264.610 717.640 1264.930 717.700 ;
        RECT 1263.690 717.500 1264.930 717.640 ;
        RECT 1263.690 717.440 1264.010 717.500 ;
        RECT 1264.610 717.440 1264.930 717.500 ;
        RECT 1262.770 596.940 1263.090 597.000 ;
        RECT 1263.705 596.940 1263.995 596.985 ;
        RECT 1262.770 596.800 1263.995 596.940 ;
        RECT 1262.770 596.740 1263.090 596.800 ;
        RECT 1263.705 596.755 1263.995 596.800 ;
        RECT 1263.690 531.660 1264.010 531.720 ;
        RECT 1263.495 531.520 1264.010 531.660 ;
        RECT 1263.690 531.460 1264.010 531.520 ;
        RECT 1263.690 200.840 1264.010 200.900 ;
        RECT 1263.495 200.700 1264.010 200.840 ;
        RECT 1263.690 200.640 1264.010 200.700 ;
        RECT 1263.705 158.340 1263.995 158.385 ;
        RECT 1264.150 158.340 1264.470 158.400 ;
        RECT 1263.705 158.200 1264.470 158.340 ;
        RECT 1263.705 158.155 1263.995 158.200 ;
        RECT 1264.150 158.140 1264.470 158.200 ;
        RECT 1264.150 144.740 1264.470 144.800 ;
        RECT 1263.955 144.600 1264.470 144.740 ;
        RECT 1264.150 144.540 1264.470 144.600 ;
        RECT 1264.150 96.800 1264.470 96.860 ;
        RECT 1263.955 96.660 1264.470 96.800 ;
        RECT 1264.150 96.600 1264.470 96.660 ;
        RECT 1263.705 62.800 1263.995 62.845 ;
        RECT 1264.150 62.800 1264.470 62.860 ;
        RECT 1263.705 62.660 1264.470 62.800 ;
        RECT 1263.705 62.615 1263.995 62.660 ;
        RECT 1264.150 62.600 1264.470 62.660 ;
        RECT 1263.690 58.720 1264.010 58.780 ;
        RECT 1263.495 58.580 1264.010 58.720 ;
        RECT 1263.690 58.520 1264.010 58.580 ;
        RECT 234.670 19.960 234.990 20.020 ;
        RECT 1263.690 19.960 1264.010 20.020 ;
        RECT 234.670 19.820 1264.010 19.960 ;
        RECT 234.670 19.760 234.990 19.820 ;
        RECT 1263.690 19.760 1264.010 19.820 ;
      LAYER via ;
        RECT 1263.720 1672.840 1263.980 1673.100 ;
        RECT 1266.480 1672.840 1266.740 1673.100 ;
        RECT 1263.720 1594.300 1263.980 1594.560 ;
        RECT 1262.800 1593.960 1263.060 1594.220 ;
        RECT 1262.800 1545.680 1263.060 1545.940 ;
        RECT 1263.720 1545.680 1263.980 1545.940 ;
        RECT 1263.720 1448.780 1263.980 1449.040 ;
        RECT 1263.720 1400.840 1263.980 1401.100 ;
        RECT 1263.720 1352.220 1263.980 1352.480 ;
        RECT 1263.720 1304.280 1263.980 1304.540 ;
        RECT 1263.720 1110.820 1263.980 1111.080 ;
        RECT 1264.640 1110.820 1264.900 1111.080 ;
        RECT 1263.720 1062.540 1263.980 1062.800 ;
        RECT 1264.180 1062.540 1264.440 1062.800 ;
        RECT 1264.180 965.980 1264.440 966.240 ;
        RECT 1265.100 965.980 1265.360 966.240 ;
        RECT 1264.180 917.700 1264.440 917.960 ;
        RECT 1265.100 917.700 1265.360 917.960 ;
        RECT 1264.180 893.900 1264.440 894.160 ;
        RECT 1263.720 869.420 1263.980 869.680 ;
        RECT 1262.800 789.860 1263.060 790.120 ;
        RECT 1263.720 789.860 1263.980 790.120 ;
        RECT 1263.720 724.580 1263.980 724.840 ;
        RECT 1264.180 724.580 1264.440 724.840 ;
        RECT 1263.720 717.440 1263.980 717.700 ;
        RECT 1264.640 717.440 1264.900 717.700 ;
        RECT 1262.800 596.740 1263.060 597.000 ;
        RECT 1263.720 531.460 1263.980 531.720 ;
        RECT 1263.720 200.640 1263.980 200.900 ;
        RECT 1264.180 158.140 1264.440 158.400 ;
        RECT 1264.180 144.540 1264.440 144.800 ;
        RECT 1264.180 96.600 1264.440 96.860 ;
        RECT 1264.180 62.600 1264.440 62.860 ;
        RECT 1263.720 58.520 1263.980 58.780 ;
        RECT 234.700 19.760 234.960 20.020 ;
        RECT 1263.720 19.760 1263.980 20.020 ;
      LAYER met2 ;
        RECT 1269.160 1700.410 1269.440 1704.000 ;
        RECT 1266.540 1700.270 1269.440 1700.410 ;
        RECT 1266.540 1673.130 1266.680 1700.270 ;
        RECT 1269.160 1700.000 1269.440 1700.270 ;
        RECT 1263.720 1672.810 1263.980 1673.130 ;
        RECT 1266.480 1672.810 1266.740 1673.130 ;
        RECT 1263.780 1594.590 1263.920 1672.810 ;
        RECT 1263.720 1594.270 1263.980 1594.590 ;
        RECT 1262.800 1593.930 1263.060 1594.250 ;
        RECT 1262.860 1545.970 1263.000 1593.930 ;
        RECT 1262.800 1545.650 1263.060 1545.970 ;
        RECT 1263.720 1545.650 1263.980 1545.970 ;
        RECT 1263.780 1449.070 1263.920 1545.650 ;
        RECT 1263.720 1448.750 1263.980 1449.070 ;
        RECT 1263.720 1400.810 1263.980 1401.130 ;
        RECT 1263.780 1352.510 1263.920 1400.810 ;
        RECT 1263.720 1352.190 1263.980 1352.510 ;
        RECT 1263.720 1304.250 1263.980 1304.570 ;
        RECT 1263.780 1207.410 1263.920 1304.250 ;
        RECT 1263.780 1207.270 1264.380 1207.410 ;
        RECT 1264.240 1159.810 1264.380 1207.270 ;
        RECT 1263.780 1159.670 1264.380 1159.810 ;
        RECT 1263.780 1159.245 1263.920 1159.670 ;
        RECT 1263.710 1158.875 1263.990 1159.245 ;
        RECT 1264.630 1158.875 1264.910 1159.245 ;
        RECT 1263.780 1111.110 1263.920 1111.265 ;
        RECT 1264.700 1111.110 1264.840 1158.875 ;
        RECT 1263.720 1110.850 1263.980 1111.110 ;
        RECT 1263.720 1110.790 1264.380 1110.850 ;
        RECT 1264.640 1110.790 1264.900 1111.110 ;
        RECT 1263.780 1110.710 1264.380 1110.790 ;
        RECT 1264.240 1062.830 1264.380 1110.710 ;
        RECT 1263.720 1062.685 1263.980 1062.830 ;
        RECT 1263.710 1062.315 1263.990 1062.685 ;
        RECT 1264.180 1062.510 1264.440 1062.830 ;
        RECT 1264.630 1062.315 1264.910 1062.685 ;
        RECT 1264.700 1027.890 1264.840 1062.315 ;
        RECT 1264.240 1027.750 1264.840 1027.890 ;
        RECT 1264.240 1014.405 1264.380 1027.750 ;
        RECT 1264.170 1014.035 1264.450 1014.405 ;
        RECT 1265.090 1014.035 1265.370 1014.405 ;
        RECT 1265.160 966.270 1265.300 1014.035 ;
        RECT 1264.180 966.125 1264.440 966.270 ;
        RECT 1265.100 966.125 1265.360 966.270 ;
        RECT 1264.170 965.755 1264.450 966.125 ;
        RECT 1265.090 965.755 1265.370 966.125 ;
        RECT 1265.160 917.990 1265.300 965.755 ;
        RECT 1264.180 917.670 1264.440 917.990 ;
        RECT 1265.100 917.670 1265.360 917.990 ;
        RECT 1264.240 894.190 1264.380 917.670 ;
        RECT 1264.180 893.870 1264.440 894.190 ;
        RECT 1263.720 869.390 1263.980 869.710 ;
        RECT 1263.780 790.150 1263.920 869.390 ;
        RECT 1262.800 789.830 1263.060 790.150 ;
        RECT 1263.720 789.830 1263.980 790.150 ;
        RECT 1262.860 766.205 1263.000 789.830 ;
        RECT 1262.790 765.835 1263.070 766.205 ;
        RECT 1264.170 765.835 1264.450 766.205 ;
        RECT 1264.240 724.870 1264.380 765.835 ;
        RECT 1263.720 724.550 1263.980 724.870 ;
        RECT 1264.180 724.550 1264.440 724.870 ;
        RECT 1263.780 717.730 1263.920 724.550 ;
        RECT 1263.720 717.410 1263.980 717.730 ;
        RECT 1264.640 717.410 1264.900 717.730 ;
        RECT 1264.700 628.165 1264.840 717.410 ;
        RECT 1264.630 627.795 1264.910 628.165 ;
        RECT 1262.790 626.435 1263.070 626.805 ;
        RECT 1262.860 597.030 1263.000 626.435 ;
        RECT 1262.800 596.710 1263.060 597.030 ;
        RECT 1263.720 531.430 1263.980 531.750 ;
        RECT 1263.780 200.930 1263.920 531.430 ;
        RECT 1263.720 200.610 1263.980 200.930 ;
        RECT 1264.180 158.110 1264.440 158.430 ;
        RECT 1264.240 144.830 1264.380 158.110 ;
        RECT 1264.180 144.510 1264.440 144.830 ;
        RECT 1264.180 96.570 1264.440 96.890 ;
        RECT 1264.240 62.890 1264.380 96.570 ;
        RECT 1264.180 62.570 1264.440 62.890 ;
        RECT 1263.720 58.490 1263.980 58.810 ;
        RECT 1263.780 20.050 1263.920 58.490 ;
        RECT 234.700 19.730 234.960 20.050 ;
        RECT 1263.720 19.730 1263.980 20.050 ;
        RECT 234.760 2.400 234.900 19.730 ;
        RECT 234.550 -4.800 235.110 2.400 ;
      LAYER via2 ;
        RECT 1263.710 1158.920 1263.990 1159.200 ;
        RECT 1264.630 1158.920 1264.910 1159.200 ;
        RECT 1263.710 1062.360 1263.990 1062.640 ;
        RECT 1264.630 1062.360 1264.910 1062.640 ;
        RECT 1264.170 1014.080 1264.450 1014.360 ;
        RECT 1265.090 1014.080 1265.370 1014.360 ;
        RECT 1264.170 965.800 1264.450 966.080 ;
        RECT 1265.090 965.800 1265.370 966.080 ;
        RECT 1262.790 765.880 1263.070 766.160 ;
        RECT 1264.170 765.880 1264.450 766.160 ;
        RECT 1264.630 627.840 1264.910 628.120 ;
        RECT 1262.790 626.480 1263.070 626.760 ;
      LAYER met3 ;
        RECT 1263.685 1159.210 1264.015 1159.225 ;
        RECT 1264.605 1159.210 1264.935 1159.225 ;
        RECT 1263.685 1158.910 1264.935 1159.210 ;
        RECT 1263.685 1158.895 1264.015 1158.910 ;
        RECT 1264.605 1158.895 1264.935 1158.910 ;
        RECT 1263.685 1062.650 1264.015 1062.665 ;
        RECT 1264.605 1062.650 1264.935 1062.665 ;
        RECT 1263.685 1062.350 1264.935 1062.650 ;
        RECT 1263.685 1062.335 1264.015 1062.350 ;
        RECT 1264.605 1062.335 1264.935 1062.350 ;
        RECT 1264.145 1014.370 1264.475 1014.385 ;
        RECT 1265.065 1014.370 1265.395 1014.385 ;
        RECT 1264.145 1014.070 1265.395 1014.370 ;
        RECT 1264.145 1014.055 1264.475 1014.070 ;
        RECT 1265.065 1014.055 1265.395 1014.070 ;
        RECT 1264.145 966.090 1264.475 966.105 ;
        RECT 1265.065 966.090 1265.395 966.105 ;
        RECT 1264.145 965.790 1265.395 966.090 ;
        RECT 1264.145 965.775 1264.475 965.790 ;
        RECT 1265.065 965.775 1265.395 965.790 ;
        RECT 1262.765 766.170 1263.095 766.185 ;
        RECT 1264.145 766.170 1264.475 766.185 ;
        RECT 1262.765 765.870 1264.475 766.170 ;
        RECT 1262.765 765.855 1263.095 765.870 ;
        RECT 1264.145 765.855 1264.475 765.870 ;
        RECT 1264.605 628.130 1264.935 628.145 ;
        RECT 1263.470 627.830 1264.935 628.130 ;
        RECT 1262.765 626.770 1263.095 626.785 ;
        RECT 1263.470 626.770 1263.770 627.830 ;
        RECT 1264.605 627.815 1264.935 627.830 ;
        RECT 1262.765 626.470 1263.770 626.770 ;
        RECT 1262.765 626.455 1263.095 626.470 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1140.485 1686.995 1140.655 1687.675 ;
        RECT 1140.485 1686.825 1141.575 1686.995 ;
      LAYER mcon ;
        RECT 1140.485 1687.505 1140.655 1687.675 ;
        RECT 1141.405 1686.825 1141.575 1686.995 ;
      LAYER met1 ;
        RECT 86.090 1687.660 86.410 1687.720 ;
        RECT 1140.425 1687.660 1140.715 1687.705 ;
        RECT 86.090 1687.520 1140.715 1687.660 ;
        RECT 86.090 1687.460 86.410 1687.520 ;
        RECT 1140.425 1687.475 1140.715 1687.520 ;
        RECT 1141.345 1686.980 1141.635 1687.025 ;
        RECT 1177.210 1686.980 1177.530 1687.040 ;
        RECT 1141.345 1686.840 1177.530 1686.980 ;
        RECT 1141.345 1686.795 1141.635 1686.840 ;
        RECT 1177.210 1686.780 1177.530 1686.840 ;
        RECT 56.190 16.560 56.510 16.620 ;
        RECT 86.090 16.560 86.410 16.620 ;
        RECT 56.190 16.420 86.410 16.560 ;
        RECT 56.190 16.360 56.510 16.420 ;
        RECT 86.090 16.360 86.410 16.420 ;
      LAYER via ;
        RECT 86.120 1687.460 86.380 1687.720 ;
        RECT 1177.240 1686.780 1177.500 1687.040 ;
        RECT 56.220 16.360 56.480 16.620 ;
        RECT 86.120 16.360 86.380 16.620 ;
      LAYER met2 ;
        RECT 1177.160 1700.000 1177.440 1704.000 ;
        RECT 86.120 1687.430 86.380 1687.750 ;
        RECT 86.180 16.650 86.320 1687.430 ;
        RECT 1177.300 1687.070 1177.440 1700.000 ;
        RECT 1177.240 1686.750 1177.500 1687.070 ;
        RECT 56.220 16.330 56.480 16.650 ;
        RECT 86.120 16.330 86.380 16.650 ;
        RECT 56.280 2.400 56.420 16.330 ;
        RECT 56.070 -4.800 56.630 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 80.110 17.580 80.430 17.640 ;
        RECT 1187.790 17.580 1188.110 17.640 ;
        RECT 80.110 17.440 1188.110 17.580 ;
        RECT 80.110 17.380 80.430 17.440 ;
        RECT 1187.790 17.380 1188.110 17.440 ;
      LAYER via ;
        RECT 80.140 17.380 80.400 17.640 ;
        RECT 1187.820 17.380 1188.080 17.640 ;
      LAYER met2 ;
        RECT 1189.580 1700.410 1189.860 1704.000 ;
        RECT 1187.880 1700.270 1189.860 1700.410 ;
        RECT 1187.880 17.670 1188.020 1700.270 ;
        RECT 1189.580 1700.000 1189.860 1700.270 ;
        RECT 80.140 17.350 80.400 17.670 ;
        RECT 1187.820 17.350 1188.080 17.670 ;
        RECT 80.200 2.400 80.340 17.350 ;
        RECT 79.990 -4.800 80.550 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1184.185 1687.845 1184.355 1688.695 ;
      LAYER mcon ;
        RECT 1184.185 1688.525 1184.355 1688.695 ;
      LAYER met1 ;
        RECT 1184.125 1688.680 1184.415 1688.725 ;
        RECT 1202.050 1688.680 1202.370 1688.740 ;
        RECT 1184.125 1688.540 1202.370 1688.680 ;
        RECT 1184.125 1688.495 1184.415 1688.540 ;
        RECT 1202.050 1688.480 1202.370 1688.540 ;
        RECT 141.290 1688.000 141.610 1688.060 ;
        RECT 1184.125 1688.000 1184.415 1688.045 ;
        RECT 141.290 1687.860 1184.415 1688.000 ;
        RECT 141.290 1687.800 141.610 1687.860 ;
        RECT 1184.125 1687.815 1184.415 1687.860 ;
        RECT 103.570 16.560 103.890 16.620 ;
        RECT 141.290 16.560 141.610 16.620 ;
        RECT 103.570 16.420 141.610 16.560 ;
        RECT 103.570 16.360 103.890 16.420 ;
        RECT 141.290 16.360 141.610 16.420 ;
      LAYER via ;
        RECT 1202.080 1688.480 1202.340 1688.740 ;
        RECT 141.320 1687.800 141.580 1688.060 ;
        RECT 103.600 16.360 103.860 16.620 ;
        RECT 141.320 16.360 141.580 16.620 ;
      LAYER met2 ;
        RECT 1202.000 1700.000 1202.280 1704.000 ;
        RECT 1202.140 1688.770 1202.280 1700.000 ;
        RECT 1202.080 1688.450 1202.340 1688.770 ;
        RECT 141.320 1687.770 141.580 1688.090 ;
        RECT 141.380 16.650 141.520 1687.770 ;
        RECT 103.600 16.330 103.860 16.650 ;
        RECT 141.320 16.330 141.580 16.650 ;
        RECT 103.660 2.400 103.800 16.330 ;
        RECT 103.450 -4.800 104.010 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1209.025 1449.165 1209.195 1497.275 ;
        RECT 1209.025 1352.605 1209.195 1400.715 ;
        RECT 1209.025 1256.045 1209.195 1304.155 ;
        RECT 1209.025 386.325 1209.195 434.775 ;
        RECT 1191.085 17.425 1191.255 18.275 ;
      LAYER mcon ;
        RECT 1209.025 1497.105 1209.195 1497.275 ;
        RECT 1209.025 1400.545 1209.195 1400.715 ;
        RECT 1209.025 1303.985 1209.195 1304.155 ;
        RECT 1209.025 434.605 1209.195 434.775 ;
        RECT 1191.085 18.105 1191.255 18.275 ;
      LAYER met1 ;
        RECT 1208.950 1642.440 1209.270 1642.500 ;
        RECT 1211.710 1642.440 1212.030 1642.500 ;
        RECT 1208.950 1642.300 1212.030 1642.440 ;
        RECT 1208.950 1642.240 1209.270 1642.300 ;
        RECT 1211.710 1642.240 1212.030 1642.300 ;
        RECT 1208.950 1497.260 1209.270 1497.320 ;
        RECT 1208.755 1497.120 1209.270 1497.260 ;
        RECT 1208.950 1497.060 1209.270 1497.120 ;
        RECT 1208.950 1449.320 1209.270 1449.380 ;
        RECT 1208.755 1449.180 1209.270 1449.320 ;
        RECT 1208.950 1449.120 1209.270 1449.180 ;
        RECT 1208.950 1400.700 1209.270 1400.760 ;
        RECT 1208.755 1400.560 1209.270 1400.700 ;
        RECT 1208.950 1400.500 1209.270 1400.560 ;
        RECT 1208.950 1352.760 1209.270 1352.820 ;
        RECT 1208.755 1352.620 1209.270 1352.760 ;
        RECT 1208.950 1352.560 1209.270 1352.620 ;
        RECT 1208.950 1304.140 1209.270 1304.200 ;
        RECT 1208.755 1304.000 1209.270 1304.140 ;
        RECT 1208.950 1303.940 1209.270 1304.000 ;
        RECT 1208.950 1256.200 1209.270 1256.260 ;
        RECT 1208.755 1256.060 1209.270 1256.200 ;
        RECT 1208.950 1256.000 1209.270 1256.060 ;
        RECT 1208.950 869.620 1209.270 869.680 ;
        RECT 1209.870 869.620 1210.190 869.680 ;
        RECT 1208.950 869.480 1210.190 869.620 ;
        RECT 1208.950 869.420 1209.270 869.480 ;
        RECT 1209.870 869.420 1210.190 869.480 ;
        RECT 1208.950 531.320 1209.270 531.380 ;
        RECT 1209.870 531.320 1210.190 531.380 ;
        RECT 1208.950 531.180 1210.190 531.320 ;
        RECT 1208.950 531.120 1209.270 531.180 ;
        RECT 1209.870 531.120 1210.190 531.180 ;
        RECT 1208.950 434.760 1209.270 434.820 ;
        RECT 1208.755 434.620 1209.270 434.760 ;
        RECT 1208.950 434.560 1209.270 434.620 ;
        RECT 1208.950 386.480 1209.270 386.540 ;
        RECT 1208.755 386.340 1209.270 386.480 ;
        RECT 1208.950 386.280 1209.270 386.340 ;
        RECT 127.490 18.260 127.810 18.320 ;
        RECT 1191.025 18.260 1191.315 18.305 ;
        RECT 127.490 18.120 1191.315 18.260 ;
        RECT 127.490 18.060 127.810 18.120 ;
        RECT 1191.025 18.075 1191.315 18.120 ;
        RECT 1191.025 17.580 1191.315 17.625 ;
        RECT 1208.950 17.580 1209.270 17.640 ;
        RECT 1191.025 17.440 1209.270 17.580 ;
        RECT 1191.025 17.395 1191.315 17.440 ;
        RECT 1208.950 17.380 1209.270 17.440 ;
      LAYER via ;
        RECT 1208.980 1642.240 1209.240 1642.500 ;
        RECT 1211.740 1642.240 1212.000 1642.500 ;
        RECT 1208.980 1497.060 1209.240 1497.320 ;
        RECT 1208.980 1449.120 1209.240 1449.380 ;
        RECT 1208.980 1400.500 1209.240 1400.760 ;
        RECT 1208.980 1352.560 1209.240 1352.820 ;
        RECT 1208.980 1303.940 1209.240 1304.200 ;
        RECT 1208.980 1256.000 1209.240 1256.260 ;
        RECT 1208.980 869.420 1209.240 869.680 ;
        RECT 1209.900 869.420 1210.160 869.680 ;
        RECT 1208.980 531.120 1209.240 531.380 ;
        RECT 1209.900 531.120 1210.160 531.380 ;
        RECT 1208.980 434.560 1209.240 434.820 ;
        RECT 1208.980 386.280 1209.240 386.540 ;
        RECT 127.520 18.060 127.780 18.320 ;
        RECT 1208.980 17.380 1209.240 17.640 ;
      LAYER met2 ;
        RECT 1213.960 1701.090 1214.240 1704.000 ;
        RECT 1211.800 1700.950 1214.240 1701.090 ;
        RECT 1211.800 1642.530 1211.940 1700.950 ;
        RECT 1213.960 1700.000 1214.240 1700.950 ;
        RECT 1208.980 1642.210 1209.240 1642.530 ;
        RECT 1211.740 1642.210 1212.000 1642.530 ;
        RECT 1209.040 1497.350 1209.180 1642.210 ;
        RECT 1208.980 1497.030 1209.240 1497.350 ;
        RECT 1208.980 1449.090 1209.240 1449.410 ;
        RECT 1209.040 1400.790 1209.180 1449.090 ;
        RECT 1208.980 1400.470 1209.240 1400.790 ;
        RECT 1208.980 1352.530 1209.240 1352.850 ;
        RECT 1209.040 1304.230 1209.180 1352.530 ;
        RECT 1208.980 1303.910 1209.240 1304.230 ;
        RECT 1208.980 1255.970 1209.240 1256.290 ;
        RECT 1209.040 917.845 1209.180 1255.970 ;
        RECT 1208.970 917.475 1209.250 917.845 ;
        RECT 1209.890 917.475 1210.170 917.845 ;
        RECT 1209.960 869.710 1210.100 917.475 ;
        RECT 1208.980 869.390 1209.240 869.710 ;
        RECT 1209.900 869.390 1210.160 869.710 ;
        RECT 1209.040 531.410 1209.180 869.390 ;
        RECT 1208.980 531.090 1209.240 531.410 ;
        RECT 1209.900 531.090 1210.160 531.410 ;
        RECT 1209.960 483.325 1210.100 531.090 ;
        RECT 1208.970 482.955 1209.250 483.325 ;
        RECT 1209.890 482.955 1210.170 483.325 ;
        RECT 1209.040 434.850 1209.180 482.955 ;
        RECT 1208.980 434.530 1209.240 434.850 ;
        RECT 1208.980 386.250 1209.240 386.570 ;
        RECT 127.520 18.030 127.780 18.350 ;
        RECT 127.580 2.400 127.720 18.030 ;
        RECT 1209.040 17.670 1209.180 386.250 ;
        RECT 1208.980 17.350 1209.240 17.670 ;
        RECT 127.370 -4.800 127.930 2.400 ;
      LAYER via2 ;
        RECT 1208.970 917.520 1209.250 917.800 ;
        RECT 1209.890 917.520 1210.170 917.800 ;
        RECT 1208.970 483.000 1209.250 483.280 ;
        RECT 1209.890 483.000 1210.170 483.280 ;
      LAYER met3 ;
        RECT 1208.945 917.810 1209.275 917.825 ;
        RECT 1209.865 917.810 1210.195 917.825 ;
        RECT 1208.945 917.510 1210.195 917.810 ;
        RECT 1208.945 917.495 1209.275 917.510 ;
        RECT 1209.865 917.495 1210.195 917.510 ;
        RECT 1208.945 483.290 1209.275 483.305 ;
        RECT 1209.865 483.290 1210.195 483.305 ;
        RECT 1208.945 482.990 1210.195 483.290 ;
        RECT 1208.945 482.975 1209.275 482.990 ;
        RECT 1209.865 482.975 1210.195 482.990 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 26.290 17.240 26.610 17.300 ;
        RECT 51.590 17.240 51.910 17.300 ;
        RECT 26.290 17.100 51.910 17.240 ;
        RECT 26.290 17.040 26.610 17.100 ;
        RECT 51.590 17.040 51.910 17.100 ;
      LAYER via ;
        RECT 26.320 17.040 26.580 17.300 ;
        RECT 51.620 17.040 51.880 17.300 ;
      LAYER met2 ;
        RECT 1161.980 1700.000 1162.260 1704.000 ;
        RECT 1162.120 1686.925 1162.260 1700.000 ;
        RECT 51.610 1686.555 51.890 1686.925 ;
        RECT 1162.050 1686.555 1162.330 1686.925 ;
        RECT 51.680 17.330 51.820 1686.555 ;
        RECT 26.320 17.010 26.580 17.330 ;
        RECT 51.620 17.010 51.880 17.330 ;
        RECT 26.380 2.400 26.520 17.010 ;
        RECT 26.170 -4.800 26.730 2.400 ;
      LAYER via2 ;
        RECT 51.610 1686.600 51.890 1686.880 ;
        RECT 1162.050 1686.600 1162.330 1686.880 ;
      LAYER met3 ;
        RECT 51.585 1686.890 51.915 1686.905 ;
        RECT 1162.025 1686.890 1162.355 1686.905 ;
        RECT 51.585 1686.590 1162.355 1686.890 ;
        RECT 51.585 1686.575 51.915 1686.590 ;
        RECT 1162.025 1686.575 1162.355 1686.590 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1161.645 1573.265 1161.815 1621.375 ;
        RECT 1161.645 1474.325 1161.815 1566.295 ;
        RECT 1162.105 1414.485 1162.275 1462.595 ;
        RECT 1160.725 1311.125 1160.895 1359.235 ;
        RECT 1159.805 186.405 1159.975 234.515 ;
        RECT 1159.345 131.325 1159.515 179.435 ;
      LAYER mcon ;
        RECT 1161.645 1621.205 1161.815 1621.375 ;
        RECT 1161.645 1566.125 1161.815 1566.295 ;
        RECT 1162.105 1462.425 1162.275 1462.595 ;
        RECT 1160.725 1359.065 1160.895 1359.235 ;
        RECT 1159.805 234.345 1159.975 234.515 ;
        RECT 1159.345 179.265 1159.515 179.435 ;
      LAYER met1 ;
        RECT 1161.110 1642.100 1161.430 1642.160 ;
        RECT 1161.570 1642.100 1161.890 1642.160 ;
        RECT 1161.110 1641.960 1161.890 1642.100 ;
        RECT 1161.110 1641.900 1161.430 1641.960 ;
        RECT 1161.570 1641.900 1161.890 1641.960 ;
        RECT 1161.570 1621.360 1161.890 1621.420 ;
        RECT 1161.375 1621.220 1161.890 1621.360 ;
        RECT 1161.570 1621.160 1161.890 1621.220 ;
        RECT 1161.585 1573.420 1161.875 1573.465 ;
        RECT 1162.030 1573.420 1162.350 1573.480 ;
        RECT 1161.585 1573.280 1162.350 1573.420 ;
        RECT 1161.585 1573.235 1161.875 1573.280 ;
        RECT 1162.030 1573.220 1162.350 1573.280 ;
        RECT 1161.570 1566.280 1161.890 1566.340 ;
        RECT 1161.375 1566.140 1161.890 1566.280 ;
        RECT 1161.570 1566.080 1161.890 1566.140 ;
        RECT 1161.570 1474.480 1161.890 1474.540 ;
        RECT 1161.375 1474.340 1161.890 1474.480 ;
        RECT 1161.570 1474.280 1161.890 1474.340 ;
        RECT 1161.570 1469.720 1161.890 1469.780 ;
        RECT 1162.030 1469.720 1162.350 1469.780 ;
        RECT 1161.570 1469.580 1162.350 1469.720 ;
        RECT 1161.570 1469.520 1161.890 1469.580 ;
        RECT 1162.030 1469.520 1162.350 1469.580 ;
        RECT 1162.030 1462.580 1162.350 1462.640 ;
        RECT 1161.835 1462.440 1162.350 1462.580 ;
        RECT 1162.030 1462.380 1162.350 1462.440 ;
        RECT 1162.030 1414.640 1162.350 1414.700 ;
        RECT 1161.835 1414.500 1162.350 1414.640 ;
        RECT 1162.030 1414.440 1162.350 1414.500 ;
        RECT 1160.650 1366.700 1160.970 1366.760 ;
        RECT 1162.030 1366.700 1162.350 1366.760 ;
        RECT 1160.650 1366.560 1162.350 1366.700 ;
        RECT 1160.650 1366.500 1160.970 1366.560 ;
        RECT 1162.030 1366.500 1162.350 1366.560 ;
        RECT 1160.650 1359.220 1160.970 1359.280 ;
        RECT 1160.455 1359.080 1160.970 1359.220 ;
        RECT 1160.650 1359.020 1160.970 1359.080 ;
        RECT 1160.665 1311.280 1160.955 1311.325 ;
        RECT 1161.570 1311.280 1161.890 1311.340 ;
        RECT 1160.665 1311.140 1161.890 1311.280 ;
        RECT 1160.665 1311.095 1160.955 1311.140 ;
        RECT 1161.570 1311.080 1161.890 1311.140 ;
        RECT 1160.650 1269.800 1160.970 1269.860 ;
        RECT 1161.570 1269.800 1161.890 1269.860 ;
        RECT 1160.650 1269.660 1161.890 1269.800 ;
        RECT 1160.650 1269.600 1160.970 1269.660 ;
        RECT 1161.570 1269.600 1161.890 1269.660 ;
        RECT 1159.730 1221.180 1160.050 1221.240 ;
        RECT 1160.650 1221.180 1160.970 1221.240 ;
        RECT 1159.730 1221.040 1160.970 1221.180 ;
        RECT 1159.730 1220.980 1160.050 1221.040 ;
        RECT 1160.650 1220.980 1160.970 1221.040 ;
        RECT 1159.270 1083.140 1159.590 1083.200 ;
        RECT 1160.190 1083.140 1160.510 1083.200 ;
        RECT 1159.270 1083.000 1160.510 1083.140 ;
        RECT 1159.270 1082.940 1159.590 1083.000 ;
        RECT 1160.190 1082.940 1160.510 1083.000 ;
        RECT 1159.730 959.040 1160.050 959.100 ;
        RECT 1160.190 959.040 1160.510 959.100 ;
        RECT 1159.730 958.900 1160.510 959.040 ;
        RECT 1159.730 958.840 1160.050 958.900 ;
        RECT 1160.190 958.840 1160.510 958.900 ;
        RECT 1159.730 910.760 1160.050 910.820 ;
        RECT 1160.650 910.760 1160.970 910.820 ;
        RECT 1159.730 910.620 1160.970 910.760 ;
        RECT 1159.730 910.560 1160.050 910.620 ;
        RECT 1160.650 910.560 1160.970 910.620 ;
        RECT 1159.730 821.340 1160.050 821.400 ;
        RECT 1160.190 821.340 1160.510 821.400 ;
        RECT 1159.730 821.200 1160.510 821.340 ;
        RECT 1159.730 821.140 1160.050 821.200 ;
        RECT 1160.190 821.140 1160.510 821.200 ;
        RECT 1160.190 786.800 1160.510 787.060 ;
        RECT 1160.280 786.660 1160.420 786.800 ;
        RECT 1160.650 786.660 1160.970 786.720 ;
        RECT 1160.280 786.520 1160.970 786.660 ;
        RECT 1160.650 786.460 1160.970 786.520 ;
        RECT 1159.270 593.540 1159.590 593.600 ;
        RECT 1160.190 593.540 1160.510 593.600 ;
        RECT 1159.270 593.400 1160.510 593.540 ;
        RECT 1159.270 593.340 1159.590 593.400 ;
        RECT 1160.190 593.340 1160.510 593.400 ;
        RECT 1159.270 507.180 1159.590 507.240 ;
        RECT 1160.190 507.180 1160.510 507.240 ;
        RECT 1159.270 507.040 1160.510 507.180 ;
        RECT 1159.270 506.980 1159.590 507.040 ;
        RECT 1160.190 506.980 1160.510 507.040 ;
        RECT 1160.190 386.280 1160.510 386.540 ;
        RECT 1160.280 385.860 1160.420 386.280 ;
        RECT 1160.190 385.600 1160.510 385.860 ;
        RECT 1159.270 337.860 1159.590 337.920 ;
        RECT 1160.190 337.860 1160.510 337.920 ;
        RECT 1159.270 337.720 1160.510 337.860 ;
        RECT 1159.270 337.660 1159.590 337.720 ;
        RECT 1160.190 337.660 1160.510 337.720 ;
        RECT 1159.730 234.500 1160.050 234.560 ;
        RECT 1159.535 234.360 1160.050 234.500 ;
        RECT 1159.730 234.300 1160.050 234.360 ;
        RECT 1159.745 186.560 1160.035 186.605 ;
        RECT 1160.190 186.560 1160.510 186.620 ;
        RECT 1159.745 186.420 1160.510 186.560 ;
        RECT 1159.745 186.375 1160.035 186.420 ;
        RECT 1160.190 186.360 1160.510 186.420 ;
        RECT 1159.285 179.420 1159.575 179.465 ;
        RECT 1160.190 179.420 1160.510 179.480 ;
        RECT 1159.285 179.280 1160.510 179.420 ;
        RECT 1159.285 179.235 1159.575 179.280 ;
        RECT 1160.190 179.220 1160.510 179.280 ;
        RECT 1159.270 131.480 1159.590 131.540 ;
        RECT 1159.075 131.340 1159.590 131.480 ;
        RECT 1159.270 131.280 1159.590 131.340 ;
        RECT 1158.810 130.800 1159.130 130.860 ;
        RECT 1159.270 130.800 1159.590 130.860 ;
        RECT 1158.810 130.660 1159.590 130.800 ;
        RECT 1158.810 130.600 1159.130 130.660 ;
        RECT 1159.270 130.600 1159.590 130.660 ;
      LAYER via ;
        RECT 1161.140 1641.900 1161.400 1642.160 ;
        RECT 1161.600 1641.900 1161.860 1642.160 ;
        RECT 1161.600 1621.160 1161.860 1621.420 ;
        RECT 1162.060 1573.220 1162.320 1573.480 ;
        RECT 1161.600 1566.080 1161.860 1566.340 ;
        RECT 1161.600 1474.280 1161.860 1474.540 ;
        RECT 1161.600 1469.520 1161.860 1469.780 ;
        RECT 1162.060 1469.520 1162.320 1469.780 ;
        RECT 1162.060 1462.380 1162.320 1462.640 ;
        RECT 1162.060 1414.440 1162.320 1414.700 ;
        RECT 1160.680 1366.500 1160.940 1366.760 ;
        RECT 1162.060 1366.500 1162.320 1366.760 ;
        RECT 1160.680 1359.020 1160.940 1359.280 ;
        RECT 1161.600 1311.080 1161.860 1311.340 ;
        RECT 1160.680 1269.600 1160.940 1269.860 ;
        RECT 1161.600 1269.600 1161.860 1269.860 ;
        RECT 1159.760 1220.980 1160.020 1221.240 ;
        RECT 1160.680 1220.980 1160.940 1221.240 ;
        RECT 1159.300 1082.940 1159.560 1083.200 ;
        RECT 1160.220 1082.940 1160.480 1083.200 ;
        RECT 1159.760 958.840 1160.020 959.100 ;
        RECT 1160.220 958.840 1160.480 959.100 ;
        RECT 1159.760 910.560 1160.020 910.820 ;
        RECT 1160.680 910.560 1160.940 910.820 ;
        RECT 1159.760 821.140 1160.020 821.400 ;
        RECT 1160.220 821.140 1160.480 821.400 ;
        RECT 1160.220 786.800 1160.480 787.060 ;
        RECT 1160.680 786.460 1160.940 786.720 ;
        RECT 1159.300 593.340 1159.560 593.600 ;
        RECT 1160.220 593.340 1160.480 593.600 ;
        RECT 1159.300 506.980 1159.560 507.240 ;
        RECT 1160.220 506.980 1160.480 507.240 ;
        RECT 1160.220 386.280 1160.480 386.540 ;
        RECT 1160.220 385.600 1160.480 385.860 ;
        RECT 1159.300 337.660 1159.560 337.920 ;
        RECT 1160.220 337.660 1160.480 337.920 ;
        RECT 1159.760 234.300 1160.020 234.560 ;
        RECT 1160.220 186.360 1160.480 186.620 ;
        RECT 1160.220 179.220 1160.480 179.480 ;
        RECT 1159.300 131.280 1159.560 131.540 ;
        RECT 1158.840 130.600 1159.100 130.860 ;
        RECT 1159.300 130.600 1159.560 130.860 ;
      LAYER met2 ;
        RECT 1165.200 1700.410 1165.480 1704.000 ;
        RECT 1163.040 1700.270 1165.480 1700.410 ;
        RECT 1163.040 1666.410 1163.180 1700.270 ;
        RECT 1165.200 1700.000 1165.480 1700.270 ;
        RECT 1161.200 1666.270 1163.180 1666.410 ;
        RECT 1161.200 1642.190 1161.340 1666.270 ;
        RECT 1161.140 1641.870 1161.400 1642.190 ;
        RECT 1161.600 1641.870 1161.860 1642.190 ;
        RECT 1161.660 1621.450 1161.800 1641.870 ;
        RECT 1161.600 1621.130 1161.860 1621.450 ;
        RECT 1162.120 1573.510 1162.260 1573.665 ;
        RECT 1162.060 1573.250 1162.320 1573.510 ;
        RECT 1161.660 1573.190 1162.320 1573.250 ;
        RECT 1161.660 1573.110 1162.260 1573.190 ;
        RECT 1161.660 1566.370 1161.800 1573.110 ;
        RECT 1161.600 1566.050 1161.860 1566.370 ;
        RECT 1161.600 1474.250 1161.860 1474.570 ;
        RECT 1161.660 1469.810 1161.800 1474.250 ;
        RECT 1161.600 1469.490 1161.860 1469.810 ;
        RECT 1162.060 1469.490 1162.320 1469.810 ;
        RECT 1162.120 1462.670 1162.260 1469.490 ;
        RECT 1162.060 1462.350 1162.320 1462.670 ;
        RECT 1162.060 1414.410 1162.320 1414.730 ;
        RECT 1162.120 1366.790 1162.260 1414.410 ;
        RECT 1160.680 1366.470 1160.940 1366.790 ;
        RECT 1162.060 1366.470 1162.320 1366.790 ;
        RECT 1160.740 1359.310 1160.880 1366.470 ;
        RECT 1160.680 1358.990 1160.940 1359.310 ;
        RECT 1161.600 1311.050 1161.860 1311.370 ;
        RECT 1161.660 1269.890 1161.800 1311.050 ;
        RECT 1160.680 1269.570 1160.940 1269.890 ;
        RECT 1161.600 1269.570 1161.860 1269.890 ;
        RECT 1160.740 1221.270 1160.880 1269.570 ;
        RECT 1159.760 1220.950 1160.020 1221.270 ;
        RECT 1160.680 1220.950 1160.940 1221.270 ;
        RECT 1159.820 1131.930 1159.960 1220.950 ;
        RECT 1159.360 1131.790 1159.960 1131.930 ;
        RECT 1159.360 1125.130 1159.500 1131.790 ;
        RECT 1159.360 1124.990 1160.880 1125.130 ;
        RECT 1160.740 1124.450 1160.880 1124.990 ;
        RECT 1160.280 1124.310 1160.880 1124.450 ;
        RECT 1160.280 1083.230 1160.420 1124.310 ;
        RECT 1159.300 1082.910 1159.560 1083.230 ;
        RECT 1160.220 1082.910 1160.480 1083.230 ;
        RECT 1159.360 1027.890 1159.500 1082.910 ;
        RECT 1159.360 1027.750 1159.960 1027.890 ;
        RECT 1159.820 980.290 1159.960 1027.750 ;
        RECT 1159.820 980.150 1160.420 980.290 ;
        RECT 1160.280 959.130 1160.420 980.150 ;
        RECT 1159.760 958.810 1160.020 959.130 ;
        RECT 1160.220 958.810 1160.480 959.130 ;
        RECT 1159.820 931.330 1159.960 958.810 ;
        RECT 1159.820 931.190 1160.420 931.330 ;
        RECT 1160.280 910.930 1160.420 931.190 ;
        RECT 1160.280 910.850 1160.880 910.930 ;
        RECT 1159.760 910.530 1160.020 910.850 ;
        RECT 1160.280 910.790 1160.940 910.850 ;
        RECT 1160.680 910.530 1160.940 910.790 ;
        RECT 1159.820 821.430 1159.960 910.530 ;
        RECT 1159.760 821.110 1160.020 821.430 ;
        RECT 1160.220 821.110 1160.480 821.430 ;
        RECT 1160.280 787.090 1160.420 821.110 ;
        RECT 1160.220 786.770 1160.480 787.090 ;
        RECT 1160.680 786.430 1160.940 786.750 ;
        RECT 1160.740 738.210 1160.880 786.430 ;
        RECT 1159.820 738.070 1160.880 738.210 ;
        RECT 1159.820 689.930 1159.960 738.070 ;
        RECT 1159.360 689.790 1159.960 689.930 ;
        RECT 1159.360 641.650 1159.500 689.790 ;
        RECT 1159.360 641.510 1160.420 641.650 ;
        RECT 1160.280 593.630 1160.420 641.510 ;
        RECT 1159.300 593.310 1159.560 593.630 ;
        RECT 1160.220 593.310 1160.480 593.630 ;
        RECT 1159.360 545.090 1159.500 593.310 ;
        RECT 1159.360 544.950 1160.420 545.090 ;
        RECT 1160.280 507.270 1160.420 544.950 ;
        RECT 1159.300 506.950 1159.560 507.270 ;
        RECT 1160.220 506.950 1160.480 507.270 ;
        RECT 1159.360 448.530 1159.500 506.950 ;
        RECT 1159.360 448.390 1160.420 448.530 ;
        RECT 1160.280 386.570 1160.420 448.390 ;
        RECT 1160.220 386.250 1160.480 386.570 ;
        RECT 1160.220 385.570 1160.480 385.890 ;
        RECT 1160.280 337.950 1160.420 385.570 ;
        RECT 1159.300 337.630 1159.560 337.950 ;
        RECT 1160.220 337.630 1160.480 337.950 ;
        RECT 1159.360 307.090 1159.500 337.630 ;
        RECT 1159.360 306.950 1160.880 307.090 ;
        RECT 1160.740 289.410 1160.880 306.950 ;
        RECT 1160.280 289.270 1160.880 289.410 ;
        RECT 1160.280 264.930 1160.420 289.270 ;
        RECT 1159.820 264.790 1160.420 264.930 ;
        RECT 1159.820 234.590 1159.960 264.790 ;
        RECT 1159.760 234.270 1160.020 234.590 ;
        RECT 1160.220 186.330 1160.480 186.650 ;
        RECT 1160.280 179.510 1160.420 186.330 ;
        RECT 1160.220 179.190 1160.480 179.510 ;
        RECT 1159.300 131.250 1159.560 131.570 ;
        RECT 1159.360 130.890 1159.500 131.250 ;
        RECT 1158.840 130.570 1159.100 130.890 ;
        RECT 1159.300 130.570 1159.560 130.890 ;
        RECT 1158.900 107.170 1159.040 130.570 ;
        RECT 1158.900 107.030 1159.500 107.170 ;
        RECT 1159.360 16.845 1159.500 107.030 ;
        RECT 32.290 16.475 32.570 16.845 ;
        RECT 1159.290 16.475 1159.570 16.845 ;
        RECT 32.360 2.400 32.500 16.475 ;
        RECT 32.150 -4.800 32.710 2.400 ;
      LAYER via2 ;
        RECT 32.290 16.520 32.570 16.800 ;
        RECT 1159.290 16.520 1159.570 16.800 ;
      LAYER met3 ;
        RECT 32.265 16.810 32.595 16.825 ;
        RECT 1159.265 16.810 1159.595 16.825 ;
        RECT 32.265 16.510 1159.595 16.810 ;
        RECT 32.265 16.495 32.595 16.510 ;
        RECT 1159.265 16.495 1159.595 16.510 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -9.980 -4.620 -6.980 3524.300 ;
        RECT 4.020 -9.220 7.020 3528.900 ;
        RECT 184.020 -9.220 187.020 3528.900 ;
        RECT 364.020 -9.220 367.020 3528.900 ;
        RECT 544.020 -9.220 547.020 3528.900 ;
        RECT 724.020 -9.220 727.020 3528.900 ;
        RECT 904.020 -9.220 907.020 3528.900 ;
        RECT 1084.020 -9.220 1087.020 3528.900 ;
        RECT 1264.020 -9.220 1267.020 3528.900 ;
        RECT 1444.020 -9.220 1447.020 3528.900 ;
        RECT 1624.020 -9.220 1627.020 3528.900 ;
        RECT 1804.020 -9.220 1807.020 3528.900 ;
        RECT 1984.020 -9.220 1987.020 3528.900 ;
        RECT 2164.020 -9.220 2167.020 3528.900 ;
        RECT 2344.020 -9.220 2347.020 3528.900 ;
        RECT 2524.020 -9.220 2527.020 3528.900 ;
        RECT 2704.020 -9.220 2707.020 3528.900 ;
        RECT 2884.020 -9.220 2887.020 3528.900 ;
        RECT 2926.600 -4.620 2929.600 3524.300 ;
      LAYER via4 ;
        RECT -9.070 3523.010 -7.890 3524.190 ;
        RECT -9.070 3521.410 -7.890 3522.590 ;
        RECT -9.070 3431.090 -7.890 3432.270 ;
        RECT -9.070 3429.490 -7.890 3430.670 ;
        RECT -9.070 3251.090 -7.890 3252.270 ;
        RECT -9.070 3249.490 -7.890 3250.670 ;
        RECT -9.070 3071.090 -7.890 3072.270 ;
        RECT -9.070 3069.490 -7.890 3070.670 ;
        RECT -9.070 2891.090 -7.890 2892.270 ;
        RECT -9.070 2889.490 -7.890 2890.670 ;
        RECT -9.070 2711.090 -7.890 2712.270 ;
        RECT -9.070 2709.490 -7.890 2710.670 ;
        RECT -9.070 2531.090 -7.890 2532.270 ;
        RECT -9.070 2529.490 -7.890 2530.670 ;
        RECT -9.070 2351.090 -7.890 2352.270 ;
        RECT -9.070 2349.490 -7.890 2350.670 ;
        RECT -9.070 2171.090 -7.890 2172.270 ;
        RECT -9.070 2169.490 -7.890 2170.670 ;
        RECT -9.070 1991.090 -7.890 1992.270 ;
        RECT -9.070 1989.490 -7.890 1990.670 ;
        RECT -9.070 1811.090 -7.890 1812.270 ;
        RECT -9.070 1809.490 -7.890 1810.670 ;
        RECT -9.070 1631.090 -7.890 1632.270 ;
        RECT -9.070 1629.490 -7.890 1630.670 ;
        RECT -9.070 1451.090 -7.890 1452.270 ;
        RECT -9.070 1449.490 -7.890 1450.670 ;
        RECT -9.070 1271.090 -7.890 1272.270 ;
        RECT -9.070 1269.490 -7.890 1270.670 ;
        RECT -9.070 1091.090 -7.890 1092.270 ;
        RECT -9.070 1089.490 -7.890 1090.670 ;
        RECT -9.070 911.090 -7.890 912.270 ;
        RECT -9.070 909.490 -7.890 910.670 ;
        RECT -9.070 731.090 -7.890 732.270 ;
        RECT -9.070 729.490 -7.890 730.670 ;
        RECT -9.070 551.090 -7.890 552.270 ;
        RECT -9.070 549.490 -7.890 550.670 ;
        RECT -9.070 371.090 -7.890 372.270 ;
        RECT -9.070 369.490 -7.890 370.670 ;
        RECT -9.070 191.090 -7.890 192.270 ;
        RECT -9.070 189.490 -7.890 190.670 ;
        RECT -9.070 11.090 -7.890 12.270 ;
        RECT -9.070 9.490 -7.890 10.670 ;
        RECT -9.070 -2.910 -7.890 -1.730 ;
        RECT -9.070 -4.510 -7.890 -3.330 ;
        RECT 4.930 3523.010 6.110 3524.190 ;
        RECT 4.930 3521.410 6.110 3522.590 ;
        RECT 4.930 3431.090 6.110 3432.270 ;
        RECT 4.930 3429.490 6.110 3430.670 ;
        RECT 4.930 3251.090 6.110 3252.270 ;
        RECT 4.930 3249.490 6.110 3250.670 ;
        RECT 4.930 3071.090 6.110 3072.270 ;
        RECT 4.930 3069.490 6.110 3070.670 ;
        RECT 4.930 2891.090 6.110 2892.270 ;
        RECT 4.930 2889.490 6.110 2890.670 ;
        RECT 4.930 2711.090 6.110 2712.270 ;
        RECT 4.930 2709.490 6.110 2710.670 ;
        RECT 4.930 2531.090 6.110 2532.270 ;
        RECT 4.930 2529.490 6.110 2530.670 ;
        RECT 4.930 2351.090 6.110 2352.270 ;
        RECT 4.930 2349.490 6.110 2350.670 ;
        RECT 4.930 2171.090 6.110 2172.270 ;
        RECT 4.930 2169.490 6.110 2170.670 ;
        RECT 4.930 1991.090 6.110 1992.270 ;
        RECT 4.930 1989.490 6.110 1990.670 ;
        RECT 4.930 1811.090 6.110 1812.270 ;
        RECT 4.930 1809.490 6.110 1810.670 ;
        RECT 4.930 1631.090 6.110 1632.270 ;
        RECT 4.930 1629.490 6.110 1630.670 ;
        RECT 4.930 1451.090 6.110 1452.270 ;
        RECT 4.930 1449.490 6.110 1450.670 ;
        RECT 4.930 1271.090 6.110 1272.270 ;
        RECT 4.930 1269.490 6.110 1270.670 ;
        RECT 4.930 1091.090 6.110 1092.270 ;
        RECT 4.930 1089.490 6.110 1090.670 ;
        RECT 4.930 911.090 6.110 912.270 ;
        RECT 4.930 909.490 6.110 910.670 ;
        RECT 4.930 731.090 6.110 732.270 ;
        RECT 4.930 729.490 6.110 730.670 ;
        RECT 4.930 551.090 6.110 552.270 ;
        RECT 4.930 549.490 6.110 550.670 ;
        RECT 4.930 371.090 6.110 372.270 ;
        RECT 4.930 369.490 6.110 370.670 ;
        RECT 4.930 191.090 6.110 192.270 ;
        RECT 4.930 189.490 6.110 190.670 ;
        RECT 4.930 11.090 6.110 12.270 ;
        RECT 4.930 9.490 6.110 10.670 ;
        RECT 4.930 -2.910 6.110 -1.730 ;
        RECT 4.930 -4.510 6.110 -3.330 ;
        RECT 184.930 3523.010 186.110 3524.190 ;
        RECT 184.930 3521.410 186.110 3522.590 ;
        RECT 184.930 3431.090 186.110 3432.270 ;
        RECT 184.930 3429.490 186.110 3430.670 ;
        RECT 184.930 3251.090 186.110 3252.270 ;
        RECT 184.930 3249.490 186.110 3250.670 ;
        RECT 184.930 3071.090 186.110 3072.270 ;
        RECT 184.930 3069.490 186.110 3070.670 ;
        RECT 184.930 2891.090 186.110 2892.270 ;
        RECT 184.930 2889.490 186.110 2890.670 ;
        RECT 184.930 2711.090 186.110 2712.270 ;
        RECT 184.930 2709.490 186.110 2710.670 ;
        RECT 184.930 2531.090 186.110 2532.270 ;
        RECT 184.930 2529.490 186.110 2530.670 ;
        RECT 184.930 2351.090 186.110 2352.270 ;
        RECT 184.930 2349.490 186.110 2350.670 ;
        RECT 184.930 2171.090 186.110 2172.270 ;
        RECT 184.930 2169.490 186.110 2170.670 ;
        RECT 184.930 1991.090 186.110 1992.270 ;
        RECT 184.930 1989.490 186.110 1990.670 ;
        RECT 184.930 1811.090 186.110 1812.270 ;
        RECT 184.930 1809.490 186.110 1810.670 ;
        RECT 184.930 1631.090 186.110 1632.270 ;
        RECT 184.930 1629.490 186.110 1630.670 ;
        RECT 184.930 1451.090 186.110 1452.270 ;
        RECT 184.930 1449.490 186.110 1450.670 ;
        RECT 184.930 1271.090 186.110 1272.270 ;
        RECT 184.930 1269.490 186.110 1270.670 ;
        RECT 184.930 1091.090 186.110 1092.270 ;
        RECT 184.930 1089.490 186.110 1090.670 ;
        RECT 184.930 911.090 186.110 912.270 ;
        RECT 184.930 909.490 186.110 910.670 ;
        RECT 184.930 731.090 186.110 732.270 ;
        RECT 184.930 729.490 186.110 730.670 ;
        RECT 184.930 551.090 186.110 552.270 ;
        RECT 184.930 549.490 186.110 550.670 ;
        RECT 184.930 371.090 186.110 372.270 ;
        RECT 184.930 369.490 186.110 370.670 ;
        RECT 184.930 191.090 186.110 192.270 ;
        RECT 184.930 189.490 186.110 190.670 ;
        RECT 184.930 11.090 186.110 12.270 ;
        RECT 184.930 9.490 186.110 10.670 ;
        RECT 184.930 -2.910 186.110 -1.730 ;
        RECT 184.930 -4.510 186.110 -3.330 ;
        RECT 364.930 3523.010 366.110 3524.190 ;
        RECT 364.930 3521.410 366.110 3522.590 ;
        RECT 364.930 3431.090 366.110 3432.270 ;
        RECT 364.930 3429.490 366.110 3430.670 ;
        RECT 364.930 3251.090 366.110 3252.270 ;
        RECT 364.930 3249.490 366.110 3250.670 ;
        RECT 364.930 3071.090 366.110 3072.270 ;
        RECT 364.930 3069.490 366.110 3070.670 ;
        RECT 364.930 2891.090 366.110 2892.270 ;
        RECT 364.930 2889.490 366.110 2890.670 ;
        RECT 364.930 2711.090 366.110 2712.270 ;
        RECT 364.930 2709.490 366.110 2710.670 ;
        RECT 364.930 2531.090 366.110 2532.270 ;
        RECT 364.930 2529.490 366.110 2530.670 ;
        RECT 364.930 2351.090 366.110 2352.270 ;
        RECT 364.930 2349.490 366.110 2350.670 ;
        RECT 364.930 2171.090 366.110 2172.270 ;
        RECT 364.930 2169.490 366.110 2170.670 ;
        RECT 364.930 1991.090 366.110 1992.270 ;
        RECT 364.930 1989.490 366.110 1990.670 ;
        RECT 364.930 1811.090 366.110 1812.270 ;
        RECT 364.930 1809.490 366.110 1810.670 ;
        RECT 364.930 1631.090 366.110 1632.270 ;
        RECT 364.930 1629.490 366.110 1630.670 ;
        RECT 364.930 1451.090 366.110 1452.270 ;
        RECT 364.930 1449.490 366.110 1450.670 ;
        RECT 364.930 1271.090 366.110 1272.270 ;
        RECT 364.930 1269.490 366.110 1270.670 ;
        RECT 364.930 1091.090 366.110 1092.270 ;
        RECT 364.930 1089.490 366.110 1090.670 ;
        RECT 364.930 911.090 366.110 912.270 ;
        RECT 364.930 909.490 366.110 910.670 ;
        RECT 364.930 731.090 366.110 732.270 ;
        RECT 364.930 729.490 366.110 730.670 ;
        RECT 364.930 551.090 366.110 552.270 ;
        RECT 364.930 549.490 366.110 550.670 ;
        RECT 364.930 371.090 366.110 372.270 ;
        RECT 364.930 369.490 366.110 370.670 ;
        RECT 364.930 191.090 366.110 192.270 ;
        RECT 364.930 189.490 366.110 190.670 ;
        RECT 364.930 11.090 366.110 12.270 ;
        RECT 364.930 9.490 366.110 10.670 ;
        RECT 364.930 -2.910 366.110 -1.730 ;
        RECT 364.930 -4.510 366.110 -3.330 ;
        RECT 544.930 3523.010 546.110 3524.190 ;
        RECT 544.930 3521.410 546.110 3522.590 ;
        RECT 544.930 3431.090 546.110 3432.270 ;
        RECT 544.930 3429.490 546.110 3430.670 ;
        RECT 544.930 3251.090 546.110 3252.270 ;
        RECT 544.930 3249.490 546.110 3250.670 ;
        RECT 544.930 3071.090 546.110 3072.270 ;
        RECT 544.930 3069.490 546.110 3070.670 ;
        RECT 544.930 2891.090 546.110 2892.270 ;
        RECT 544.930 2889.490 546.110 2890.670 ;
        RECT 544.930 2711.090 546.110 2712.270 ;
        RECT 544.930 2709.490 546.110 2710.670 ;
        RECT 544.930 2531.090 546.110 2532.270 ;
        RECT 544.930 2529.490 546.110 2530.670 ;
        RECT 544.930 2351.090 546.110 2352.270 ;
        RECT 544.930 2349.490 546.110 2350.670 ;
        RECT 544.930 2171.090 546.110 2172.270 ;
        RECT 544.930 2169.490 546.110 2170.670 ;
        RECT 544.930 1991.090 546.110 1992.270 ;
        RECT 544.930 1989.490 546.110 1990.670 ;
        RECT 544.930 1811.090 546.110 1812.270 ;
        RECT 544.930 1809.490 546.110 1810.670 ;
        RECT 544.930 1631.090 546.110 1632.270 ;
        RECT 544.930 1629.490 546.110 1630.670 ;
        RECT 544.930 1451.090 546.110 1452.270 ;
        RECT 544.930 1449.490 546.110 1450.670 ;
        RECT 544.930 1271.090 546.110 1272.270 ;
        RECT 544.930 1269.490 546.110 1270.670 ;
        RECT 544.930 1091.090 546.110 1092.270 ;
        RECT 544.930 1089.490 546.110 1090.670 ;
        RECT 544.930 911.090 546.110 912.270 ;
        RECT 544.930 909.490 546.110 910.670 ;
        RECT 544.930 731.090 546.110 732.270 ;
        RECT 544.930 729.490 546.110 730.670 ;
        RECT 544.930 551.090 546.110 552.270 ;
        RECT 544.930 549.490 546.110 550.670 ;
        RECT 544.930 371.090 546.110 372.270 ;
        RECT 544.930 369.490 546.110 370.670 ;
        RECT 544.930 191.090 546.110 192.270 ;
        RECT 544.930 189.490 546.110 190.670 ;
        RECT 544.930 11.090 546.110 12.270 ;
        RECT 544.930 9.490 546.110 10.670 ;
        RECT 544.930 -2.910 546.110 -1.730 ;
        RECT 544.930 -4.510 546.110 -3.330 ;
        RECT 724.930 3523.010 726.110 3524.190 ;
        RECT 724.930 3521.410 726.110 3522.590 ;
        RECT 724.930 3431.090 726.110 3432.270 ;
        RECT 724.930 3429.490 726.110 3430.670 ;
        RECT 724.930 3251.090 726.110 3252.270 ;
        RECT 724.930 3249.490 726.110 3250.670 ;
        RECT 724.930 3071.090 726.110 3072.270 ;
        RECT 724.930 3069.490 726.110 3070.670 ;
        RECT 724.930 2891.090 726.110 2892.270 ;
        RECT 724.930 2889.490 726.110 2890.670 ;
        RECT 724.930 2711.090 726.110 2712.270 ;
        RECT 724.930 2709.490 726.110 2710.670 ;
        RECT 724.930 2531.090 726.110 2532.270 ;
        RECT 724.930 2529.490 726.110 2530.670 ;
        RECT 724.930 2351.090 726.110 2352.270 ;
        RECT 724.930 2349.490 726.110 2350.670 ;
        RECT 724.930 2171.090 726.110 2172.270 ;
        RECT 724.930 2169.490 726.110 2170.670 ;
        RECT 724.930 1991.090 726.110 1992.270 ;
        RECT 724.930 1989.490 726.110 1990.670 ;
        RECT 724.930 1811.090 726.110 1812.270 ;
        RECT 724.930 1809.490 726.110 1810.670 ;
        RECT 724.930 1631.090 726.110 1632.270 ;
        RECT 724.930 1629.490 726.110 1630.670 ;
        RECT 724.930 1451.090 726.110 1452.270 ;
        RECT 724.930 1449.490 726.110 1450.670 ;
        RECT 724.930 1271.090 726.110 1272.270 ;
        RECT 724.930 1269.490 726.110 1270.670 ;
        RECT 724.930 1091.090 726.110 1092.270 ;
        RECT 724.930 1089.490 726.110 1090.670 ;
        RECT 724.930 911.090 726.110 912.270 ;
        RECT 724.930 909.490 726.110 910.670 ;
        RECT 724.930 731.090 726.110 732.270 ;
        RECT 724.930 729.490 726.110 730.670 ;
        RECT 724.930 551.090 726.110 552.270 ;
        RECT 724.930 549.490 726.110 550.670 ;
        RECT 724.930 371.090 726.110 372.270 ;
        RECT 724.930 369.490 726.110 370.670 ;
        RECT 724.930 191.090 726.110 192.270 ;
        RECT 724.930 189.490 726.110 190.670 ;
        RECT 724.930 11.090 726.110 12.270 ;
        RECT 724.930 9.490 726.110 10.670 ;
        RECT 724.930 -2.910 726.110 -1.730 ;
        RECT 724.930 -4.510 726.110 -3.330 ;
        RECT 904.930 3523.010 906.110 3524.190 ;
        RECT 904.930 3521.410 906.110 3522.590 ;
        RECT 904.930 3431.090 906.110 3432.270 ;
        RECT 904.930 3429.490 906.110 3430.670 ;
        RECT 904.930 3251.090 906.110 3252.270 ;
        RECT 904.930 3249.490 906.110 3250.670 ;
        RECT 904.930 3071.090 906.110 3072.270 ;
        RECT 904.930 3069.490 906.110 3070.670 ;
        RECT 904.930 2891.090 906.110 2892.270 ;
        RECT 904.930 2889.490 906.110 2890.670 ;
        RECT 904.930 2711.090 906.110 2712.270 ;
        RECT 904.930 2709.490 906.110 2710.670 ;
        RECT 904.930 2531.090 906.110 2532.270 ;
        RECT 904.930 2529.490 906.110 2530.670 ;
        RECT 904.930 2351.090 906.110 2352.270 ;
        RECT 904.930 2349.490 906.110 2350.670 ;
        RECT 904.930 2171.090 906.110 2172.270 ;
        RECT 904.930 2169.490 906.110 2170.670 ;
        RECT 904.930 1991.090 906.110 1992.270 ;
        RECT 904.930 1989.490 906.110 1990.670 ;
        RECT 904.930 1811.090 906.110 1812.270 ;
        RECT 904.930 1809.490 906.110 1810.670 ;
        RECT 904.930 1631.090 906.110 1632.270 ;
        RECT 904.930 1629.490 906.110 1630.670 ;
        RECT 904.930 1451.090 906.110 1452.270 ;
        RECT 904.930 1449.490 906.110 1450.670 ;
        RECT 904.930 1271.090 906.110 1272.270 ;
        RECT 904.930 1269.490 906.110 1270.670 ;
        RECT 904.930 1091.090 906.110 1092.270 ;
        RECT 904.930 1089.490 906.110 1090.670 ;
        RECT 904.930 911.090 906.110 912.270 ;
        RECT 904.930 909.490 906.110 910.670 ;
        RECT 904.930 731.090 906.110 732.270 ;
        RECT 904.930 729.490 906.110 730.670 ;
        RECT 904.930 551.090 906.110 552.270 ;
        RECT 904.930 549.490 906.110 550.670 ;
        RECT 904.930 371.090 906.110 372.270 ;
        RECT 904.930 369.490 906.110 370.670 ;
        RECT 904.930 191.090 906.110 192.270 ;
        RECT 904.930 189.490 906.110 190.670 ;
        RECT 904.930 11.090 906.110 12.270 ;
        RECT 904.930 9.490 906.110 10.670 ;
        RECT 904.930 -2.910 906.110 -1.730 ;
        RECT 904.930 -4.510 906.110 -3.330 ;
        RECT 1084.930 3523.010 1086.110 3524.190 ;
        RECT 1084.930 3521.410 1086.110 3522.590 ;
        RECT 1084.930 3431.090 1086.110 3432.270 ;
        RECT 1084.930 3429.490 1086.110 3430.670 ;
        RECT 1084.930 3251.090 1086.110 3252.270 ;
        RECT 1084.930 3249.490 1086.110 3250.670 ;
        RECT 1084.930 3071.090 1086.110 3072.270 ;
        RECT 1084.930 3069.490 1086.110 3070.670 ;
        RECT 1084.930 2891.090 1086.110 2892.270 ;
        RECT 1084.930 2889.490 1086.110 2890.670 ;
        RECT 1084.930 2711.090 1086.110 2712.270 ;
        RECT 1084.930 2709.490 1086.110 2710.670 ;
        RECT 1084.930 2531.090 1086.110 2532.270 ;
        RECT 1084.930 2529.490 1086.110 2530.670 ;
        RECT 1084.930 2351.090 1086.110 2352.270 ;
        RECT 1084.930 2349.490 1086.110 2350.670 ;
        RECT 1084.930 2171.090 1086.110 2172.270 ;
        RECT 1084.930 2169.490 1086.110 2170.670 ;
        RECT 1084.930 1991.090 1086.110 1992.270 ;
        RECT 1084.930 1989.490 1086.110 1990.670 ;
        RECT 1084.930 1811.090 1086.110 1812.270 ;
        RECT 1084.930 1809.490 1086.110 1810.670 ;
        RECT 1084.930 1631.090 1086.110 1632.270 ;
        RECT 1084.930 1629.490 1086.110 1630.670 ;
        RECT 1084.930 1451.090 1086.110 1452.270 ;
        RECT 1084.930 1449.490 1086.110 1450.670 ;
        RECT 1084.930 1271.090 1086.110 1272.270 ;
        RECT 1084.930 1269.490 1086.110 1270.670 ;
        RECT 1084.930 1091.090 1086.110 1092.270 ;
        RECT 1084.930 1089.490 1086.110 1090.670 ;
        RECT 1084.930 911.090 1086.110 912.270 ;
        RECT 1084.930 909.490 1086.110 910.670 ;
        RECT 1084.930 731.090 1086.110 732.270 ;
        RECT 1084.930 729.490 1086.110 730.670 ;
        RECT 1084.930 551.090 1086.110 552.270 ;
        RECT 1084.930 549.490 1086.110 550.670 ;
        RECT 1084.930 371.090 1086.110 372.270 ;
        RECT 1084.930 369.490 1086.110 370.670 ;
        RECT 1084.930 191.090 1086.110 192.270 ;
        RECT 1084.930 189.490 1086.110 190.670 ;
        RECT 1084.930 11.090 1086.110 12.270 ;
        RECT 1084.930 9.490 1086.110 10.670 ;
        RECT 1084.930 -2.910 1086.110 -1.730 ;
        RECT 1084.930 -4.510 1086.110 -3.330 ;
        RECT 1264.930 3523.010 1266.110 3524.190 ;
        RECT 1264.930 3521.410 1266.110 3522.590 ;
        RECT 1264.930 3431.090 1266.110 3432.270 ;
        RECT 1264.930 3429.490 1266.110 3430.670 ;
        RECT 1264.930 3251.090 1266.110 3252.270 ;
        RECT 1264.930 3249.490 1266.110 3250.670 ;
        RECT 1264.930 3071.090 1266.110 3072.270 ;
        RECT 1264.930 3069.490 1266.110 3070.670 ;
        RECT 1264.930 2891.090 1266.110 2892.270 ;
        RECT 1264.930 2889.490 1266.110 2890.670 ;
        RECT 1264.930 2711.090 1266.110 2712.270 ;
        RECT 1264.930 2709.490 1266.110 2710.670 ;
        RECT 1264.930 2531.090 1266.110 2532.270 ;
        RECT 1264.930 2529.490 1266.110 2530.670 ;
        RECT 1264.930 2351.090 1266.110 2352.270 ;
        RECT 1264.930 2349.490 1266.110 2350.670 ;
        RECT 1264.930 2171.090 1266.110 2172.270 ;
        RECT 1264.930 2169.490 1266.110 2170.670 ;
        RECT 1264.930 1991.090 1266.110 1992.270 ;
        RECT 1264.930 1989.490 1266.110 1990.670 ;
        RECT 1264.930 1811.090 1266.110 1812.270 ;
        RECT 1264.930 1809.490 1266.110 1810.670 ;
        RECT 1264.930 1631.090 1266.110 1632.270 ;
        RECT 1264.930 1629.490 1266.110 1630.670 ;
        RECT 1264.930 1451.090 1266.110 1452.270 ;
        RECT 1264.930 1449.490 1266.110 1450.670 ;
        RECT 1264.930 1271.090 1266.110 1272.270 ;
        RECT 1264.930 1269.490 1266.110 1270.670 ;
        RECT 1264.930 1091.090 1266.110 1092.270 ;
        RECT 1264.930 1089.490 1266.110 1090.670 ;
        RECT 1264.930 911.090 1266.110 912.270 ;
        RECT 1264.930 909.490 1266.110 910.670 ;
        RECT 1264.930 731.090 1266.110 732.270 ;
        RECT 1264.930 729.490 1266.110 730.670 ;
        RECT 1264.930 551.090 1266.110 552.270 ;
        RECT 1264.930 549.490 1266.110 550.670 ;
        RECT 1264.930 371.090 1266.110 372.270 ;
        RECT 1264.930 369.490 1266.110 370.670 ;
        RECT 1264.930 191.090 1266.110 192.270 ;
        RECT 1264.930 189.490 1266.110 190.670 ;
        RECT 1264.930 11.090 1266.110 12.270 ;
        RECT 1264.930 9.490 1266.110 10.670 ;
        RECT 1264.930 -2.910 1266.110 -1.730 ;
        RECT 1264.930 -4.510 1266.110 -3.330 ;
        RECT 1444.930 3523.010 1446.110 3524.190 ;
        RECT 1444.930 3521.410 1446.110 3522.590 ;
        RECT 1444.930 3431.090 1446.110 3432.270 ;
        RECT 1444.930 3429.490 1446.110 3430.670 ;
        RECT 1444.930 3251.090 1446.110 3252.270 ;
        RECT 1444.930 3249.490 1446.110 3250.670 ;
        RECT 1444.930 3071.090 1446.110 3072.270 ;
        RECT 1444.930 3069.490 1446.110 3070.670 ;
        RECT 1444.930 2891.090 1446.110 2892.270 ;
        RECT 1444.930 2889.490 1446.110 2890.670 ;
        RECT 1444.930 2711.090 1446.110 2712.270 ;
        RECT 1444.930 2709.490 1446.110 2710.670 ;
        RECT 1444.930 2531.090 1446.110 2532.270 ;
        RECT 1444.930 2529.490 1446.110 2530.670 ;
        RECT 1444.930 2351.090 1446.110 2352.270 ;
        RECT 1444.930 2349.490 1446.110 2350.670 ;
        RECT 1444.930 2171.090 1446.110 2172.270 ;
        RECT 1444.930 2169.490 1446.110 2170.670 ;
        RECT 1444.930 1991.090 1446.110 1992.270 ;
        RECT 1444.930 1989.490 1446.110 1990.670 ;
        RECT 1444.930 1811.090 1446.110 1812.270 ;
        RECT 1444.930 1809.490 1446.110 1810.670 ;
        RECT 1444.930 1631.090 1446.110 1632.270 ;
        RECT 1444.930 1629.490 1446.110 1630.670 ;
        RECT 1444.930 1451.090 1446.110 1452.270 ;
        RECT 1444.930 1449.490 1446.110 1450.670 ;
        RECT 1444.930 1271.090 1446.110 1272.270 ;
        RECT 1444.930 1269.490 1446.110 1270.670 ;
        RECT 1444.930 1091.090 1446.110 1092.270 ;
        RECT 1444.930 1089.490 1446.110 1090.670 ;
        RECT 1444.930 911.090 1446.110 912.270 ;
        RECT 1444.930 909.490 1446.110 910.670 ;
        RECT 1444.930 731.090 1446.110 732.270 ;
        RECT 1444.930 729.490 1446.110 730.670 ;
        RECT 1444.930 551.090 1446.110 552.270 ;
        RECT 1444.930 549.490 1446.110 550.670 ;
        RECT 1444.930 371.090 1446.110 372.270 ;
        RECT 1444.930 369.490 1446.110 370.670 ;
        RECT 1444.930 191.090 1446.110 192.270 ;
        RECT 1444.930 189.490 1446.110 190.670 ;
        RECT 1444.930 11.090 1446.110 12.270 ;
        RECT 1444.930 9.490 1446.110 10.670 ;
        RECT 1444.930 -2.910 1446.110 -1.730 ;
        RECT 1444.930 -4.510 1446.110 -3.330 ;
        RECT 1624.930 3523.010 1626.110 3524.190 ;
        RECT 1624.930 3521.410 1626.110 3522.590 ;
        RECT 1624.930 3431.090 1626.110 3432.270 ;
        RECT 1624.930 3429.490 1626.110 3430.670 ;
        RECT 1624.930 3251.090 1626.110 3252.270 ;
        RECT 1624.930 3249.490 1626.110 3250.670 ;
        RECT 1624.930 3071.090 1626.110 3072.270 ;
        RECT 1624.930 3069.490 1626.110 3070.670 ;
        RECT 1624.930 2891.090 1626.110 2892.270 ;
        RECT 1624.930 2889.490 1626.110 2890.670 ;
        RECT 1624.930 2711.090 1626.110 2712.270 ;
        RECT 1624.930 2709.490 1626.110 2710.670 ;
        RECT 1624.930 2531.090 1626.110 2532.270 ;
        RECT 1624.930 2529.490 1626.110 2530.670 ;
        RECT 1624.930 2351.090 1626.110 2352.270 ;
        RECT 1624.930 2349.490 1626.110 2350.670 ;
        RECT 1624.930 2171.090 1626.110 2172.270 ;
        RECT 1624.930 2169.490 1626.110 2170.670 ;
        RECT 1624.930 1991.090 1626.110 1992.270 ;
        RECT 1624.930 1989.490 1626.110 1990.670 ;
        RECT 1624.930 1811.090 1626.110 1812.270 ;
        RECT 1624.930 1809.490 1626.110 1810.670 ;
        RECT 1624.930 1631.090 1626.110 1632.270 ;
        RECT 1624.930 1629.490 1626.110 1630.670 ;
        RECT 1624.930 1451.090 1626.110 1452.270 ;
        RECT 1624.930 1449.490 1626.110 1450.670 ;
        RECT 1624.930 1271.090 1626.110 1272.270 ;
        RECT 1624.930 1269.490 1626.110 1270.670 ;
        RECT 1624.930 1091.090 1626.110 1092.270 ;
        RECT 1624.930 1089.490 1626.110 1090.670 ;
        RECT 1624.930 911.090 1626.110 912.270 ;
        RECT 1624.930 909.490 1626.110 910.670 ;
        RECT 1624.930 731.090 1626.110 732.270 ;
        RECT 1624.930 729.490 1626.110 730.670 ;
        RECT 1624.930 551.090 1626.110 552.270 ;
        RECT 1624.930 549.490 1626.110 550.670 ;
        RECT 1624.930 371.090 1626.110 372.270 ;
        RECT 1624.930 369.490 1626.110 370.670 ;
        RECT 1624.930 191.090 1626.110 192.270 ;
        RECT 1624.930 189.490 1626.110 190.670 ;
        RECT 1624.930 11.090 1626.110 12.270 ;
        RECT 1624.930 9.490 1626.110 10.670 ;
        RECT 1624.930 -2.910 1626.110 -1.730 ;
        RECT 1624.930 -4.510 1626.110 -3.330 ;
        RECT 1804.930 3523.010 1806.110 3524.190 ;
        RECT 1804.930 3521.410 1806.110 3522.590 ;
        RECT 1804.930 3431.090 1806.110 3432.270 ;
        RECT 1804.930 3429.490 1806.110 3430.670 ;
        RECT 1804.930 3251.090 1806.110 3252.270 ;
        RECT 1804.930 3249.490 1806.110 3250.670 ;
        RECT 1804.930 3071.090 1806.110 3072.270 ;
        RECT 1804.930 3069.490 1806.110 3070.670 ;
        RECT 1804.930 2891.090 1806.110 2892.270 ;
        RECT 1804.930 2889.490 1806.110 2890.670 ;
        RECT 1804.930 2711.090 1806.110 2712.270 ;
        RECT 1804.930 2709.490 1806.110 2710.670 ;
        RECT 1804.930 2531.090 1806.110 2532.270 ;
        RECT 1804.930 2529.490 1806.110 2530.670 ;
        RECT 1804.930 2351.090 1806.110 2352.270 ;
        RECT 1804.930 2349.490 1806.110 2350.670 ;
        RECT 1804.930 2171.090 1806.110 2172.270 ;
        RECT 1804.930 2169.490 1806.110 2170.670 ;
        RECT 1804.930 1991.090 1806.110 1992.270 ;
        RECT 1804.930 1989.490 1806.110 1990.670 ;
        RECT 1804.930 1811.090 1806.110 1812.270 ;
        RECT 1804.930 1809.490 1806.110 1810.670 ;
        RECT 1804.930 1631.090 1806.110 1632.270 ;
        RECT 1804.930 1629.490 1806.110 1630.670 ;
        RECT 1804.930 1451.090 1806.110 1452.270 ;
        RECT 1804.930 1449.490 1806.110 1450.670 ;
        RECT 1804.930 1271.090 1806.110 1272.270 ;
        RECT 1804.930 1269.490 1806.110 1270.670 ;
        RECT 1804.930 1091.090 1806.110 1092.270 ;
        RECT 1804.930 1089.490 1806.110 1090.670 ;
        RECT 1804.930 911.090 1806.110 912.270 ;
        RECT 1804.930 909.490 1806.110 910.670 ;
        RECT 1804.930 731.090 1806.110 732.270 ;
        RECT 1804.930 729.490 1806.110 730.670 ;
        RECT 1804.930 551.090 1806.110 552.270 ;
        RECT 1804.930 549.490 1806.110 550.670 ;
        RECT 1804.930 371.090 1806.110 372.270 ;
        RECT 1804.930 369.490 1806.110 370.670 ;
        RECT 1804.930 191.090 1806.110 192.270 ;
        RECT 1804.930 189.490 1806.110 190.670 ;
        RECT 1804.930 11.090 1806.110 12.270 ;
        RECT 1804.930 9.490 1806.110 10.670 ;
        RECT 1804.930 -2.910 1806.110 -1.730 ;
        RECT 1804.930 -4.510 1806.110 -3.330 ;
        RECT 1984.930 3523.010 1986.110 3524.190 ;
        RECT 1984.930 3521.410 1986.110 3522.590 ;
        RECT 1984.930 3431.090 1986.110 3432.270 ;
        RECT 1984.930 3429.490 1986.110 3430.670 ;
        RECT 1984.930 3251.090 1986.110 3252.270 ;
        RECT 1984.930 3249.490 1986.110 3250.670 ;
        RECT 1984.930 3071.090 1986.110 3072.270 ;
        RECT 1984.930 3069.490 1986.110 3070.670 ;
        RECT 1984.930 2891.090 1986.110 2892.270 ;
        RECT 1984.930 2889.490 1986.110 2890.670 ;
        RECT 1984.930 2711.090 1986.110 2712.270 ;
        RECT 1984.930 2709.490 1986.110 2710.670 ;
        RECT 1984.930 2531.090 1986.110 2532.270 ;
        RECT 1984.930 2529.490 1986.110 2530.670 ;
        RECT 1984.930 2351.090 1986.110 2352.270 ;
        RECT 1984.930 2349.490 1986.110 2350.670 ;
        RECT 1984.930 2171.090 1986.110 2172.270 ;
        RECT 1984.930 2169.490 1986.110 2170.670 ;
        RECT 1984.930 1991.090 1986.110 1992.270 ;
        RECT 1984.930 1989.490 1986.110 1990.670 ;
        RECT 1984.930 1811.090 1986.110 1812.270 ;
        RECT 1984.930 1809.490 1986.110 1810.670 ;
        RECT 1984.930 1631.090 1986.110 1632.270 ;
        RECT 1984.930 1629.490 1986.110 1630.670 ;
        RECT 1984.930 1451.090 1986.110 1452.270 ;
        RECT 1984.930 1449.490 1986.110 1450.670 ;
        RECT 1984.930 1271.090 1986.110 1272.270 ;
        RECT 1984.930 1269.490 1986.110 1270.670 ;
        RECT 1984.930 1091.090 1986.110 1092.270 ;
        RECT 1984.930 1089.490 1986.110 1090.670 ;
        RECT 1984.930 911.090 1986.110 912.270 ;
        RECT 1984.930 909.490 1986.110 910.670 ;
        RECT 1984.930 731.090 1986.110 732.270 ;
        RECT 1984.930 729.490 1986.110 730.670 ;
        RECT 1984.930 551.090 1986.110 552.270 ;
        RECT 1984.930 549.490 1986.110 550.670 ;
        RECT 1984.930 371.090 1986.110 372.270 ;
        RECT 1984.930 369.490 1986.110 370.670 ;
        RECT 1984.930 191.090 1986.110 192.270 ;
        RECT 1984.930 189.490 1986.110 190.670 ;
        RECT 1984.930 11.090 1986.110 12.270 ;
        RECT 1984.930 9.490 1986.110 10.670 ;
        RECT 1984.930 -2.910 1986.110 -1.730 ;
        RECT 1984.930 -4.510 1986.110 -3.330 ;
        RECT 2164.930 3523.010 2166.110 3524.190 ;
        RECT 2164.930 3521.410 2166.110 3522.590 ;
        RECT 2164.930 3431.090 2166.110 3432.270 ;
        RECT 2164.930 3429.490 2166.110 3430.670 ;
        RECT 2164.930 3251.090 2166.110 3252.270 ;
        RECT 2164.930 3249.490 2166.110 3250.670 ;
        RECT 2164.930 3071.090 2166.110 3072.270 ;
        RECT 2164.930 3069.490 2166.110 3070.670 ;
        RECT 2164.930 2891.090 2166.110 2892.270 ;
        RECT 2164.930 2889.490 2166.110 2890.670 ;
        RECT 2164.930 2711.090 2166.110 2712.270 ;
        RECT 2164.930 2709.490 2166.110 2710.670 ;
        RECT 2164.930 2531.090 2166.110 2532.270 ;
        RECT 2164.930 2529.490 2166.110 2530.670 ;
        RECT 2164.930 2351.090 2166.110 2352.270 ;
        RECT 2164.930 2349.490 2166.110 2350.670 ;
        RECT 2164.930 2171.090 2166.110 2172.270 ;
        RECT 2164.930 2169.490 2166.110 2170.670 ;
        RECT 2164.930 1991.090 2166.110 1992.270 ;
        RECT 2164.930 1989.490 2166.110 1990.670 ;
        RECT 2164.930 1811.090 2166.110 1812.270 ;
        RECT 2164.930 1809.490 2166.110 1810.670 ;
        RECT 2164.930 1631.090 2166.110 1632.270 ;
        RECT 2164.930 1629.490 2166.110 1630.670 ;
        RECT 2164.930 1451.090 2166.110 1452.270 ;
        RECT 2164.930 1449.490 2166.110 1450.670 ;
        RECT 2164.930 1271.090 2166.110 1272.270 ;
        RECT 2164.930 1269.490 2166.110 1270.670 ;
        RECT 2164.930 1091.090 2166.110 1092.270 ;
        RECT 2164.930 1089.490 2166.110 1090.670 ;
        RECT 2164.930 911.090 2166.110 912.270 ;
        RECT 2164.930 909.490 2166.110 910.670 ;
        RECT 2164.930 731.090 2166.110 732.270 ;
        RECT 2164.930 729.490 2166.110 730.670 ;
        RECT 2164.930 551.090 2166.110 552.270 ;
        RECT 2164.930 549.490 2166.110 550.670 ;
        RECT 2164.930 371.090 2166.110 372.270 ;
        RECT 2164.930 369.490 2166.110 370.670 ;
        RECT 2164.930 191.090 2166.110 192.270 ;
        RECT 2164.930 189.490 2166.110 190.670 ;
        RECT 2164.930 11.090 2166.110 12.270 ;
        RECT 2164.930 9.490 2166.110 10.670 ;
        RECT 2164.930 -2.910 2166.110 -1.730 ;
        RECT 2164.930 -4.510 2166.110 -3.330 ;
        RECT 2344.930 3523.010 2346.110 3524.190 ;
        RECT 2344.930 3521.410 2346.110 3522.590 ;
        RECT 2344.930 3431.090 2346.110 3432.270 ;
        RECT 2344.930 3429.490 2346.110 3430.670 ;
        RECT 2344.930 3251.090 2346.110 3252.270 ;
        RECT 2344.930 3249.490 2346.110 3250.670 ;
        RECT 2344.930 3071.090 2346.110 3072.270 ;
        RECT 2344.930 3069.490 2346.110 3070.670 ;
        RECT 2344.930 2891.090 2346.110 2892.270 ;
        RECT 2344.930 2889.490 2346.110 2890.670 ;
        RECT 2344.930 2711.090 2346.110 2712.270 ;
        RECT 2344.930 2709.490 2346.110 2710.670 ;
        RECT 2344.930 2531.090 2346.110 2532.270 ;
        RECT 2344.930 2529.490 2346.110 2530.670 ;
        RECT 2344.930 2351.090 2346.110 2352.270 ;
        RECT 2344.930 2349.490 2346.110 2350.670 ;
        RECT 2344.930 2171.090 2346.110 2172.270 ;
        RECT 2344.930 2169.490 2346.110 2170.670 ;
        RECT 2344.930 1991.090 2346.110 1992.270 ;
        RECT 2344.930 1989.490 2346.110 1990.670 ;
        RECT 2344.930 1811.090 2346.110 1812.270 ;
        RECT 2344.930 1809.490 2346.110 1810.670 ;
        RECT 2344.930 1631.090 2346.110 1632.270 ;
        RECT 2344.930 1629.490 2346.110 1630.670 ;
        RECT 2344.930 1451.090 2346.110 1452.270 ;
        RECT 2344.930 1449.490 2346.110 1450.670 ;
        RECT 2344.930 1271.090 2346.110 1272.270 ;
        RECT 2344.930 1269.490 2346.110 1270.670 ;
        RECT 2344.930 1091.090 2346.110 1092.270 ;
        RECT 2344.930 1089.490 2346.110 1090.670 ;
        RECT 2344.930 911.090 2346.110 912.270 ;
        RECT 2344.930 909.490 2346.110 910.670 ;
        RECT 2344.930 731.090 2346.110 732.270 ;
        RECT 2344.930 729.490 2346.110 730.670 ;
        RECT 2344.930 551.090 2346.110 552.270 ;
        RECT 2344.930 549.490 2346.110 550.670 ;
        RECT 2344.930 371.090 2346.110 372.270 ;
        RECT 2344.930 369.490 2346.110 370.670 ;
        RECT 2344.930 191.090 2346.110 192.270 ;
        RECT 2344.930 189.490 2346.110 190.670 ;
        RECT 2344.930 11.090 2346.110 12.270 ;
        RECT 2344.930 9.490 2346.110 10.670 ;
        RECT 2344.930 -2.910 2346.110 -1.730 ;
        RECT 2344.930 -4.510 2346.110 -3.330 ;
        RECT 2524.930 3523.010 2526.110 3524.190 ;
        RECT 2524.930 3521.410 2526.110 3522.590 ;
        RECT 2524.930 3431.090 2526.110 3432.270 ;
        RECT 2524.930 3429.490 2526.110 3430.670 ;
        RECT 2524.930 3251.090 2526.110 3252.270 ;
        RECT 2524.930 3249.490 2526.110 3250.670 ;
        RECT 2524.930 3071.090 2526.110 3072.270 ;
        RECT 2524.930 3069.490 2526.110 3070.670 ;
        RECT 2524.930 2891.090 2526.110 2892.270 ;
        RECT 2524.930 2889.490 2526.110 2890.670 ;
        RECT 2524.930 2711.090 2526.110 2712.270 ;
        RECT 2524.930 2709.490 2526.110 2710.670 ;
        RECT 2524.930 2531.090 2526.110 2532.270 ;
        RECT 2524.930 2529.490 2526.110 2530.670 ;
        RECT 2524.930 2351.090 2526.110 2352.270 ;
        RECT 2524.930 2349.490 2526.110 2350.670 ;
        RECT 2524.930 2171.090 2526.110 2172.270 ;
        RECT 2524.930 2169.490 2526.110 2170.670 ;
        RECT 2524.930 1991.090 2526.110 1992.270 ;
        RECT 2524.930 1989.490 2526.110 1990.670 ;
        RECT 2524.930 1811.090 2526.110 1812.270 ;
        RECT 2524.930 1809.490 2526.110 1810.670 ;
        RECT 2524.930 1631.090 2526.110 1632.270 ;
        RECT 2524.930 1629.490 2526.110 1630.670 ;
        RECT 2524.930 1451.090 2526.110 1452.270 ;
        RECT 2524.930 1449.490 2526.110 1450.670 ;
        RECT 2524.930 1271.090 2526.110 1272.270 ;
        RECT 2524.930 1269.490 2526.110 1270.670 ;
        RECT 2524.930 1091.090 2526.110 1092.270 ;
        RECT 2524.930 1089.490 2526.110 1090.670 ;
        RECT 2524.930 911.090 2526.110 912.270 ;
        RECT 2524.930 909.490 2526.110 910.670 ;
        RECT 2524.930 731.090 2526.110 732.270 ;
        RECT 2524.930 729.490 2526.110 730.670 ;
        RECT 2524.930 551.090 2526.110 552.270 ;
        RECT 2524.930 549.490 2526.110 550.670 ;
        RECT 2524.930 371.090 2526.110 372.270 ;
        RECT 2524.930 369.490 2526.110 370.670 ;
        RECT 2524.930 191.090 2526.110 192.270 ;
        RECT 2524.930 189.490 2526.110 190.670 ;
        RECT 2524.930 11.090 2526.110 12.270 ;
        RECT 2524.930 9.490 2526.110 10.670 ;
        RECT 2524.930 -2.910 2526.110 -1.730 ;
        RECT 2524.930 -4.510 2526.110 -3.330 ;
        RECT 2704.930 3523.010 2706.110 3524.190 ;
        RECT 2704.930 3521.410 2706.110 3522.590 ;
        RECT 2704.930 3431.090 2706.110 3432.270 ;
        RECT 2704.930 3429.490 2706.110 3430.670 ;
        RECT 2704.930 3251.090 2706.110 3252.270 ;
        RECT 2704.930 3249.490 2706.110 3250.670 ;
        RECT 2704.930 3071.090 2706.110 3072.270 ;
        RECT 2704.930 3069.490 2706.110 3070.670 ;
        RECT 2704.930 2891.090 2706.110 2892.270 ;
        RECT 2704.930 2889.490 2706.110 2890.670 ;
        RECT 2704.930 2711.090 2706.110 2712.270 ;
        RECT 2704.930 2709.490 2706.110 2710.670 ;
        RECT 2704.930 2531.090 2706.110 2532.270 ;
        RECT 2704.930 2529.490 2706.110 2530.670 ;
        RECT 2704.930 2351.090 2706.110 2352.270 ;
        RECT 2704.930 2349.490 2706.110 2350.670 ;
        RECT 2704.930 2171.090 2706.110 2172.270 ;
        RECT 2704.930 2169.490 2706.110 2170.670 ;
        RECT 2704.930 1991.090 2706.110 1992.270 ;
        RECT 2704.930 1989.490 2706.110 1990.670 ;
        RECT 2704.930 1811.090 2706.110 1812.270 ;
        RECT 2704.930 1809.490 2706.110 1810.670 ;
        RECT 2704.930 1631.090 2706.110 1632.270 ;
        RECT 2704.930 1629.490 2706.110 1630.670 ;
        RECT 2704.930 1451.090 2706.110 1452.270 ;
        RECT 2704.930 1449.490 2706.110 1450.670 ;
        RECT 2704.930 1271.090 2706.110 1272.270 ;
        RECT 2704.930 1269.490 2706.110 1270.670 ;
        RECT 2704.930 1091.090 2706.110 1092.270 ;
        RECT 2704.930 1089.490 2706.110 1090.670 ;
        RECT 2704.930 911.090 2706.110 912.270 ;
        RECT 2704.930 909.490 2706.110 910.670 ;
        RECT 2704.930 731.090 2706.110 732.270 ;
        RECT 2704.930 729.490 2706.110 730.670 ;
        RECT 2704.930 551.090 2706.110 552.270 ;
        RECT 2704.930 549.490 2706.110 550.670 ;
        RECT 2704.930 371.090 2706.110 372.270 ;
        RECT 2704.930 369.490 2706.110 370.670 ;
        RECT 2704.930 191.090 2706.110 192.270 ;
        RECT 2704.930 189.490 2706.110 190.670 ;
        RECT 2704.930 11.090 2706.110 12.270 ;
        RECT 2704.930 9.490 2706.110 10.670 ;
        RECT 2704.930 -2.910 2706.110 -1.730 ;
        RECT 2704.930 -4.510 2706.110 -3.330 ;
        RECT 2884.930 3523.010 2886.110 3524.190 ;
        RECT 2884.930 3521.410 2886.110 3522.590 ;
        RECT 2884.930 3431.090 2886.110 3432.270 ;
        RECT 2884.930 3429.490 2886.110 3430.670 ;
        RECT 2884.930 3251.090 2886.110 3252.270 ;
        RECT 2884.930 3249.490 2886.110 3250.670 ;
        RECT 2884.930 3071.090 2886.110 3072.270 ;
        RECT 2884.930 3069.490 2886.110 3070.670 ;
        RECT 2884.930 2891.090 2886.110 2892.270 ;
        RECT 2884.930 2889.490 2886.110 2890.670 ;
        RECT 2884.930 2711.090 2886.110 2712.270 ;
        RECT 2884.930 2709.490 2886.110 2710.670 ;
        RECT 2884.930 2531.090 2886.110 2532.270 ;
        RECT 2884.930 2529.490 2886.110 2530.670 ;
        RECT 2884.930 2351.090 2886.110 2352.270 ;
        RECT 2884.930 2349.490 2886.110 2350.670 ;
        RECT 2884.930 2171.090 2886.110 2172.270 ;
        RECT 2884.930 2169.490 2886.110 2170.670 ;
        RECT 2884.930 1991.090 2886.110 1992.270 ;
        RECT 2884.930 1989.490 2886.110 1990.670 ;
        RECT 2884.930 1811.090 2886.110 1812.270 ;
        RECT 2884.930 1809.490 2886.110 1810.670 ;
        RECT 2884.930 1631.090 2886.110 1632.270 ;
        RECT 2884.930 1629.490 2886.110 1630.670 ;
        RECT 2884.930 1451.090 2886.110 1452.270 ;
        RECT 2884.930 1449.490 2886.110 1450.670 ;
        RECT 2884.930 1271.090 2886.110 1272.270 ;
        RECT 2884.930 1269.490 2886.110 1270.670 ;
        RECT 2884.930 1091.090 2886.110 1092.270 ;
        RECT 2884.930 1089.490 2886.110 1090.670 ;
        RECT 2884.930 911.090 2886.110 912.270 ;
        RECT 2884.930 909.490 2886.110 910.670 ;
        RECT 2884.930 731.090 2886.110 732.270 ;
        RECT 2884.930 729.490 2886.110 730.670 ;
        RECT 2884.930 551.090 2886.110 552.270 ;
        RECT 2884.930 549.490 2886.110 550.670 ;
        RECT 2884.930 371.090 2886.110 372.270 ;
        RECT 2884.930 369.490 2886.110 370.670 ;
        RECT 2884.930 191.090 2886.110 192.270 ;
        RECT 2884.930 189.490 2886.110 190.670 ;
        RECT 2884.930 11.090 2886.110 12.270 ;
        RECT 2884.930 9.490 2886.110 10.670 ;
        RECT 2884.930 -2.910 2886.110 -1.730 ;
        RECT 2884.930 -4.510 2886.110 -3.330 ;
        RECT 2927.510 3523.010 2928.690 3524.190 ;
        RECT 2927.510 3521.410 2928.690 3522.590 ;
        RECT 2927.510 3431.090 2928.690 3432.270 ;
        RECT 2927.510 3429.490 2928.690 3430.670 ;
        RECT 2927.510 3251.090 2928.690 3252.270 ;
        RECT 2927.510 3249.490 2928.690 3250.670 ;
        RECT 2927.510 3071.090 2928.690 3072.270 ;
        RECT 2927.510 3069.490 2928.690 3070.670 ;
        RECT 2927.510 2891.090 2928.690 2892.270 ;
        RECT 2927.510 2889.490 2928.690 2890.670 ;
        RECT 2927.510 2711.090 2928.690 2712.270 ;
        RECT 2927.510 2709.490 2928.690 2710.670 ;
        RECT 2927.510 2531.090 2928.690 2532.270 ;
        RECT 2927.510 2529.490 2928.690 2530.670 ;
        RECT 2927.510 2351.090 2928.690 2352.270 ;
        RECT 2927.510 2349.490 2928.690 2350.670 ;
        RECT 2927.510 2171.090 2928.690 2172.270 ;
        RECT 2927.510 2169.490 2928.690 2170.670 ;
        RECT 2927.510 1991.090 2928.690 1992.270 ;
        RECT 2927.510 1989.490 2928.690 1990.670 ;
        RECT 2927.510 1811.090 2928.690 1812.270 ;
        RECT 2927.510 1809.490 2928.690 1810.670 ;
        RECT 2927.510 1631.090 2928.690 1632.270 ;
        RECT 2927.510 1629.490 2928.690 1630.670 ;
        RECT 2927.510 1451.090 2928.690 1452.270 ;
        RECT 2927.510 1449.490 2928.690 1450.670 ;
        RECT 2927.510 1271.090 2928.690 1272.270 ;
        RECT 2927.510 1269.490 2928.690 1270.670 ;
        RECT 2927.510 1091.090 2928.690 1092.270 ;
        RECT 2927.510 1089.490 2928.690 1090.670 ;
        RECT 2927.510 911.090 2928.690 912.270 ;
        RECT 2927.510 909.490 2928.690 910.670 ;
        RECT 2927.510 731.090 2928.690 732.270 ;
        RECT 2927.510 729.490 2928.690 730.670 ;
        RECT 2927.510 551.090 2928.690 552.270 ;
        RECT 2927.510 549.490 2928.690 550.670 ;
        RECT 2927.510 371.090 2928.690 372.270 ;
        RECT 2927.510 369.490 2928.690 370.670 ;
        RECT 2927.510 191.090 2928.690 192.270 ;
        RECT 2927.510 189.490 2928.690 190.670 ;
        RECT 2927.510 11.090 2928.690 12.270 ;
        RECT 2927.510 9.490 2928.690 10.670 ;
        RECT 2927.510 -2.910 2928.690 -1.730 ;
        RECT 2927.510 -4.510 2928.690 -3.330 ;
      LAYER met5 ;
        RECT -9.980 3524.300 -6.980 3524.310 ;
        RECT 4.020 3524.300 7.020 3524.310 ;
        RECT 184.020 3524.300 187.020 3524.310 ;
        RECT 364.020 3524.300 367.020 3524.310 ;
        RECT 544.020 3524.300 547.020 3524.310 ;
        RECT 724.020 3524.300 727.020 3524.310 ;
        RECT 904.020 3524.300 907.020 3524.310 ;
        RECT 1084.020 3524.300 1087.020 3524.310 ;
        RECT 1264.020 3524.300 1267.020 3524.310 ;
        RECT 1444.020 3524.300 1447.020 3524.310 ;
        RECT 1624.020 3524.300 1627.020 3524.310 ;
        RECT 1804.020 3524.300 1807.020 3524.310 ;
        RECT 1984.020 3524.300 1987.020 3524.310 ;
        RECT 2164.020 3524.300 2167.020 3524.310 ;
        RECT 2344.020 3524.300 2347.020 3524.310 ;
        RECT 2524.020 3524.300 2527.020 3524.310 ;
        RECT 2704.020 3524.300 2707.020 3524.310 ;
        RECT 2884.020 3524.300 2887.020 3524.310 ;
        RECT 2926.600 3524.300 2929.600 3524.310 ;
        RECT -9.980 3521.300 2929.600 3524.300 ;
        RECT -9.980 3521.290 -6.980 3521.300 ;
        RECT 4.020 3521.290 7.020 3521.300 ;
        RECT 184.020 3521.290 187.020 3521.300 ;
        RECT 364.020 3521.290 367.020 3521.300 ;
        RECT 544.020 3521.290 547.020 3521.300 ;
        RECT 724.020 3521.290 727.020 3521.300 ;
        RECT 904.020 3521.290 907.020 3521.300 ;
        RECT 1084.020 3521.290 1087.020 3521.300 ;
        RECT 1264.020 3521.290 1267.020 3521.300 ;
        RECT 1444.020 3521.290 1447.020 3521.300 ;
        RECT 1624.020 3521.290 1627.020 3521.300 ;
        RECT 1804.020 3521.290 1807.020 3521.300 ;
        RECT 1984.020 3521.290 1987.020 3521.300 ;
        RECT 2164.020 3521.290 2167.020 3521.300 ;
        RECT 2344.020 3521.290 2347.020 3521.300 ;
        RECT 2524.020 3521.290 2527.020 3521.300 ;
        RECT 2704.020 3521.290 2707.020 3521.300 ;
        RECT 2884.020 3521.290 2887.020 3521.300 ;
        RECT 2926.600 3521.290 2929.600 3521.300 ;
        RECT -9.980 3432.380 -6.980 3432.390 ;
        RECT 4.020 3432.380 7.020 3432.390 ;
        RECT 184.020 3432.380 187.020 3432.390 ;
        RECT 364.020 3432.380 367.020 3432.390 ;
        RECT 544.020 3432.380 547.020 3432.390 ;
        RECT 724.020 3432.380 727.020 3432.390 ;
        RECT 904.020 3432.380 907.020 3432.390 ;
        RECT 1084.020 3432.380 1087.020 3432.390 ;
        RECT 1264.020 3432.380 1267.020 3432.390 ;
        RECT 1444.020 3432.380 1447.020 3432.390 ;
        RECT 1624.020 3432.380 1627.020 3432.390 ;
        RECT 1804.020 3432.380 1807.020 3432.390 ;
        RECT 1984.020 3432.380 1987.020 3432.390 ;
        RECT 2164.020 3432.380 2167.020 3432.390 ;
        RECT 2344.020 3432.380 2347.020 3432.390 ;
        RECT 2524.020 3432.380 2527.020 3432.390 ;
        RECT 2704.020 3432.380 2707.020 3432.390 ;
        RECT 2884.020 3432.380 2887.020 3432.390 ;
        RECT 2926.600 3432.380 2929.600 3432.390 ;
        RECT -14.580 3429.380 2934.200 3432.380 ;
        RECT -9.980 3429.370 -6.980 3429.380 ;
        RECT 4.020 3429.370 7.020 3429.380 ;
        RECT 184.020 3429.370 187.020 3429.380 ;
        RECT 364.020 3429.370 367.020 3429.380 ;
        RECT 544.020 3429.370 547.020 3429.380 ;
        RECT 724.020 3429.370 727.020 3429.380 ;
        RECT 904.020 3429.370 907.020 3429.380 ;
        RECT 1084.020 3429.370 1087.020 3429.380 ;
        RECT 1264.020 3429.370 1267.020 3429.380 ;
        RECT 1444.020 3429.370 1447.020 3429.380 ;
        RECT 1624.020 3429.370 1627.020 3429.380 ;
        RECT 1804.020 3429.370 1807.020 3429.380 ;
        RECT 1984.020 3429.370 1987.020 3429.380 ;
        RECT 2164.020 3429.370 2167.020 3429.380 ;
        RECT 2344.020 3429.370 2347.020 3429.380 ;
        RECT 2524.020 3429.370 2527.020 3429.380 ;
        RECT 2704.020 3429.370 2707.020 3429.380 ;
        RECT 2884.020 3429.370 2887.020 3429.380 ;
        RECT 2926.600 3429.370 2929.600 3429.380 ;
        RECT -9.980 3252.380 -6.980 3252.390 ;
        RECT 4.020 3252.380 7.020 3252.390 ;
        RECT 184.020 3252.380 187.020 3252.390 ;
        RECT 364.020 3252.380 367.020 3252.390 ;
        RECT 544.020 3252.380 547.020 3252.390 ;
        RECT 724.020 3252.380 727.020 3252.390 ;
        RECT 904.020 3252.380 907.020 3252.390 ;
        RECT 1084.020 3252.380 1087.020 3252.390 ;
        RECT 1264.020 3252.380 1267.020 3252.390 ;
        RECT 1444.020 3252.380 1447.020 3252.390 ;
        RECT 1624.020 3252.380 1627.020 3252.390 ;
        RECT 1804.020 3252.380 1807.020 3252.390 ;
        RECT 1984.020 3252.380 1987.020 3252.390 ;
        RECT 2164.020 3252.380 2167.020 3252.390 ;
        RECT 2344.020 3252.380 2347.020 3252.390 ;
        RECT 2524.020 3252.380 2527.020 3252.390 ;
        RECT 2704.020 3252.380 2707.020 3252.390 ;
        RECT 2884.020 3252.380 2887.020 3252.390 ;
        RECT 2926.600 3252.380 2929.600 3252.390 ;
        RECT -14.580 3249.380 2934.200 3252.380 ;
        RECT -9.980 3249.370 -6.980 3249.380 ;
        RECT 4.020 3249.370 7.020 3249.380 ;
        RECT 184.020 3249.370 187.020 3249.380 ;
        RECT 364.020 3249.370 367.020 3249.380 ;
        RECT 544.020 3249.370 547.020 3249.380 ;
        RECT 724.020 3249.370 727.020 3249.380 ;
        RECT 904.020 3249.370 907.020 3249.380 ;
        RECT 1084.020 3249.370 1087.020 3249.380 ;
        RECT 1264.020 3249.370 1267.020 3249.380 ;
        RECT 1444.020 3249.370 1447.020 3249.380 ;
        RECT 1624.020 3249.370 1627.020 3249.380 ;
        RECT 1804.020 3249.370 1807.020 3249.380 ;
        RECT 1984.020 3249.370 1987.020 3249.380 ;
        RECT 2164.020 3249.370 2167.020 3249.380 ;
        RECT 2344.020 3249.370 2347.020 3249.380 ;
        RECT 2524.020 3249.370 2527.020 3249.380 ;
        RECT 2704.020 3249.370 2707.020 3249.380 ;
        RECT 2884.020 3249.370 2887.020 3249.380 ;
        RECT 2926.600 3249.370 2929.600 3249.380 ;
        RECT -9.980 3072.380 -6.980 3072.390 ;
        RECT 4.020 3072.380 7.020 3072.390 ;
        RECT 184.020 3072.380 187.020 3072.390 ;
        RECT 364.020 3072.380 367.020 3072.390 ;
        RECT 544.020 3072.380 547.020 3072.390 ;
        RECT 724.020 3072.380 727.020 3072.390 ;
        RECT 904.020 3072.380 907.020 3072.390 ;
        RECT 1084.020 3072.380 1087.020 3072.390 ;
        RECT 1264.020 3072.380 1267.020 3072.390 ;
        RECT 1444.020 3072.380 1447.020 3072.390 ;
        RECT 1624.020 3072.380 1627.020 3072.390 ;
        RECT 1804.020 3072.380 1807.020 3072.390 ;
        RECT 1984.020 3072.380 1987.020 3072.390 ;
        RECT 2164.020 3072.380 2167.020 3072.390 ;
        RECT 2344.020 3072.380 2347.020 3072.390 ;
        RECT 2524.020 3072.380 2527.020 3072.390 ;
        RECT 2704.020 3072.380 2707.020 3072.390 ;
        RECT 2884.020 3072.380 2887.020 3072.390 ;
        RECT 2926.600 3072.380 2929.600 3072.390 ;
        RECT -14.580 3069.380 2934.200 3072.380 ;
        RECT -9.980 3069.370 -6.980 3069.380 ;
        RECT 4.020 3069.370 7.020 3069.380 ;
        RECT 184.020 3069.370 187.020 3069.380 ;
        RECT 364.020 3069.370 367.020 3069.380 ;
        RECT 544.020 3069.370 547.020 3069.380 ;
        RECT 724.020 3069.370 727.020 3069.380 ;
        RECT 904.020 3069.370 907.020 3069.380 ;
        RECT 1084.020 3069.370 1087.020 3069.380 ;
        RECT 1264.020 3069.370 1267.020 3069.380 ;
        RECT 1444.020 3069.370 1447.020 3069.380 ;
        RECT 1624.020 3069.370 1627.020 3069.380 ;
        RECT 1804.020 3069.370 1807.020 3069.380 ;
        RECT 1984.020 3069.370 1987.020 3069.380 ;
        RECT 2164.020 3069.370 2167.020 3069.380 ;
        RECT 2344.020 3069.370 2347.020 3069.380 ;
        RECT 2524.020 3069.370 2527.020 3069.380 ;
        RECT 2704.020 3069.370 2707.020 3069.380 ;
        RECT 2884.020 3069.370 2887.020 3069.380 ;
        RECT 2926.600 3069.370 2929.600 3069.380 ;
        RECT -9.980 2892.380 -6.980 2892.390 ;
        RECT 4.020 2892.380 7.020 2892.390 ;
        RECT 184.020 2892.380 187.020 2892.390 ;
        RECT 364.020 2892.380 367.020 2892.390 ;
        RECT 544.020 2892.380 547.020 2892.390 ;
        RECT 724.020 2892.380 727.020 2892.390 ;
        RECT 904.020 2892.380 907.020 2892.390 ;
        RECT 1084.020 2892.380 1087.020 2892.390 ;
        RECT 1264.020 2892.380 1267.020 2892.390 ;
        RECT 1444.020 2892.380 1447.020 2892.390 ;
        RECT 1624.020 2892.380 1627.020 2892.390 ;
        RECT 1804.020 2892.380 1807.020 2892.390 ;
        RECT 1984.020 2892.380 1987.020 2892.390 ;
        RECT 2164.020 2892.380 2167.020 2892.390 ;
        RECT 2344.020 2892.380 2347.020 2892.390 ;
        RECT 2524.020 2892.380 2527.020 2892.390 ;
        RECT 2704.020 2892.380 2707.020 2892.390 ;
        RECT 2884.020 2892.380 2887.020 2892.390 ;
        RECT 2926.600 2892.380 2929.600 2892.390 ;
        RECT -14.580 2889.380 2934.200 2892.380 ;
        RECT -9.980 2889.370 -6.980 2889.380 ;
        RECT 4.020 2889.370 7.020 2889.380 ;
        RECT 184.020 2889.370 187.020 2889.380 ;
        RECT 364.020 2889.370 367.020 2889.380 ;
        RECT 544.020 2889.370 547.020 2889.380 ;
        RECT 724.020 2889.370 727.020 2889.380 ;
        RECT 904.020 2889.370 907.020 2889.380 ;
        RECT 1084.020 2889.370 1087.020 2889.380 ;
        RECT 1264.020 2889.370 1267.020 2889.380 ;
        RECT 1444.020 2889.370 1447.020 2889.380 ;
        RECT 1624.020 2889.370 1627.020 2889.380 ;
        RECT 1804.020 2889.370 1807.020 2889.380 ;
        RECT 1984.020 2889.370 1987.020 2889.380 ;
        RECT 2164.020 2889.370 2167.020 2889.380 ;
        RECT 2344.020 2889.370 2347.020 2889.380 ;
        RECT 2524.020 2889.370 2527.020 2889.380 ;
        RECT 2704.020 2889.370 2707.020 2889.380 ;
        RECT 2884.020 2889.370 2887.020 2889.380 ;
        RECT 2926.600 2889.370 2929.600 2889.380 ;
        RECT -9.980 2712.380 -6.980 2712.390 ;
        RECT 4.020 2712.380 7.020 2712.390 ;
        RECT 184.020 2712.380 187.020 2712.390 ;
        RECT 364.020 2712.380 367.020 2712.390 ;
        RECT 544.020 2712.380 547.020 2712.390 ;
        RECT 724.020 2712.380 727.020 2712.390 ;
        RECT 904.020 2712.380 907.020 2712.390 ;
        RECT 1084.020 2712.380 1087.020 2712.390 ;
        RECT 1264.020 2712.380 1267.020 2712.390 ;
        RECT 1444.020 2712.380 1447.020 2712.390 ;
        RECT 1624.020 2712.380 1627.020 2712.390 ;
        RECT 1804.020 2712.380 1807.020 2712.390 ;
        RECT 1984.020 2712.380 1987.020 2712.390 ;
        RECT 2164.020 2712.380 2167.020 2712.390 ;
        RECT 2344.020 2712.380 2347.020 2712.390 ;
        RECT 2524.020 2712.380 2527.020 2712.390 ;
        RECT 2704.020 2712.380 2707.020 2712.390 ;
        RECT 2884.020 2712.380 2887.020 2712.390 ;
        RECT 2926.600 2712.380 2929.600 2712.390 ;
        RECT -14.580 2709.380 2934.200 2712.380 ;
        RECT -9.980 2709.370 -6.980 2709.380 ;
        RECT 4.020 2709.370 7.020 2709.380 ;
        RECT 184.020 2709.370 187.020 2709.380 ;
        RECT 364.020 2709.370 367.020 2709.380 ;
        RECT 544.020 2709.370 547.020 2709.380 ;
        RECT 724.020 2709.370 727.020 2709.380 ;
        RECT 904.020 2709.370 907.020 2709.380 ;
        RECT 1084.020 2709.370 1087.020 2709.380 ;
        RECT 1264.020 2709.370 1267.020 2709.380 ;
        RECT 1444.020 2709.370 1447.020 2709.380 ;
        RECT 1624.020 2709.370 1627.020 2709.380 ;
        RECT 1804.020 2709.370 1807.020 2709.380 ;
        RECT 1984.020 2709.370 1987.020 2709.380 ;
        RECT 2164.020 2709.370 2167.020 2709.380 ;
        RECT 2344.020 2709.370 2347.020 2709.380 ;
        RECT 2524.020 2709.370 2527.020 2709.380 ;
        RECT 2704.020 2709.370 2707.020 2709.380 ;
        RECT 2884.020 2709.370 2887.020 2709.380 ;
        RECT 2926.600 2709.370 2929.600 2709.380 ;
        RECT -9.980 2532.380 -6.980 2532.390 ;
        RECT 4.020 2532.380 7.020 2532.390 ;
        RECT 184.020 2532.380 187.020 2532.390 ;
        RECT 364.020 2532.380 367.020 2532.390 ;
        RECT 544.020 2532.380 547.020 2532.390 ;
        RECT 724.020 2532.380 727.020 2532.390 ;
        RECT 904.020 2532.380 907.020 2532.390 ;
        RECT 1084.020 2532.380 1087.020 2532.390 ;
        RECT 1264.020 2532.380 1267.020 2532.390 ;
        RECT 1444.020 2532.380 1447.020 2532.390 ;
        RECT 1624.020 2532.380 1627.020 2532.390 ;
        RECT 1804.020 2532.380 1807.020 2532.390 ;
        RECT 1984.020 2532.380 1987.020 2532.390 ;
        RECT 2164.020 2532.380 2167.020 2532.390 ;
        RECT 2344.020 2532.380 2347.020 2532.390 ;
        RECT 2524.020 2532.380 2527.020 2532.390 ;
        RECT 2704.020 2532.380 2707.020 2532.390 ;
        RECT 2884.020 2532.380 2887.020 2532.390 ;
        RECT 2926.600 2532.380 2929.600 2532.390 ;
        RECT -14.580 2529.380 2934.200 2532.380 ;
        RECT -9.980 2529.370 -6.980 2529.380 ;
        RECT 4.020 2529.370 7.020 2529.380 ;
        RECT 184.020 2529.370 187.020 2529.380 ;
        RECT 364.020 2529.370 367.020 2529.380 ;
        RECT 544.020 2529.370 547.020 2529.380 ;
        RECT 724.020 2529.370 727.020 2529.380 ;
        RECT 904.020 2529.370 907.020 2529.380 ;
        RECT 1084.020 2529.370 1087.020 2529.380 ;
        RECT 1264.020 2529.370 1267.020 2529.380 ;
        RECT 1444.020 2529.370 1447.020 2529.380 ;
        RECT 1624.020 2529.370 1627.020 2529.380 ;
        RECT 1804.020 2529.370 1807.020 2529.380 ;
        RECT 1984.020 2529.370 1987.020 2529.380 ;
        RECT 2164.020 2529.370 2167.020 2529.380 ;
        RECT 2344.020 2529.370 2347.020 2529.380 ;
        RECT 2524.020 2529.370 2527.020 2529.380 ;
        RECT 2704.020 2529.370 2707.020 2529.380 ;
        RECT 2884.020 2529.370 2887.020 2529.380 ;
        RECT 2926.600 2529.370 2929.600 2529.380 ;
        RECT -9.980 2352.380 -6.980 2352.390 ;
        RECT 4.020 2352.380 7.020 2352.390 ;
        RECT 184.020 2352.380 187.020 2352.390 ;
        RECT 364.020 2352.380 367.020 2352.390 ;
        RECT 544.020 2352.380 547.020 2352.390 ;
        RECT 724.020 2352.380 727.020 2352.390 ;
        RECT 904.020 2352.380 907.020 2352.390 ;
        RECT 1084.020 2352.380 1087.020 2352.390 ;
        RECT 1264.020 2352.380 1267.020 2352.390 ;
        RECT 1444.020 2352.380 1447.020 2352.390 ;
        RECT 1624.020 2352.380 1627.020 2352.390 ;
        RECT 1804.020 2352.380 1807.020 2352.390 ;
        RECT 1984.020 2352.380 1987.020 2352.390 ;
        RECT 2164.020 2352.380 2167.020 2352.390 ;
        RECT 2344.020 2352.380 2347.020 2352.390 ;
        RECT 2524.020 2352.380 2527.020 2352.390 ;
        RECT 2704.020 2352.380 2707.020 2352.390 ;
        RECT 2884.020 2352.380 2887.020 2352.390 ;
        RECT 2926.600 2352.380 2929.600 2352.390 ;
        RECT -14.580 2349.380 2934.200 2352.380 ;
        RECT -9.980 2349.370 -6.980 2349.380 ;
        RECT 4.020 2349.370 7.020 2349.380 ;
        RECT 184.020 2349.370 187.020 2349.380 ;
        RECT 364.020 2349.370 367.020 2349.380 ;
        RECT 544.020 2349.370 547.020 2349.380 ;
        RECT 724.020 2349.370 727.020 2349.380 ;
        RECT 904.020 2349.370 907.020 2349.380 ;
        RECT 1084.020 2349.370 1087.020 2349.380 ;
        RECT 1264.020 2349.370 1267.020 2349.380 ;
        RECT 1444.020 2349.370 1447.020 2349.380 ;
        RECT 1624.020 2349.370 1627.020 2349.380 ;
        RECT 1804.020 2349.370 1807.020 2349.380 ;
        RECT 1984.020 2349.370 1987.020 2349.380 ;
        RECT 2164.020 2349.370 2167.020 2349.380 ;
        RECT 2344.020 2349.370 2347.020 2349.380 ;
        RECT 2524.020 2349.370 2527.020 2349.380 ;
        RECT 2704.020 2349.370 2707.020 2349.380 ;
        RECT 2884.020 2349.370 2887.020 2349.380 ;
        RECT 2926.600 2349.370 2929.600 2349.380 ;
        RECT -9.980 2172.380 -6.980 2172.390 ;
        RECT 4.020 2172.380 7.020 2172.390 ;
        RECT 184.020 2172.380 187.020 2172.390 ;
        RECT 364.020 2172.380 367.020 2172.390 ;
        RECT 544.020 2172.380 547.020 2172.390 ;
        RECT 724.020 2172.380 727.020 2172.390 ;
        RECT 904.020 2172.380 907.020 2172.390 ;
        RECT 1084.020 2172.380 1087.020 2172.390 ;
        RECT 1264.020 2172.380 1267.020 2172.390 ;
        RECT 1444.020 2172.380 1447.020 2172.390 ;
        RECT 1624.020 2172.380 1627.020 2172.390 ;
        RECT 1804.020 2172.380 1807.020 2172.390 ;
        RECT 1984.020 2172.380 1987.020 2172.390 ;
        RECT 2164.020 2172.380 2167.020 2172.390 ;
        RECT 2344.020 2172.380 2347.020 2172.390 ;
        RECT 2524.020 2172.380 2527.020 2172.390 ;
        RECT 2704.020 2172.380 2707.020 2172.390 ;
        RECT 2884.020 2172.380 2887.020 2172.390 ;
        RECT 2926.600 2172.380 2929.600 2172.390 ;
        RECT -14.580 2169.380 2934.200 2172.380 ;
        RECT -9.980 2169.370 -6.980 2169.380 ;
        RECT 4.020 2169.370 7.020 2169.380 ;
        RECT 184.020 2169.370 187.020 2169.380 ;
        RECT 364.020 2169.370 367.020 2169.380 ;
        RECT 544.020 2169.370 547.020 2169.380 ;
        RECT 724.020 2169.370 727.020 2169.380 ;
        RECT 904.020 2169.370 907.020 2169.380 ;
        RECT 1084.020 2169.370 1087.020 2169.380 ;
        RECT 1264.020 2169.370 1267.020 2169.380 ;
        RECT 1444.020 2169.370 1447.020 2169.380 ;
        RECT 1624.020 2169.370 1627.020 2169.380 ;
        RECT 1804.020 2169.370 1807.020 2169.380 ;
        RECT 1984.020 2169.370 1987.020 2169.380 ;
        RECT 2164.020 2169.370 2167.020 2169.380 ;
        RECT 2344.020 2169.370 2347.020 2169.380 ;
        RECT 2524.020 2169.370 2527.020 2169.380 ;
        RECT 2704.020 2169.370 2707.020 2169.380 ;
        RECT 2884.020 2169.370 2887.020 2169.380 ;
        RECT 2926.600 2169.370 2929.600 2169.380 ;
        RECT -9.980 1992.380 -6.980 1992.390 ;
        RECT 4.020 1992.380 7.020 1992.390 ;
        RECT 184.020 1992.380 187.020 1992.390 ;
        RECT 364.020 1992.380 367.020 1992.390 ;
        RECT 544.020 1992.380 547.020 1992.390 ;
        RECT 724.020 1992.380 727.020 1992.390 ;
        RECT 904.020 1992.380 907.020 1992.390 ;
        RECT 1084.020 1992.380 1087.020 1992.390 ;
        RECT 1264.020 1992.380 1267.020 1992.390 ;
        RECT 1444.020 1992.380 1447.020 1992.390 ;
        RECT 1624.020 1992.380 1627.020 1992.390 ;
        RECT 1804.020 1992.380 1807.020 1992.390 ;
        RECT 1984.020 1992.380 1987.020 1992.390 ;
        RECT 2164.020 1992.380 2167.020 1992.390 ;
        RECT 2344.020 1992.380 2347.020 1992.390 ;
        RECT 2524.020 1992.380 2527.020 1992.390 ;
        RECT 2704.020 1992.380 2707.020 1992.390 ;
        RECT 2884.020 1992.380 2887.020 1992.390 ;
        RECT 2926.600 1992.380 2929.600 1992.390 ;
        RECT -14.580 1989.380 2934.200 1992.380 ;
        RECT -9.980 1989.370 -6.980 1989.380 ;
        RECT 4.020 1989.370 7.020 1989.380 ;
        RECT 184.020 1989.370 187.020 1989.380 ;
        RECT 364.020 1989.370 367.020 1989.380 ;
        RECT 544.020 1989.370 547.020 1989.380 ;
        RECT 724.020 1989.370 727.020 1989.380 ;
        RECT 904.020 1989.370 907.020 1989.380 ;
        RECT 1084.020 1989.370 1087.020 1989.380 ;
        RECT 1264.020 1989.370 1267.020 1989.380 ;
        RECT 1444.020 1989.370 1447.020 1989.380 ;
        RECT 1624.020 1989.370 1627.020 1989.380 ;
        RECT 1804.020 1989.370 1807.020 1989.380 ;
        RECT 1984.020 1989.370 1987.020 1989.380 ;
        RECT 2164.020 1989.370 2167.020 1989.380 ;
        RECT 2344.020 1989.370 2347.020 1989.380 ;
        RECT 2524.020 1989.370 2527.020 1989.380 ;
        RECT 2704.020 1989.370 2707.020 1989.380 ;
        RECT 2884.020 1989.370 2887.020 1989.380 ;
        RECT 2926.600 1989.370 2929.600 1989.380 ;
        RECT -9.980 1812.380 -6.980 1812.390 ;
        RECT 4.020 1812.380 7.020 1812.390 ;
        RECT 184.020 1812.380 187.020 1812.390 ;
        RECT 364.020 1812.380 367.020 1812.390 ;
        RECT 544.020 1812.380 547.020 1812.390 ;
        RECT 724.020 1812.380 727.020 1812.390 ;
        RECT 904.020 1812.380 907.020 1812.390 ;
        RECT 1084.020 1812.380 1087.020 1812.390 ;
        RECT 1264.020 1812.380 1267.020 1812.390 ;
        RECT 1444.020 1812.380 1447.020 1812.390 ;
        RECT 1624.020 1812.380 1627.020 1812.390 ;
        RECT 1804.020 1812.380 1807.020 1812.390 ;
        RECT 1984.020 1812.380 1987.020 1812.390 ;
        RECT 2164.020 1812.380 2167.020 1812.390 ;
        RECT 2344.020 1812.380 2347.020 1812.390 ;
        RECT 2524.020 1812.380 2527.020 1812.390 ;
        RECT 2704.020 1812.380 2707.020 1812.390 ;
        RECT 2884.020 1812.380 2887.020 1812.390 ;
        RECT 2926.600 1812.380 2929.600 1812.390 ;
        RECT -14.580 1809.380 2934.200 1812.380 ;
        RECT -9.980 1809.370 -6.980 1809.380 ;
        RECT 4.020 1809.370 7.020 1809.380 ;
        RECT 184.020 1809.370 187.020 1809.380 ;
        RECT 364.020 1809.370 367.020 1809.380 ;
        RECT 544.020 1809.370 547.020 1809.380 ;
        RECT 724.020 1809.370 727.020 1809.380 ;
        RECT 904.020 1809.370 907.020 1809.380 ;
        RECT 1084.020 1809.370 1087.020 1809.380 ;
        RECT 1264.020 1809.370 1267.020 1809.380 ;
        RECT 1444.020 1809.370 1447.020 1809.380 ;
        RECT 1624.020 1809.370 1627.020 1809.380 ;
        RECT 1804.020 1809.370 1807.020 1809.380 ;
        RECT 1984.020 1809.370 1987.020 1809.380 ;
        RECT 2164.020 1809.370 2167.020 1809.380 ;
        RECT 2344.020 1809.370 2347.020 1809.380 ;
        RECT 2524.020 1809.370 2527.020 1809.380 ;
        RECT 2704.020 1809.370 2707.020 1809.380 ;
        RECT 2884.020 1809.370 2887.020 1809.380 ;
        RECT 2926.600 1809.370 2929.600 1809.380 ;
        RECT -9.980 1632.380 -6.980 1632.390 ;
        RECT 4.020 1632.380 7.020 1632.390 ;
        RECT 184.020 1632.380 187.020 1632.390 ;
        RECT 364.020 1632.380 367.020 1632.390 ;
        RECT 544.020 1632.380 547.020 1632.390 ;
        RECT 724.020 1632.380 727.020 1632.390 ;
        RECT 904.020 1632.380 907.020 1632.390 ;
        RECT 1084.020 1632.380 1087.020 1632.390 ;
        RECT 1264.020 1632.380 1267.020 1632.390 ;
        RECT 1444.020 1632.380 1447.020 1632.390 ;
        RECT 1624.020 1632.380 1627.020 1632.390 ;
        RECT 1804.020 1632.380 1807.020 1632.390 ;
        RECT 1984.020 1632.380 1987.020 1632.390 ;
        RECT 2164.020 1632.380 2167.020 1632.390 ;
        RECT 2344.020 1632.380 2347.020 1632.390 ;
        RECT 2524.020 1632.380 2527.020 1632.390 ;
        RECT 2704.020 1632.380 2707.020 1632.390 ;
        RECT 2884.020 1632.380 2887.020 1632.390 ;
        RECT 2926.600 1632.380 2929.600 1632.390 ;
        RECT -14.580 1629.380 2934.200 1632.380 ;
        RECT -9.980 1629.370 -6.980 1629.380 ;
        RECT 4.020 1629.370 7.020 1629.380 ;
        RECT 184.020 1629.370 187.020 1629.380 ;
        RECT 364.020 1629.370 367.020 1629.380 ;
        RECT 544.020 1629.370 547.020 1629.380 ;
        RECT 724.020 1629.370 727.020 1629.380 ;
        RECT 904.020 1629.370 907.020 1629.380 ;
        RECT 1084.020 1629.370 1087.020 1629.380 ;
        RECT 1264.020 1629.370 1267.020 1629.380 ;
        RECT 1444.020 1629.370 1447.020 1629.380 ;
        RECT 1624.020 1629.370 1627.020 1629.380 ;
        RECT 1804.020 1629.370 1807.020 1629.380 ;
        RECT 1984.020 1629.370 1987.020 1629.380 ;
        RECT 2164.020 1629.370 2167.020 1629.380 ;
        RECT 2344.020 1629.370 2347.020 1629.380 ;
        RECT 2524.020 1629.370 2527.020 1629.380 ;
        RECT 2704.020 1629.370 2707.020 1629.380 ;
        RECT 2884.020 1629.370 2887.020 1629.380 ;
        RECT 2926.600 1629.370 2929.600 1629.380 ;
        RECT -9.980 1452.380 -6.980 1452.390 ;
        RECT 4.020 1452.380 7.020 1452.390 ;
        RECT 184.020 1452.380 187.020 1452.390 ;
        RECT 364.020 1452.380 367.020 1452.390 ;
        RECT 544.020 1452.380 547.020 1452.390 ;
        RECT 724.020 1452.380 727.020 1452.390 ;
        RECT 904.020 1452.380 907.020 1452.390 ;
        RECT 1084.020 1452.380 1087.020 1452.390 ;
        RECT 1264.020 1452.380 1267.020 1452.390 ;
        RECT 1444.020 1452.380 1447.020 1452.390 ;
        RECT 1624.020 1452.380 1627.020 1452.390 ;
        RECT 1804.020 1452.380 1807.020 1452.390 ;
        RECT 1984.020 1452.380 1987.020 1452.390 ;
        RECT 2164.020 1452.380 2167.020 1452.390 ;
        RECT 2344.020 1452.380 2347.020 1452.390 ;
        RECT 2524.020 1452.380 2527.020 1452.390 ;
        RECT 2704.020 1452.380 2707.020 1452.390 ;
        RECT 2884.020 1452.380 2887.020 1452.390 ;
        RECT 2926.600 1452.380 2929.600 1452.390 ;
        RECT -14.580 1449.380 2934.200 1452.380 ;
        RECT -9.980 1449.370 -6.980 1449.380 ;
        RECT 4.020 1449.370 7.020 1449.380 ;
        RECT 184.020 1449.370 187.020 1449.380 ;
        RECT 364.020 1449.370 367.020 1449.380 ;
        RECT 544.020 1449.370 547.020 1449.380 ;
        RECT 724.020 1449.370 727.020 1449.380 ;
        RECT 904.020 1449.370 907.020 1449.380 ;
        RECT 1084.020 1449.370 1087.020 1449.380 ;
        RECT 1264.020 1449.370 1267.020 1449.380 ;
        RECT 1444.020 1449.370 1447.020 1449.380 ;
        RECT 1624.020 1449.370 1627.020 1449.380 ;
        RECT 1804.020 1449.370 1807.020 1449.380 ;
        RECT 1984.020 1449.370 1987.020 1449.380 ;
        RECT 2164.020 1449.370 2167.020 1449.380 ;
        RECT 2344.020 1449.370 2347.020 1449.380 ;
        RECT 2524.020 1449.370 2527.020 1449.380 ;
        RECT 2704.020 1449.370 2707.020 1449.380 ;
        RECT 2884.020 1449.370 2887.020 1449.380 ;
        RECT 2926.600 1449.370 2929.600 1449.380 ;
        RECT -9.980 1272.380 -6.980 1272.390 ;
        RECT 4.020 1272.380 7.020 1272.390 ;
        RECT 184.020 1272.380 187.020 1272.390 ;
        RECT 364.020 1272.380 367.020 1272.390 ;
        RECT 544.020 1272.380 547.020 1272.390 ;
        RECT 724.020 1272.380 727.020 1272.390 ;
        RECT 904.020 1272.380 907.020 1272.390 ;
        RECT 1084.020 1272.380 1087.020 1272.390 ;
        RECT 1264.020 1272.380 1267.020 1272.390 ;
        RECT 1444.020 1272.380 1447.020 1272.390 ;
        RECT 1624.020 1272.380 1627.020 1272.390 ;
        RECT 1804.020 1272.380 1807.020 1272.390 ;
        RECT 1984.020 1272.380 1987.020 1272.390 ;
        RECT 2164.020 1272.380 2167.020 1272.390 ;
        RECT 2344.020 1272.380 2347.020 1272.390 ;
        RECT 2524.020 1272.380 2527.020 1272.390 ;
        RECT 2704.020 1272.380 2707.020 1272.390 ;
        RECT 2884.020 1272.380 2887.020 1272.390 ;
        RECT 2926.600 1272.380 2929.600 1272.390 ;
        RECT -14.580 1269.380 2934.200 1272.380 ;
        RECT -9.980 1269.370 -6.980 1269.380 ;
        RECT 4.020 1269.370 7.020 1269.380 ;
        RECT 184.020 1269.370 187.020 1269.380 ;
        RECT 364.020 1269.370 367.020 1269.380 ;
        RECT 544.020 1269.370 547.020 1269.380 ;
        RECT 724.020 1269.370 727.020 1269.380 ;
        RECT 904.020 1269.370 907.020 1269.380 ;
        RECT 1084.020 1269.370 1087.020 1269.380 ;
        RECT 1264.020 1269.370 1267.020 1269.380 ;
        RECT 1444.020 1269.370 1447.020 1269.380 ;
        RECT 1624.020 1269.370 1627.020 1269.380 ;
        RECT 1804.020 1269.370 1807.020 1269.380 ;
        RECT 1984.020 1269.370 1987.020 1269.380 ;
        RECT 2164.020 1269.370 2167.020 1269.380 ;
        RECT 2344.020 1269.370 2347.020 1269.380 ;
        RECT 2524.020 1269.370 2527.020 1269.380 ;
        RECT 2704.020 1269.370 2707.020 1269.380 ;
        RECT 2884.020 1269.370 2887.020 1269.380 ;
        RECT 2926.600 1269.370 2929.600 1269.380 ;
        RECT -9.980 1092.380 -6.980 1092.390 ;
        RECT 4.020 1092.380 7.020 1092.390 ;
        RECT 184.020 1092.380 187.020 1092.390 ;
        RECT 364.020 1092.380 367.020 1092.390 ;
        RECT 544.020 1092.380 547.020 1092.390 ;
        RECT 724.020 1092.380 727.020 1092.390 ;
        RECT 904.020 1092.380 907.020 1092.390 ;
        RECT 1084.020 1092.380 1087.020 1092.390 ;
        RECT 1264.020 1092.380 1267.020 1092.390 ;
        RECT 1444.020 1092.380 1447.020 1092.390 ;
        RECT 1624.020 1092.380 1627.020 1092.390 ;
        RECT 1804.020 1092.380 1807.020 1092.390 ;
        RECT 1984.020 1092.380 1987.020 1092.390 ;
        RECT 2164.020 1092.380 2167.020 1092.390 ;
        RECT 2344.020 1092.380 2347.020 1092.390 ;
        RECT 2524.020 1092.380 2527.020 1092.390 ;
        RECT 2704.020 1092.380 2707.020 1092.390 ;
        RECT 2884.020 1092.380 2887.020 1092.390 ;
        RECT 2926.600 1092.380 2929.600 1092.390 ;
        RECT -14.580 1089.380 2934.200 1092.380 ;
        RECT -9.980 1089.370 -6.980 1089.380 ;
        RECT 4.020 1089.370 7.020 1089.380 ;
        RECT 184.020 1089.370 187.020 1089.380 ;
        RECT 364.020 1089.370 367.020 1089.380 ;
        RECT 544.020 1089.370 547.020 1089.380 ;
        RECT 724.020 1089.370 727.020 1089.380 ;
        RECT 904.020 1089.370 907.020 1089.380 ;
        RECT 1084.020 1089.370 1087.020 1089.380 ;
        RECT 1264.020 1089.370 1267.020 1089.380 ;
        RECT 1444.020 1089.370 1447.020 1089.380 ;
        RECT 1624.020 1089.370 1627.020 1089.380 ;
        RECT 1804.020 1089.370 1807.020 1089.380 ;
        RECT 1984.020 1089.370 1987.020 1089.380 ;
        RECT 2164.020 1089.370 2167.020 1089.380 ;
        RECT 2344.020 1089.370 2347.020 1089.380 ;
        RECT 2524.020 1089.370 2527.020 1089.380 ;
        RECT 2704.020 1089.370 2707.020 1089.380 ;
        RECT 2884.020 1089.370 2887.020 1089.380 ;
        RECT 2926.600 1089.370 2929.600 1089.380 ;
        RECT -9.980 912.380 -6.980 912.390 ;
        RECT 4.020 912.380 7.020 912.390 ;
        RECT 184.020 912.380 187.020 912.390 ;
        RECT 364.020 912.380 367.020 912.390 ;
        RECT 544.020 912.380 547.020 912.390 ;
        RECT 724.020 912.380 727.020 912.390 ;
        RECT 904.020 912.380 907.020 912.390 ;
        RECT 1084.020 912.380 1087.020 912.390 ;
        RECT 1264.020 912.380 1267.020 912.390 ;
        RECT 1444.020 912.380 1447.020 912.390 ;
        RECT 1624.020 912.380 1627.020 912.390 ;
        RECT 1804.020 912.380 1807.020 912.390 ;
        RECT 1984.020 912.380 1987.020 912.390 ;
        RECT 2164.020 912.380 2167.020 912.390 ;
        RECT 2344.020 912.380 2347.020 912.390 ;
        RECT 2524.020 912.380 2527.020 912.390 ;
        RECT 2704.020 912.380 2707.020 912.390 ;
        RECT 2884.020 912.380 2887.020 912.390 ;
        RECT 2926.600 912.380 2929.600 912.390 ;
        RECT -14.580 909.380 2934.200 912.380 ;
        RECT -9.980 909.370 -6.980 909.380 ;
        RECT 4.020 909.370 7.020 909.380 ;
        RECT 184.020 909.370 187.020 909.380 ;
        RECT 364.020 909.370 367.020 909.380 ;
        RECT 544.020 909.370 547.020 909.380 ;
        RECT 724.020 909.370 727.020 909.380 ;
        RECT 904.020 909.370 907.020 909.380 ;
        RECT 1084.020 909.370 1087.020 909.380 ;
        RECT 1264.020 909.370 1267.020 909.380 ;
        RECT 1444.020 909.370 1447.020 909.380 ;
        RECT 1624.020 909.370 1627.020 909.380 ;
        RECT 1804.020 909.370 1807.020 909.380 ;
        RECT 1984.020 909.370 1987.020 909.380 ;
        RECT 2164.020 909.370 2167.020 909.380 ;
        RECT 2344.020 909.370 2347.020 909.380 ;
        RECT 2524.020 909.370 2527.020 909.380 ;
        RECT 2704.020 909.370 2707.020 909.380 ;
        RECT 2884.020 909.370 2887.020 909.380 ;
        RECT 2926.600 909.370 2929.600 909.380 ;
        RECT -9.980 732.380 -6.980 732.390 ;
        RECT 4.020 732.380 7.020 732.390 ;
        RECT 184.020 732.380 187.020 732.390 ;
        RECT 364.020 732.380 367.020 732.390 ;
        RECT 544.020 732.380 547.020 732.390 ;
        RECT 724.020 732.380 727.020 732.390 ;
        RECT 904.020 732.380 907.020 732.390 ;
        RECT 1084.020 732.380 1087.020 732.390 ;
        RECT 1264.020 732.380 1267.020 732.390 ;
        RECT 1444.020 732.380 1447.020 732.390 ;
        RECT 1624.020 732.380 1627.020 732.390 ;
        RECT 1804.020 732.380 1807.020 732.390 ;
        RECT 1984.020 732.380 1987.020 732.390 ;
        RECT 2164.020 732.380 2167.020 732.390 ;
        RECT 2344.020 732.380 2347.020 732.390 ;
        RECT 2524.020 732.380 2527.020 732.390 ;
        RECT 2704.020 732.380 2707.020 732.390 ;
        RECT 2884.020 732.380 2887.020 732.390 ;
        RECT 2926.600 732.380 2929.600 732.390 ;
        RECT -14.580 729.380 2934.200 732.380 ;
        RECT -9.980 729.370 -6.980 729.380 ;
        RECT 4.020 729.370 7.020 729.380 ;
        RECT 184.020 729.370 187.020 729.380 ;
        RECT 364.020 729.370 367.020 729.380 ;
        RECT 544.020 729.370 547.020 729.380 ;
        RECT 724.020 729.370 727.020 729.380 ;
        RECT 904.020 729.370 907.020 729.380 ;
        RECT 1084.020 729.370 1087.020 729.380 ;
        RECT 1264.020 729.370 1267.020 729.380 ;
        RECT 1444.020 729.370 1447.020 729.380 ;
        RECT 1624.020 729.370 1627.020 729.380 ;
        RECT 1804.020 729.370 1807.020 729.380 ;
        RECT 1984.020 729.370 1987.020 729.380 ;
        RECT 2164.020 729.370 2167.020 729.380 ;
        RECT 2344.020 729.370 2347.020 729.380 ;
        RECT 2524.020 729.370 2527.020 729.380 ;
        RECT 2704.020 729.370 2707.020 729.380 ;
        RECT 2884.020 729.370 2887.020 729.380 ;
        RECT 2926.600 729.370 2929.600 729.380 ;
        RECT -9.980 552.380 -6.980 552.390 ;
        RECT 4.020 552.380 7.020 552.390 ;
        RECT 184.020 552.380 187.020 552.390 ;
        RECT 364.020 552.380 367.020 552.390 ;
        RECT 544.020 552.380 547.020 552.390 ;
        RECT 724.020 552.380 727.020 552.390 ;
        RECT 904.020 552.380 907.020 552.390 ;
        RECT 1084.020 552.380 1087.020 552.390 ;
        RECT 1264.020 552.380 1267.020 552.390 ;
        RECT 1444.020 552.380 1447.020 552.390 ;
        RECT 1624.020 552.380 1627.020 552.390 ;
        RECT 1804.020 552.380 1807.020 552.390 ;
        RECT 1984.020 552.380 1987.020 552.390 ;
        RECT 2164.020 552.380 2167.020 552.390 ;
        RECT 2344.020 552.380 2347.020 552.390 ;
        RECT 2524.020 552.380 2527.020 552.390 ;
        RECT 2704.020 552.380 2707.020 552.390 ;
        RECT 2884.020 552.380 2887.020 552.390 ;
        RECT 2926.600 552.380 2929.600 552.390 ;
        RECT -14.580 549.380 2934.200 552.380 ;
        RECT -9.980 549.370 -6.980 549.380 ;
        RECT 4.020 549.370 7.020 549.380 ;
        RECT 184.020 549.370 187.020 549.380 ;
        RECT 364.020 549.370 367.020 549.380 ;
        RECT 544.020 549.370 547.020 549.380 ;
        RECT 724.020 549.370 727.020 549.380 ;
        RECT 904.020 549.370 907.020 549.380 ;
        RECT 1084.020 549.370 1087.020 549.380 ;
        RECT 1264.020 549.370 1267.020 549.380 ;
        RECT 1444.020 549.370 1447.020 549.380 ;
        RECT 1624.020 549.370 1627.020 549.380 ;
        RECT 1804.020 549.370 1807.020 549.380 ;
        RECT 1984.020 549.370 1987.020 549.380 ;
        RECT 2164.020 549.370 2167.020 549.380 ;
        RECT 2344.020 549.370 2347.020 549.380 ;
        RECT 2524.020 549.370 2527.020 549.380 ;
        RECT 2704.020 549.370 2707.020 549.380 ;
        RECT 2884.020 549.370 2887.020 549.380 ;
        RECT 2926.600 549.370 2929.600 549.380 ;
        RECT -9.980 372.380 -6.980 372.390 ;
        RECT 4.020 372.380 7.020 372.390 ;
        RECT 184.020 372.380 187.020 372.390 ;
        RECT 364.020 372.380 367.020 372.390 ;
        RECT 544.020 372.380 547.020 372.390 ;
        RECT 724.020 372.380 727.020 372.390 ;
        RECT 904.020 372.380 907.020 372.390 ;
        RECT 1084.020 372.380 1087.020 372.390 ;
        RECT 1264.020 372.380 1267.020 372.390 ;
        RECT 1444.020 372.380 1447.020 372.390 ;
        RECT 1624.020 372.380 1627.020 372.390 ;
        RECT 1804.020 372.380 1807.020 372.390 ;
        RECT 1984.020 372.380 1987.020 372.390 ;
        RECT 2164.020 372.380 2167.020 372.390 ;
        RECT 2344.020 372.380 2347.020 372.390 ;
        RECT 2524.020 372.380 2527.020 372.390 ;
        RECT 2704.020 372.380 2707.020 372.390 ;
        RECT 2884.020 372.380 2887.020 372.390 ;
        RECT 2926.600 372.380 2929.600 372.390 ;
        RECT -14.580 369.380 2934.200 372.380 ;
        RECT -9.980 369.370 -6.980 369.380 ;
        RECT 4.020 369.370 7.020 369.380 ;
        RECT 184.020 369.370 187.020 369.380 ;
        RECT 364.020 369.370 367.020 369.380 ;
        RECT 544.020 369.370 547.020 369.380 ;
        RECT 724.020 369.370 727.020 369.380 ;
        RECT 904.020 369.370 907.020 369.380 ;
        RECT 1084.020 369.370 1087.020 369.380 ;
        RECT 1264.020 369.370 1267.020 369.380 ;
        RECT 1444.020 369.370 1447.020 369.380 ;
        RECT 1624.020 369.370 1627.020 369.380 ;
        RECT 1804.020 369.370 1807.020 369.380 ;
        RECT 1984.020 369.370 1987.020 369.380 ;
        RECT 2164.020 369.370 2167.020 369.380 ;
        RECT 2344.020 369.370 2347.020 369.380 ;
        RECT 2524.020 369.370 2527.020 369.380 ;
        RECT 2704.020 369.370 2707.020 369.380 ;
        RECT 2884.020 369.370 2887.020 369.380 ;
        RECT 2926.600 369.370 2929.600 369.380 ;
        RECT -9.980 192.380 -6.980 192.390 ;
        RECT 4.020 192.380 7.020 192.390 ;
        RECT 184.020 192.380 187.020 192.390 ;
        RECT 364.020 192.380 367.020 192.390 ;
        RECT 544.020 192.380 547.020 192.390 ;
        RECT 724.020 192.380 727.020 192.390 ;
        RECT 904.020 192.380 907.020 192.390 ;
        RECT 1084.020 192.380 1087.020 192.390 ;
        RECT 1264.020 192.380 1267.020 192.390 ;
        RECT 1444.020 192.380 1447.020 192.390 ;
        RECT 1624.020 192.380 1627.020 192.390 ;
        RECT 1804.020 192.380 1807.020 192.390 ;
        RECT 1984.020 192.380 1987.020 192.390 ;
        RECT 2164.020 192.380 2167.020 192.390 ;
        RECT 2344.020 192.380 2347.020 192.390 ;
        RECT 2524.020 192.380 2527.020 192.390 ;
        RECT 2704.020 192.380 2707.020 192.390 ;
        RECT 2884.020 192.380 2887.020 192.390 ;
        RECT 2926.600 192.380 2929.600 192.390 ;
        RECT -14.580 189.380 2934.200 192.380 ;
        RECT -9.980 189.370 -6.980 189.380 ;
        RECT 4.020 189.370 7.020 189.380 ;
        RECT 184.020 189.370 187.020 189.380 ;
        RECT 364.020 189.370 367.020 189.380 ;
        RECT 544.020 189.370 547.020 189.380 ;
        RECT 724.020 189.370 727.020 189.380 ;
        RECT 904.020 189.370 907.020 189.380 ;
        RECT 1084.020 189.370 1087.020 189.380 ;
        RECT 1264.020 189.370 1267.020 189.380 ;
        RECT 1444.020 189.370 1447.020 189.380 ;
        RECT 1624.020 189.370 1627.020 189.380 ;
        RECT 1804.020 189.370 1807.020 189.380 ;
        RECT 1984.020 189.370 1987.020 189.380 ;
        RECT 2164.020 189.370 2167.020 189.380 ;
        RECT 2344.020 189.370 2347.020 189.380 ;
        RECT 2524.020 189.370 2527.020 189.380 ;
        RECT 2704.020 189.370 2707.020 189.380 ;
        RECT 2884.020 189.370 2887.020 189.380 ;
        RECT 2926.600 189.370 2929.600 189.380 ;
        RECT -9.980 12.380 -6.980 12.390 ;
        RECT 4.020 12.380 7.020 12.390 ;
        RECT 184.020 12.380 187.020 12.390 ;
        RECT 364.020 12.380 367.020 12.390 ;
        RECT 544.020 12.380 547.020 12.390 ;
        RECT 724.020 12.380 727.020 12.390 ;
        RECT 904.020 12.380 907.020 12.390 ;
        RECT 1084.020 12.380 1087.020 12.390 ;
        RECT 1264.020 12.380 1267.020 12.390 ;
        RECT 1444.020 12.380 1447.020 12.390 ;
        RECT 1624.020 12.380 1627.020 12.390 ;
        RECT 1804.020 12.380 1807.020 12.390 ;
        RECT 1984.020 12.380 1987.020 12.390 ;
        RECT 2164.020 12.380 2167.020 12.390 ;
        RECT 2344.020 12.380 2347.020 12.390 ;
        RECT 2524.020 12.380 2527.020 12.390 ;
        RECT 2704.020 12.380 2707.020 12.390 ;
        RECT 2884.020 12.380 2887.020 12.390 ;
        RECT 2926.600 12.380 2929.600 12.390 ;
        RECT -14.580 9.380 2934.200 12.380 ;
        RECT -9.980 9.370 -6.980 9.380 ;
        RECT 4.020 9.370 7.020 9.380 ;
        RECT 184.020 9.370 187.020 9.380 ;
        RECT 364.020 9.370 367.020 9.380 ;
        RECT 544.020 9.370 547.020 9.380 ;
        RECT 724.020 9.370 727.020 9.380 ;
        RECT 904.020 9.370 907.020 9.380 ;
        RECT 1084.020 9.370 1087.020 9.380 ;
        RECT 1264.020 9.370 1267.020 9.380 ;
        RECT 1444.020 9.370 1447.020 9.380 ;
        RECT 1624.020 9.370 1627.020 9.380 ;
        RECT 1804.020 9.370 1807.020 9.380 ;
        RECT 1984.020 9.370 1987.020 9.380 ;
        RECT 2164.020 9.370 2167.020 9.380 ;
        RECT 2344.020 9.370 2347.020 9.380 ;
        RECT 2524.020 9.370 2527.020 9.380 ;
        RECT 2704.020 9.370 2707.020 9.380 ;
        RECT 2884.020 9.370 2887.020 9.380 ;
        RECT 2926.600 9.370 2929.600 9.380 ;
        RECT -9.980 -1.620 -6.980 -1.610 ;
        RECT 4.020 -1.620 7.020 -1.610 ;
        RECT 184.020 -1.620 187.020 -1.610 ;
        RECT 364.020 -1.620 367.020 -1.610 ;
        RECT 544.020 -1.620 547.020 -1.610 ;
        RECT 724.020 -1.620 727.020 -1.610 ;
        RECT 904.020 -1.620 907.020 -1.610 ;
        RECT 1084.020 -1.620 1087.020 -1.610 ;
        RECT 1264.020 -1.620 1267.020 -1.610 ;
        RECT 1444.020 -1.620 1447.020 -1.610 ;
        RECT 1624.020 -1.620 1627.020 -1.610 ;
        RECT 1804.020 -1.620 1807.020 -1.610 ;
        RECT 1984.020 -1.620 1987.020 -1.610 ;
        RECT 2164.020 -1.620 2167.020 -1.610 ;
        RECT 2344.020 -1.620 2347.020 -1.610 ;
        RECT 2524.020 -1.620 2527.020 -1.610 ;
        RECT 2704.020 -1.620 2707.020 -1.610 ;
        RECT 2884.020 -1.620 2887.020 -1.610 ;
        RECT 2926.600 -1.620 2929.600 -1.610 ;
        RECT -9.980 -4.620 2929.600 -1.620 ;
        RECT -9.980 -4.630 -6.980 -4.620 ;
        RECT 4.020 -4.630 7.020 -4.620 ;
        RECT 184.020 -4.630 187.020 -4.620 ;
        RECT 364.020 -4.630 367.020 -4.620 ;
        RECT 544.020 -4.630 547.020 -4.620 ;
        RECT 724.020 -4.630 727.020 -4.620 ;
        RECT 904.020 -4.630 907.020 -4.620 ;
        RECT 1084.020 -4.630 1087.020 -4.620 ;
        RECT 1264.020 -4.630 1267.020 -4.620 ;
        RECT 1444.020 -4.630 1447.020 -4.620 ;
        RECT 1624.020 -4.630 1627.020 -4.620 ;
        RECT 1804.020 -4.630 1807.020 -4.620 ;
        RECT 1984.020 -4.630 1987.020 -4.620 ;
        RECT 2164.020 -4.630 2167.020 -4.620 ;
        RECT 2344.020 -4.630 2347.020 -4.620 ;
        RECT 2524.020 -4.630 2527.020 -4.620 ;
        RECT 2704.020 -4.630 2707.020 -4.620 ;
        RECT 2884.020 -4.630 2887.020 -4.620 ;
        RECT 2926.600 -4.630 2929.600 -4.620 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -14.580 -9.220 -11.580 3528.900 ;
        RECT 94.020 -9.220 97.020 3528.900 ;
        RECT 274.020 -9.220 277.020 3528.900 ;
        RECT 454.020 -9.220 457.020 3528.900 ;
        RECT 634.020 -9.220 637.020 3528.900 ;
        RECT 814.020 -9.220 817.020 3528.900 ;
        RECT 994.020 -9.220 997.020 3528.900 ;
        RECT 1174.020 -9.220 1177.020 3528.900 ;
        RECT 1354.020 -9.220 1357.020 3528.900 ;
        RECT 1534.020 -9.220 1537.020 3528.900 ;
        RECT 1714.020 -9.220 1717.020 3528.900 ;
        RECT 1894.020 -9.220 1897.020 3528.900 ;
        RECT 2074.020 -9.220 2077.020 3528.900 ;
        RECT 2254.020 -9.220 2257.020 3528.900 ;
        RECT 2434.020 -9.220 2437.020 3528.900 ;
        RECT 2614.020 -9.220 2617.020 3528.900 ;
        RECT 2794.020 -9.220 2797.020 3528.900 ;
        RECT 2931.200 -9.220 2934.200 3528.900 ;
      LAYER via4 ;
        RECT -13.670 3527.610 -12.490 3528.790 ;
        RECT -13.670 3526.010 -12.490 3527.190 ;
        RECT -13.670 3341.090 -12.490 3342.270 ;
        RECT -13.670 3339.490 -12.490 3340.670 ;
        RECT -13.670 3161.090 -12.490 3162.270 ;
        RECT -13.670 3159.490 -12.490 3160.670 ;
        RECT -13.670 2981.090 -12.490 2982.270 ;
        RECT -13.670 2979.490 -12.490 2980.670 ;
        RECT -13.670 2801.090 -12.490 2802.270 ;
        RECT -13.670 2799.490 -12.490 2800.670 ;
        RECT -13.670 2621.090 -12.490 2622.270 ;
        RECT -13.670 2619.490 -12.490 2620.670 ;
        RECT -13.670 2441.090 -12.490 2442.270 ;
        RECT -13.670 2439.490 -12.490 2440.670 ;
        RECT -13.670 2261.090 -12.490 2262.270 ;
        RECT -13.670 2259.490 -12.490 2260.670 ;
        RECT -13.670 2081.090 -12.490 2082.270 ;
        RECT -13.670 2079.490 -12.490 2080.670 ;
        RECT -13.670 1901.090 -12.490 1902.270 ;
        RECT -13.670 1899.490 -12.490 1900.670 ;
        RECT -13.670 1721.090 -12.490 1722.270 ;
        RECT -13.670 1719.490 -12.490 1720.670 ;
        RECT -13.670 1541.090 -12.490 1542.270 ;
        RECT -13.670 1539.490 -12.490 1540.670 ;
        RECT -13.670 1361.090 -12.490 1362.270 ;
        RECT -13.670 1359.490 -12.490 1360.670 ;
        RECT -13.670 1181.090 -12.490 1182.270 ;
        RECT -13.670 1179.490 -12.490 1180.670 ;
        RECT -13.670 1001.090 -12.490 1002.270 ;
        RECT -13.670 999.490 -12.490 1000.670 ;
        RECT -13.670 821.090 -12.490 822.270 ;
        RECT -13.670 819.490 -12.490 820.670 ;
        RECT -13.670 641.090 -12.490 642.270 ;
        RECT -13.670 639.490 -12.490 640.670 ;
        RECT -13.670 461.090 -12.490 462.270 ;
        RECT -13.670 459.490 -12.490 460.670 ;
        RECT -13.670 281.090 -12.490 282.270 ;
        RECT -13.670 279.490 -12.490 280.670 ;
        RECT -13.670 101.090 -12.490 102.270 ;
        RECT -13.670 99.490 -12.490 100.670 ;
        RECT -13.670 -7.510 -12.490 -6.330 ;
        RECT -13.670 -9.110 -12.490 -7.930 ;
        RECT 94.930 3527.610 96.110 3528.790 ;
        RECT 94.930 3526.010 96.110 3527.190 ;
        RECT 94.930 3341.090 96.110 3342.270 ;
        RECT 94.930 3339.490 96.110 3340.670 ;
        RECT 94.930 3161.090 96.110 3162.270 ;
        RECT 94.930 3159.490 96.110 3160.670 ;
        RECT 94.930 2981.090 96.110 2982.270 ;
        RECT 94.930 2979.490 96.110 2980.670 ;
        RECT 94.930 2801.090 96.110 2802.270 ;
        RECT 94.930 2799.490 96.110 2800.670 ;
        RECT 94.930 2621.090 96.110 2622.270 ;
        RECT 94.930 2619.490 96.110 2620.670 ;
        RECT 94.930 2441.090 96.110 2442.270 ;
        RECT 94.930 2439.490 96.110 2440.670 ;
        RECT 94.930 2261.090 96.110 2262.270 ;
        RECT 94.930 2259.490 96.110 2260.670 ;
        RECT 94.930 2081.090 96.110 2082.270 ;
        RECT 94.930 2079.490 96.110 2080.670 ;
        RECT 94.930 1901.090 96.110 1902.270 ;
        RECT 94.930 1899.490 96.110 1900.670 ;
        RECT 94.930 1721.090 96.110 1722.270 ;
        RECT 94.930 1719.490 96.110 1720.670 ;
        RECT 94.930 1541.090 96.110 1542.270 ;
        RECT 94.930 1539.490 96.110 1540.670 ;
        RECT 94.930 1361.090 96.110 1362.270 ;
        RECT 94.930 1359.490 96.110 1360.670 ;
        RECT 94.930 1181.090 96.110 1182.270 ;
        RECT 94.930 1179.490 96.110 1180.670 ;
        RECT 94.930 1001.090 96.110 1002.270 ;
        RECT 94.930 999.490 96.110 1000.670 ;
        RECT 94.930 821.090 96.110 822.270 ;
        RECT 94.930 819.490 96.110 820.670 ;
        RECT 94.930 641.090 96.110 642.270 ;
        RECT 94.930 639.490 96.110 640.670 ;
        RECT 94.930 461.090 96.110 462.270 ;
        RECT 94.930 459.490 96.110 460.670 ;
        RECT 94.930 281.090 96.110 282.270 ;
        RECT 94.930 279.490 96.110 280.670 ;
        RECT 94.930 101.090 96.110 102.270 ;
        RECT 94.930 99.490 96.110 100.670 ;
        RECT 94.930 -7.510 96.110 -6.330 ;
        RECT 94.930 -9.110 96.110 -7.930 ;
        RECT 274.930 3527.610 276.110 3528.790 ;
        RECT 274.930 3526.010 276.110 3527.190 ;
        RECT 274.930 3341.090 276.110 3342.270 ;
        RECT 274.930 3339.490 276.110 3340.670 ;
        RECT 274.930 3161.090 276.110 3162.270 ;
        RECT 274.930 3159.490 276.110 3160.670 ;
        RECT 274.930 2981.090 276.110 2982.270 ;
        RECT 274.930 2979.490 276.110 2980.670 ;
        RECT 274.930 2801.090 276.110 2802.270 ;
        RECT 274.930 2799.490 276.110 2800.670 ;
        RECT 274.930 2621.090 276.110 2622.270 ;
        RECT 274.930 2619.490 276.110 2620.670 ;
        RECT 274.930 2441.090 276.110 2442.270 ;
        RECT 274.930 2439.490 276.110 2440.670 ;
        RECT 274.930 2261.090 276.110 2262.270 ;
        RECT 274.930 2259.490 276.110 2260.670 ;
        RECT 274.930 2081.090 276.110 2082.270 ;
        RECT 274.930 2079.490 276.110 2080.670 ;
        RECT 274.930 1901.090 276.110 1902.270 ;
        RECT 274.930 1899.490 276.110 1900.670 ;
        RECT 274.930 1721.090 276.110 1722.270 ;
        RECT 274.930 1719.490 276.110 1720.670 ;
        RECT 274.930 1541.090 276.110 1542.270 ;
        RECT 274.930 1539.490 276.110 1540.670 ;
        RECT 274.930 1361.090 276.110 1362.270 ;
        RECT 274.930 1359.490 276.110 1360.670 ;
        RECT 274.930 1181.090 276.110 1182.270 ;
        RECT 274.930 1179.490 276.110 1180.670 ;
        RECT 274.930 1001.090 276.110 1002.270 ;
        RECT 274.930 999.490 276.110 1000.670 ;
        RECT 274.930 821.090 276.110 822.270 ;
        RECT 274.930 819.490 276.110 820.670 ;
        RECT 274.930 641.090 276.110 642.270 ;
        RECT 274.930 639.490 276.110 640.670 ;
        RECT 274.930 461.090 276.110 462.270 ;
        RECT 274.930 459.490 276.110 460.670 ;
        RECT 274.930 281.090 276.110 282.270 ;
        RECT 274.930 279.490 276.110 280.670 ;
        RECT 274.930 101.090 276.110 102.270 ;
        RECT 274.930 99.490 276.110 100.670 ;
        RECT 274.930 -7.510 276.110 -6.330 ;
        RECT 274.930 -9.110 276.110 -7.930 ;
        RECT 454.930 3527.610 456.110 3528.790 ;
        RECT 454.930 3526.010 456.110 3527.190 ;
        RECT 454.930 3341.090 456.110 3342.270 ;
        RECT 454.930 3339.490 456.110 3340.670 ;
        RECT 454.930 3161.090 456.110 3162.270 ;
        RECT 454.930 3159.490 456.110 3160.670 ;
        RECT 454.930 2981.090 456.110 2982.270 ;
        RECT 454.930 2979.490 456.110 2980.670 ;
        RECT 454.930 2801.090 456.110 2802.270 ;
        RECT 454.930 2799.490 456.110 2800.670 ;
        RECT 454.930 2621.090 456.110 2622.270 ;
        RECT 454.930 2619.490 456.110 2620.670 ;
        RECT 454.930 2441.090 456.110 2442.270 ;
        RECT 454.930 2439.490 456.110 2440.670 ;
        RECT 454.930 2261.090 456.110 2262.270 ;
        RECT 454.930 2259.490 456.110 2260.670 ;
        RECT 454.930 2081.090 456.110 2082.270 ;
        RECT 454.930 2079.490 456.110 2080.670 ;
        RECT 454.930 1901.090 456.110 1902.270 ;
        RECT 454.930 1899.490 456.110 1900.670 ;
        RECT 454.930 1721.090 456.110 1722.270 ;
        RECT 454.930 1719.490 456.110 1720.670 ;
        RECT 454.930 1541.090 456.110 1542.270 ;
        RECT 454.930 1539.490 456.110 1540.670 ;
        RECT 454.930 1361.090 456.110 1362.270 ;
        RECT 454.930 1359.490 456.110 1360.670 ;
        RECT 454.930 1181.090 456.110 1182.270 ;
        RECT 454.930 1179.490 456.110 1180.670 ;
        RECT 454.930 1001.090 456.110 1002.270 ;
        RECT 454.930 999.490 456.110 1000.670 ;
        RECT 454.930 821.090 456.110 822.270 ;
        RECT 454.930 819.490 456.110 820.670 ;
        RECT 454.930 641.090 456.110 642.270 ;
        RECT 454.930 639.490 456.110 640.670 ;
        RECT 454.930 461.090 456.110 462.270 ;
        RECT 454.930 459.490 456.110 460.670 ;
        RECT 454.930 281.090 456.110 282.270 ;
        RECT 454.930 279.490 456.110 280.670 ;
        RECT 454.930 101.090 456.110 102.270 ;
        RECT 454.930 99.490 456.110 100.670 ;
        RECT 454.930 -7.510 456.110 -6.330 ;
        RECT 454.930 -9.110 456.110 -7.930 ;
        RECT 634.930 3527.610 636.110 3528.790 ;
        RECT 634.930 3526.010 636.110 3527.190 ;
        RECT 634.930 3341.090 636.110 3342.270 ;
        RECT 634.930 3339.490 636.110 3340.670 ;
        RECT 634.930 3161.090 636.110 3162.270 ;
        RECT 634.930 3159.490 636.110 3160.670 ;
        RECT 634.930 2981.090 636.110 2982.270 ;
        RECT 634.930 2979.490 636.110 2980.670 ;
        RECT 634.930 2801.090 636.110 2802.270 ;
        RECT 634.930 2799.490 636.110 2800.670 ;
        RECT 634.930 2621.090 636.110 2622.270 ;
        RECT 634.930 2619.490 636.110 2620.670 ;
        RECT 634.930 2441.090 636.110 2442.270 ;
        RECT 634.930 2439.490 636.110 2440.670 ;
        RECT 634.930 2261.090 636.110 2262.270 ;
        RECT 634.930 2259.490 636.110 2260.670 ;
        RECT 634.930 2081.090 636.110 2082.270 ;
        RECT 634.930 2079.490 636.110 2080.670 ;
        RECT 634.930 1901.090 636.110 1902.270 ;
        RECT 634.930 1899.490 636.110 1900.670 ;
        RECT 634.930 1721.090 636.110 1722.270 ;
        RECT 634.930 1719.490 636.110 1720.670 ;
        RECT 634.930 1541.090 636.110 1542.270 ;
        RECT 634.930 1539.490 636.110 1540.670 ;
        RECT 634.930 1361.090 636.110 1362.270 ;
        RECT 634.930 1359.490 636.110 1360.670 ;
        RECT 634.930 1181.090 636.110 1182.270 ;
        RECT 634.930 1179.490 636.110 1180.670 ;
        RECT 634.930 1001.090 636.110 1002.270 ;
        RECT 634.930 999.490 636.110 1000.670 ;
        RECT 634.930 821.090 636.110 822.270 ;
        RECT 634.930 819.490 636.110 820.670 ;
        RECT 634.930 641.090 636.110 642.270 ;
        RECT 634.930 639.490 636.110 640.670 ;
        RECT 634.930 461.090 636.110 462.270 ;
        RECT 634.930 459.490 636.110 460.670 ;
        RECT 634.930 281.090 636.110 282.270 ;
        RECT 634.930 279.490 636.110 280.670 ;
        RECT 634.930 101.090 636.110 102.270 ;
        RECT 634.930 99.490 636.110 100.670 ;
        RECT 634.930 -7.510 636.110 -6.330 ;
        RECT 634.930 -9.110 636.110 -7.930 ;
        RECT 814.930 3527.610 816.110 3528.790 ;
        RECT 814.930 3526.010 816.110 3527.190 ;
        RECT 814.930 3341.090 816.110 3342.270 ;
        RECT 814.930 3339.490 816.110 3340.670 ;
        RECT 814.930 3161.090 816.110 3162.270 ;
        RECT 814.930 3159.490 816.110 3160.670 ;
        RECT 814.930 2981.090 816.110 2982.270 ;
        RECT 814.930 2979.490 816.110 2980.670 ;
        RECT 814.930 2801.090 816.110 2802.270 ;
        RECT 814.930 2799.490 816.110 2800.670 ;
        RECT 814.930 2621.090 816.110 2622.270 ;
        RECT 814.930 2619.490 816.110 2620.670 ;
        RECT 814.930 2441.090 816.110 2442.270 ;
        RECT 814.930 2439.490 816.110 2440.670 ;
        RECT 814.930 2261.090 816.110 2262.270 ;
        RECT 814.930 2259.490 816.110 2260.670 ;
        RECT 814.930 2081.090 816.110 2082.270 ;
        RECT 814.930 2079.490 816.110 2080.670 ;
        RECT 814.930 1901.090 816.110 1902.270 ;
        RECT 814.930 1899.490 816.110 1900.670 ;
        RECT 814.930 1721.090 816.110 1722.270 ;
        RECT 814.930 1719.490 816.110 1720.670 ;
        RECT 814.930 1541.090 816.110 1542.270 ;
        RECT 814.930 1539.490 816.110 1540.670 ;
        RECT 814.930 1361.090 816.110 1362.270 ;
        RECT 814.930 1359.490 816.110 1360.670 ;
        RECT 814.930 1181.090 816.110 1182.270 ;
        RECT 814.930 1179.490 816.110 1180.670 ;
        RECT 814.930 1001.090 816.110 1002.270 ;
        RECT 814.930 999.490 816.110 1000.670 ;
        RECT 814.930 821.090 816.110 822.270 ;
        RECT 814.930 819.490 816.110 820.670 ;
        RECT 814.930 641.090 816.110 642.270 ;
        RECT 814.930 639.490 816.110 640.670 ;
        RECT 814.930 461.090 816.110 462.270 ;
        RECT 814.930 459.490 816.110 460.670 ;
        RECT 814.930 281.090 816.110 282.270 ;
        RECT 814.930 279.490 816.110 280.670 ;
        RECT 814.930 101.090 816.110 102.270 ;
        RECT 814.930 99.490 816.110 100.670 ;
        RECT 814.930 -7.510 816.110 -6.330 ;
        RECT 814.930 -9.110 816.110 -7.930 ;
        RECT 994.930 3527.610 996.110 3528.790 ;
        RECT 994.930 3526.010 996.110 3527.190 ;
        RECT 994.930 3341.090 996.110 3342.270 ;
        RECT 994.930 3339.490 996.110 3340.670 ;
        RECT 994.930 3161.090 996.110 3162.270 ;
        RECT 994.930 3159.490 996.110 3160.670 ;
        RECT 994.930 2981.090 996.110 2982.270 ;
        RECT 994.930 2979.490 996.110 2980.670 ;
        RECT 994.930 2801.090 996.110 2802.270 ;
        RECT 994.930 2799.490 996.110 2800.670 ;
        RECT 994.930 2621.090 996.110 2622.270 ;
        RECT 994.930 2619.490 996.110 2620.670 ;
        RECT 994.930 2441.090 996.110 2442.270 ;
        RECT 994.930 2439.490 996.110 2440.670 ;
        RECT 994.930 2261.090 996.110 2262.270 ;
        RECT 994.930 2259.490 996.110 2260.670 ;
        RECT 994.930 2081.090 996.110 2082.270 ;
        RECT 994.930 2079.490 996.110 2080.670 ;
        RECT 994.930 1901.090 996.110 1902.270 ;
        RECT 994.930 1899.490 996.110 1900.670 ;
        RECT 994.930 1721.090 996.110 1722.270 ;
        RECT 994.930 1719.490 996.110 1720.670 ;
        RECT 994.930 1541.090 996.110 1542.270 ;
        RECT 994.930 1539.490 996.110 1540.670 ;
        RECT 994.930 1361.090 996.110 1362.270 ;
        RECT 994.930 1359.490 996.110 1360.670 ;
        RECT 994.930 1181.090 996.110 1182.270 ;
        RECT 994.930 1179.490 996.110 1180.670 ;
        RECT 994.930 1001.090 996.110 1002.270 ;
        RECT 994.930 999.490 996.110 1000.670 ;
        RECT 994.930 821.090 996.110 822.270 ;
        RECT 994.930 819.490 996.110 820.670 ;
        RECT 994.930 641.090 996.110 642.270 ;
        RECT 994.930 639.490 996.110 640.670 ;
        RECT 994.930 461.090 996.110 462.270 ;
        RECT 994.930 459.490 996.110 460.670 ;
        RECT 994.930 281.090 996.110 282.270 ;
        RECT 994.930 279.490 996.110 280.670 ;
        RECT 994.930 101.090 996.110 102.270 ;
        RECT 994.930 99.490 996.110 100.670 ;
        RECT 994.930 -7.510 996.110 -6.330 ;
        RECT 994.930 -9.110 996.110 -7.930 ;
        RECT 1174.930 3527.610 1176.110 3528.790 ;
        RECT 1174.930 3526.010 1176.110 3527.190 ;
        RECT 1174.930 3341.090 1176.110 3342.270 ;
        RECT 1174.930 3339.490 1176.110 3340.670 ;
        RECT 1174.930 3161.090 1176.110 3162.270 ;
        RECT 1174.930 3159.490 1176.110 3160.670 ;
        RECT 1174.930 2981.090 1176.110 2982.270 ;
        RECT 1174.930 2979.490 1176.110 2980.670 ;
        RECT 1174.930 2801.090 1176.110 2802.270 ;
        RECT 1174.930 2799.490 1176.110 2800.670 ;
        RECT 1174.930 2621.090 1176.110 2622.270 ;
        RECT 1174.930 2619.490 1176.110 2620.670 ;
        RECT 1174.930 2441.090 1176.110 2442.270 ;
        RECT 1174.930 2439.490 1176.110 2440.670 ;
        RECT 1174.930 2261.090 1176.110 2262.270 ;
        RECT 1174.930 2259.490 1176.110 2260.670 ;
        RECT 1174.930 2081.090 1176.110 2082.270 ;
        RECT 1174.930 2079.490 1176.110 2080.670 ;
        RECT 1174.930 1901.090 1176.110 1902.270 ;
        RECT 1174.930 1899.490 1176.110 1900.670 ;
        RECT 1174.930 1721.090 1176.110 1722.270 ;
        RECT 1174.930 1719.490 1176.110 1720.670 ;
        RECT 1174.930 1541.090 1176.110 1542.270 ;
        RECT 1174.930 1539.490 1176.110 1540.670 ;
        RECT 1174.930 1361.090 1176.110 1362.270 ;
        RECT 1174.930 1359.490 1176.110 1360.670 ;
        RECT 1174.930 1181.090 1176.110 1182.270 ;
        RECT 1174.930 1179.490 1176.110 1180.670 ;
        RECT 1174.930 1001.090 1176.110 1002.270 ;
        RECT 1174.930 999.490 1176.110 1000.670 ;
        RECT 1174.930 821.090 1176.110 822.270 ;
        RECT 1174.930 819.490 1176.110 820.670 ;
        RECT 1174.930 641.090 1176.110 642.270 ;
        RECT 1174.930 639.490 1176.110 640.670 ;
        RECT 1174.930 461.090 1176.110 462.270 ;
        RECT 1174.930 459.490 1176.110 460.670 ;
        RECT 1174.930 281.090 1176.110 282.270 ;
        RECT 1174.930 279.490 1176.110 280.670 ;
        RECT 1174.930 101.090 1176.110 102.270 ;
        RECT 1174.930 99.490 1176.110 100.670 ;
        RECT 1174.930 -7.510 1176.110 -6.330 ;
        RECT 1174.930 -9.110 1176.110 -7.930 ;
        RECT 1354.930 3527.610 1356.110 3528.790 ;
        RECT 1354.930 3526.010 1356.110 3527.190 ;
        RECT 1354.930 3341.090 1356.110 3342.270 ;
        RECT 1354.930 3339.490 1356.110 3340.670 ;
        RECT 1354.930 3161.090 1356.110 3162.270 ;
        RECT 1354.930 3159.490 1356.110 3160.670 ;
        RECT 1354.930 2981.090 1356.110 2982.270 ;
        RECT 1354.930 2979.490 1356.110 2980.670 ;
        RECT 1354.930 2801.090 1356.110 2802.270 ;
        RECT 1354.930 2799.490 1356.110 2800.670 ;
        RECT 1354.930 2621.090 1356.110 2622.270 ;
        RECT 1354.930 2619.490 1356.110 2620.670 ;
        RECT 1354.930 2441.090 1356.110 2442.270 ;
        RECT 1354.930 2439.490 1356.110 2440.670 ;
        RECT 1354.930 2261.090 1356.110 2262.270 ;
        RECT 1354.930 2259.490 1356.110 2260.670 ;
        RECT 1354.930 2081.090 1356.110 2082.270 ;
        RECT 1354.930 2079.490 1356.110 2080.670 ;
        RECT 1354.930 1901.090 1356.110 1902.270 ;
        RECT 1354.930 1899.490 1356.110 1900.670 ;
        RECT 1354.930 1721.090 1356.110 1722.270 ;
        RECT 1354.930 1719.490 1356.110 1720.670 ;
        RECT 1354.930 1541.090 1356.110 1542.270 ;
        RECT 1354.930 1539.490 1356.110 1540.670 ;
        RECT 1354.930 1361.090 1356.110 1362.270 ;
        RECT 1354.930 1359.490 1356.110 1360.670 ;
        RECT 1354.930 1181.090 1356.110 1182.270 ;
        RECT 1354.930 1179.490 1356.110 1180.670 ;
        RECT 1354.930 1001.090 1356.110 1002.270 ;
        RECT 1354.930 999.490 1356.110 1000.670 ;
        RECT 1354.930 821.090 1356.110 822.270 ;
        RECT 1354.930 819.490 1356.110 820.670 ;
        RECT 1354.930 641.090 1356.110 642.270 ;
        RECT 1354.930 639.490 1356.110 640.670 ;
        RECT 1354.930 461.090 1356.110 462.270 ;
        RECT 1354.930 459.490 1356.110 460.670 ;
        RECT 1354.930 281.090 1356.110 282.270 ;
        RECT 1354.930 279.490 1356.110 280.670 ;
        RECT 1354.930 101.090 1356.110 102.270 ;
        RECT 1354.930 99.490 1356.110 100.670 ;
        RECT 1354.930 -7.510 1356.110 -6.330 ;
        RECT 1354.930 -9.110 1356.110 -7.930 ;
        RECT 1534.930 3527.610 1536.110 3528.790 ;
        RECT 1534.930 3526.010 1536.110 3527.190 ;
        RECT 1534.930 3341.090 1536.110 3342.270 ;
        RECT 1534.930 3339.490 1536.110 3340.670 ;
        RECT 1534.930 3161.090 1536.110 3162.270 ;
        RECT 1534.930 3159.490 1536.110 3160.670 ;
        RECT 1534.930 2981.090 1536.110 2982.270 ;
        RECT 1534.930 2979.490 1536.110 2980.670 ;
        RECT 1534.930 2801.090 1536.110 2802.270 ;
        RECT 1534.930 2799.490 1536.110 2800.670 ;
        RECT 1534.930 2621.090 1536.110 2622.270 ;
        RECT 1534.930 2619.490 1536.110 2620.670 ;
        RECT 1534.930 2441.090 1536.110 2442.270 ;
        RECT 1534.930 2439.490 1536.110 2440.670 ;
        RECT 1534.930 2261.090 1536.110 2262.270 ;
        RECT 1534.930 2259.490 1536.110 2260.670 ;
        RECT 1534.930 2081.090 1536.110 2082.270 ;
        RECT 1534.930 2079.490 1536.110 2080.670 ;
        RECT 1534.930 1901.090 1536.110 1902.270 ;
        RECT 1534.930 1899.490 1536.110 1900.670 ;
        RECT 1534.930 1721.090 1536.110 1722.270 ;
        RECT 1534.930 1719.490 1536.110 1720.670 ;
        RECT 1534.930 1541.090 1536.110 1542.270 ;
        RECT 1534.930 1539.490 1536.110 1540.670 ;
        RECT 1534.930 1361.090 1536.110 1362.270 ;
        RECT 1534.930 1359.490 1536.110 1360.670 ;
        RECT 1534.930 1181.090 1536.110 1182.270 ;
        RECT 1534.930 1179.490 1536.110 1180.670 ;
        RECT 1534.930 1001.090 1536.110 1002.270 ;
        RECT 1534.930 999.490 1536.110 1000.670 ;
        RECT 1534.930 821.090 1536.110 822.270 ;
        RECT 1534.930 819.490 1536.110 820.670 ;
        RECT 1534.930 641.090 1536.110 642.270 ;
        RECT 1534.930 639.490 1536.110 640.670 ;
        RECT 1534.930 461.090 1536.110 462.270 ;
        RECT 1534.930 459.490 1536.110 460.670 ;
        RECT 1534.930 281.090 1536.110 282.270 ;
        RECT 1534.930 279.490 1536.110 280.670 ;
        RECT 1534.930 101.090 1536.110 102.270 ;
        RECT 1534.930 99.490 1536.110 100.670 ;
        RECT 1534.930 -7.510 1536.110 -6.330 ;
        RECT 1534.930 -9.110 1536.110 -7.930 ;
        RECT 1714.930 3527.610 1716.110 3528.790 ;
        RECT 1714.930 3526.010 1716.110 3527.190 ;
        RECT 1714.930 3341.090 1716.110 3342.270 ;
        RECT 1714.930 3339.490 1716.110 3340.670 ;
        RECT 1714.930 3161.090 1716.110 3162.270 ;
        RECT 1714.930 3159.490 1716.110 3160.670 ;
        RECT 1714.930 2981.090 1716.110 2982.270 ;
        RECT 1714.930 2979.490 1716.110 2980.670 ;
        RECT 1714.930 2801.090 1716.110 2802.270 ;
        RECT 1714.930 2799.490 1716.110 2800.670 ;
        RECT 1714.930 2621.090 1716.110 2622.270 ;
        RECT 1714.930 2619.490 1716.110 2620.670 ;
        RECT 1714.930 2441.090 1716.110 2442.270 ;
        RECT 1714.930 2439.490 1716.110 2440.670 ;
        RECT 1714.930 2261.090 1716.110 2262.270 ;
        RECT 1714.930 2259.490 1716.110 2260.670 ;
        RECT 1714.930 2081.090 1716.110 2082.270 ;
        RECT 1714.930 2079.490 1716.110 2080.670 ;
        RECT 1714.930 1901.090 1716.110 1902.270 ;
        RECT 1714.930 1899.490 1716.110 1900.670 ;
        RECT 1714.930 1721.090 1716.110 1722.270 ;
        RECT 1714.930 1719.490 1716.110 1720.670 ;
        RECT 1714.930 1541.090 1716.110 1542.270 ;
        RECT 1714.930 1539.490 1716.110 1540.670 ;
        RECT 1714.930 1361.090 1716.110 1362.270 ;
        RECT 1714.930 1359.490 1716.110 1360.670 ;
        RECT 1714.930 1181.090 1716.110 1182.270 ;
        RECT 1714.930 1179.490 1716.110 1180.670 ;
        RECT 1714.930 1001.090 1716.110 1002.270 ;
        RECT 1714.930 999.490 1716.110 1000.670 ;
        RECT 1714.930 821.090 1716.110 822.270 ;
        RECT 1714.930 819.490 1716.110 820.670 ;
        RECT 1714.930 641.090 1716.110 642.270 ;
        RECT 1714.930 639.490 1716.110 640.670 ;
        RECT 1714.930 461.090 1716.110 462.270 ;
        RECT 1714.930 459.490 1716.110 460.670 ;
        RECT 1714.930 281.090 1716.110 282.270 ;
        RECT 1714.930 279.490 1716.110 280.670 ;
        RECT 1714.930 101.090 1716.110 102.270 ;
        RECT 1714.930 99.490 1716.110 100.670 ;
        RECT 1714.930 -7.510 1716.110 -6.330 ;
        RECT 1714.930 -9.110 1716.110 -7.930 ;
        RECT 1894.930 3527.610 1896.110 3528.790 ;
        RECT 1894.930 3526.010 1896.110 3527.190 ;
        RECT 1894.930 3341.090 1896.110 3342.270 ;
        RECT 1894.930 3339.490 1896.110 3340.670 ;
        RECT 1894.930 3161.090 1896.110 3162.270 ;
        RECT 1894.930 3159.490 1896.110 3160.670 ;
        RECT 1894.930 2981.090 1896.110 2982.270 ;
        RECT 1894.930 2979.490 1896.110 2980.670 ;
        RECT 1894.930 2801.090 1896.110 2802.270 ;
        RECT 1894.930 2799.490 1896.110 2800.670 ;
        RECT 1894.930 2621.090 1896.110 2622.270 ;
        RECT 1894.930 2619.490 1896.110 2620.670 ;
        RECT 1894.930 2441.090 1896.110 2442.270 ;
        RECT 1894.930 2439.490 1896.110 2440.670 ;
        RECT 1894.930 2261.090 1896.110 2262.270 ;
        RECT 1894.930 2259.490 1896.110 2260.670 ;
        RECT 1894.930 2081.090 1896.110 2082.270 ;
        RECT 1894.930 2079.490 1896.110 2080.670 ;
        RECT 1894.930 1901.090 1896.110 1902.270 ;
        RECT 1894.930 1899.490 1896.110 1900.670 ;
        RECT 1894.930 1721.090 1896.110 1722.270 ;
        RECT 1894.930 1719.490 1896.110 1720.670 ;
        RECT 1894.930 1541.090 1896.110 1542.270 ;
        RECT 1894.930 1539.490 1896.110 1540.670 ;
        RECT 1894.930 1361.090 1896.110 1362.270 ;
        RECT 1894.930 1359.490 1896.110 1360.670 ;
        RECT 1894.930 1181.090 1896.110 1182.270 ;
        RECT 1894.930 1179.490 1896.110 1180.670 ;
        RECT 1894.930 1001.090 1896.110 1002.270 ;
        RECT 1894.930 999.490 1896.110 1000.670 ;
        RECT 1894.930 821.090 1896.110 822.270 ;
        RECT 1894.930 819.490 1896.110 820.670 ;
        RECT 1894.930 641.090 1896.110 642.270 ;
        RECT 1894.930 639.490 1896.110 640.670 ;
        RECT 1894.930 461.090 1896.110 462.270 ;
        RECT 1894.930 459.490 1896.110 460.670 ;
        RECT 1894.930 281.090 1896.110 282.270 ;
        RECT 1894.930 279.490 1896.110 280.670 ;
        RECT 1894.930 101.090 1896.110 102.270 ;
        RECT 1894.930 99.490 1896.110 100.670 ;
        RECT 1894.930 -7.510 1896.110 -6.330 ;
        RECT 1894.930 -9.110 1896.110 -7.930 ;
        RECT 2074.930 3527.610 2076.110 3528.790 ;
        RECT 2074.930 3526.010 2076.110 3527.190 ;
        RECT 2074.930 3341.090 2076.110 3342.270 ;
        RECT 2074.930 3339.490 2076.110 3340.670 ;
        RECT 2074.930 3161.090 2076.110 3162.270 ;
        RECT 2074.930 3159.490 2076.110 3160.670 ;
        RECT 2074.930 2981.090 2076.110 2982.270 ;
        RECT 2074.930 2979.490 2076.110 2980.670 ;
        RECT 2074.930 2801.090 2076.110 2802.270 ;
        RECT 2074.930 2799.490 2076.110 2800.670 ;
        RECT 2074.930 2621.090 2076.110 2622.270 ;
        RECT 2074.930 2619.490 2076.110 2620.670 ;
        RECT 2074.930 2441.090 2076.110 2442.270 ;
        RECT 2074.930 2439.490 2076.110 2440.670 ;
        RECT 2074.930 2261.090 2076.110 2262.270 ;
        RECT 2074.930 2259.490 2076.110 2260.670 ;
        RECT 2074.930 2081.090 2076.110 2082.270 ;
        RECT 2074.930 2079.490 2076.110 2080.670 ;
        RECT 2074.930 1901.090 2076.110 1902.270 ;
        RECT 2074.930 1899.490 2076.110 1900.670 ;
        RECT 2074.930 1721.090 2076.110 1722.270 ;
        RECT 2074.930 1719.490 2076.110 1720.670 ;
        RECT 2074.930 1541.090 2076.110 1542.270 ;
        RECT 2074.930 1539.490 2076.110 1540.670 ;
        RECT 2074.930 1361.090 2076.110 1362.270 ;
        RECT 2074.930 1359.490 2076.110 1360.670 ;
        RECT 2074.930 1181.090 2076.110 1182.270 ;
        RECT 2074.930 1179.490 2076.110 1180.670 ;
        RECT 2074.930 1001.090 2076.110 1002.270 ;
        RECT 2074.930 999.490 2076.110 1000.670 ;
        RECT 2074.930 821.090 2076.110 822.270 ;
        RECT 2074.930 819.490 2076.110 820.670 ;
        RECT 2074.930 641.090 2076.110 642.270 ;
        RECT 2074.930 639.490 2076.110 640.670 ;
        RECT 2074.930 461.090 2076.110 462.270 ;
        RECT 2074.930 459.490 2076.110 460.670 ;
        RECT 2074.930 281.090 2076.110 282.270 ;
        RECT 2074.930 279.490 2076.110 280.670 ;
        RECT 2074.930 101.090 2076.110 102.270 ;
        RECT 2074.930 99.490 2076.110 100.670 ;
        RECT 2074.930 -7.510 2076.110 -6.330 ;
        RECT 2074.930 -9.110 2076.110 -7.930 ;
        RECT 2254.930 3527.610 2256.110 3528.790 ;
        RECT 2254.930 3526.010 2256.110 3527.190 ;
        RECT 2254.930 3341.090 2256.110 3342.270 ;
        RECT 2254.930 3339.490 2256.110 3340.670 ;
        RECT 2254.930 3161.090 2256.110 3162.270 ;
        RECT 2254.930 3159.490 2256.110 3160.670 ;
        RECT 2254.930 2981.090 2256.110 2982.270 ;
        RECT 2254.930 2979.490 2256.110 2980.670 ;
        RECT 2254.930 2801.090 2256.110 2802.270 ;
        RECT 2254.930 2799.490 2256.110 2800.670 ;
        RECT 2254.930 2621.090 2256.110 2622.270 ;
        RECT 2254.930 2619.490 2256.110 2620.670 ;
        RECT 2254.930 2441.090 2256.110 2442.270 ;
        RECT 2254.930 2439.490 2256.110 2440.670 ;
        RECT 2254.930 2261.090 2256.110 2262.270 ;
        RECT 2254.930 2259.490 2256.110 2260.670 ;
        RECT 2254.930 2081.090 2256.110 2082.270 ;
        RECT 2254.930 2079.490 2256.110 2080.670 ;
        RECT 2254.930 1901.090 2256.110 1902.270 ;
        RECT 2254.930 1899.490 2256.110 1900.670 ;
        RECT 2254.930 1721.090 2256.110 1722.270 ;
        RECT 2254.930 1719.490 2256.110 1720.670 ;
        RECT 2254.930 1541.090 2256.110 1542.270 ;
        RECT 2254.930 1539.490 2256.110 1540.670 ;
        RECT 2254.930 1361.090 2256.110 1362.270 ;
        RECT 2254.930 1359.490 2256.110 1360.670 ;
        RECT 2254.930 1181.090 2256.110 1182.270 ;
        RECT 2254.930 1179.490 2256.110 1180.670 ;
        RECT 2254.930 1001.090 2256.110 1002.270 ;
        RECT 2254.930 999.490 2256.110 1000.670 ;
        RECT 2254.930 821.090 2256.110 822.270 ;
        RECT 2254.930 819.490 2256.110 820.670 ;
        RECT 2254.930 641.090 2256.110 642.270 ;
        RECT 2254.930 639.490 2256.110 640.670 ;
        RECT 2254.930 461.090 2256.110 462.270 ;
        RECT 2254.930 459.490 2256.110 460.670 ;
        RECT 2254.930 281.090 2256.110 282.270 ;
        RECT 2254.930 279.490 2256.110 280.670 ;
        RECT 2254.930 101.090 2256.110 102.270 ;
        RECT 2254.930 99.490 2256.110 100.670 ;
        RECT 2254.930 -7.510 2256.110 -6.330 ;
        RECT 2254.930 -9.110 2256.110 -7.930 ;
        RECT 2434.930 3527.610 2436.110 3528.790 ;
        RECT 2434.930 3526.010 2436.110 3527.190 ;
        RECT 2434.930 3341.090 2436.110 3342.270 ;
        RECT 2434.930 3339.490 2436.110 3340.670 ;
        RECT 2434.930 3161.090 2436.110 3162.270 ;
        RECT 2434.930 3159.490 2436.110 3160.670 ;
        RECT 2434.930 2981.090 2436.110 2982.270 ;
        RECT 2434.930 2979.490 2436.110 2980.670 ;
        RECT 2434.930 2801.090 2436.110 2802.270 ;
        RECT 2434.930 2799.490 2436.110 2800.670 ;
        RECT 2434.930 2621.090 2436.110 2622.270 ;
        RECT 2434.930 2619.490 2436.110 2620.670 ;
        RECT 2434.930 2441.090 2436.110 2442.270 ;
        RECT 2434.930 2439.490 2436.110 2440.670 ;
        RECT 2434.930 2261.090 2436.110 2262.270 ;
        RECT 2434.930 2259.490 2436.110 2260.670 ;
        RECT 2434.930 2081.090 2436.110 2082.270 ;
        RECT 2434.930 2079.490 2436.110 2080.670 ;
        RECT 2434.930 1901.090 2436.110 1902.270 ;
        RECT 2434.930 1899.490 2436.110 1900.670 ;
        RECT 2434.930 1721.090 2436.110 1722.270 ;
        RECT 2434.930 1719.490 2436.110 1720.670 ;
        RECT 2434.930 1541.090 2436.110 1542.270 ;
        RECT 2434.930 1539.490 2436.110 1540.670 ;
        RECT 2434.930 1361.090 2436.110 1362.270 ;
        RECT 2434.930 1359.490 2436.110 1360.670 ;
        RECT 2434.930 1181.090 2436.110 1182.270 ;
        RECT 2434.930 1179.490 2436.110 1180.670 ;
        RECT 2434.930 1001.090 2436.110 1002.270 ;
        RECT 2434.930 999.490 2436.110 1000.670 ;
        RECT 2434.930 821.090 2436.110 822.270 ;
        RECT 2434.930 819.490 2436.110 820.670 ;
        RECT 2434.930 641.090 2436.110 642.270 ;
        RECT 2434.930 639.490 2436.110 640.670 ;
        RECT 2434.930 461.090 2436.110 462.270 ;
        RECT 2434.930 459.490 2436.110 460.670 ;
        RECT 2434.930 281.090 2436.110 282.270 ;
        RECT 2434.930 279.490 2436.110 280.670 ;
        RECT 2434.930 101.090 2436.110 102.270 ;
        RECT 2434.930 99.490 2436.110 100.670 ;
        RECT 2434.930 -7.510 2436.110 -6.330 ;
        RECT 2434.930 -9.110 2436.110 -7.930 ;
        RECT 2614.930 3527.610 2616.110 3528.790 ;
        RECT 2614.930 3526.010 2616.110 3527.190 ;
        RECT 2614.930 3341.090 2616.110 3342.270 ;
        RECT 2614.930 3339.490 2616.110 3340.670 ;
        RECT 2614.930 3161.090 2616.110 3162.270 ;
        RECT 2614.930 3159.490 2616.110 3160.670 ;
        RECT 2614.930 2981.090 2616.110 2982.270 ;
        RECT 2614.930 2979.490 2616.110 2980.670 ;
        RECT 2614.930 2801.090 2616.110 2802.270 ;
        RECT 2614.930 2799.490 2616.110 2800.670 ;
        RECT 2614.930 2621.090 2616.110 2622.270 ;
        RECT 2614.930 2619.490 2616.110 2620.670 ;
        RECT 2614.930 2441.090 2616.110 2442.270 ;
        RECT 2614.930 2439.490 2616.110 2440.670 ;
        RECT 2614.930 2261.090 2616.110 2262.270 ;
        RECT 2614.930 2259.490 2616.110 2260.670 ;
        RECT 2614.930 2081.090 2616.110 2082.270 ;
        RECT 2614.930 2079.490 2616.110 2080.670 ;
        RECT 2614.930 1901.090 2616.110 1902.270 ;
        RECT 2614.930 1899.490 2616.110 1900.670 ;
        RECT 2614.930 1721.090 2616.110 1722.270 ;
        RECT 2614.930 1719.490 2616.110 1720.670 ;
        RECT 2614.930 1541.090 2616.110 1542.270 ;
        RECT 2614.930 1539.490 2616.110 1540.670 ;
        RECT 2614.930 1361.090 2616.110 1362.270 ;
        RECT 2614.930 1359.490 2616.110 1360.670 ;
        RECT 2614.930 1181.090 2616.110 1182.270 ;
        RECT 2614.930 1179.490 2616.110 1180.670 ;
        RECT 2614.930 1001.090 2616.110 1002.270 ;
        RECT 2614.930 999.490 2616.110 1000.670 ;
        RECT 2614.930 821.090 2616.110 822.270 ;
        RECT 2614.930 819.490 2616.110 820.670 ;
        RECT 2614.930 641.090 2616.110 642.270 ;
        RECT 2614.930 639.490 2616.110 640.670 ;
        RECT 2614.930 461.090 2616.110 462.270 ;
        RECT 2614.930 459.490 2616.110 460.670 ;
        RECT 2614.930 281.090 2616.110 282.270 ;
        RECT 2614.930 279.490 2616.110 280.670 ;
        RECT 2614.930 101.090 2616.110 102.270 ;
        RECT 2614.930 99.490 2616.110 100.670 ;
        RECT 2614.930 -7.510 2616.110 -6.330 ;
        RECT 2614.930 -9.110 2616.110 -7.930 ;
        RECT 2794.930 3527.610 2796.110 3528.790 ;
        RECT 2794.930 3526.010 2796.110 3527.190 ;
        RECT 2794.930 3341.090 2796.110 3342.270 ;
        RECT 2794.930 3339.490 2796.110 3340.670 ;
        RECT 2794.930 3161.090 2796.110 3162.270 ;
        RECT 2794.930 3159.490 2796.110 3160.670 ;
        RECT 2794.930 2981.090 2796.110 2982.270 ;
        RECT 2794.930 2979.490 2796.110 2980.670 ;
        RECT 2794.930 2801.090 2796.110 2802.270 ;
        RECT 2794.930 2799.490 2796.110 2800.670 ;
        RECT 2794.930 2621.090 2796.110 2622.270 ;
        RECT 2794.930 2619.490 2796.110 2620.670 ;
        RECT 2794.930 2441.090 2796.110 2442.270 ;
        RECT 2794.930 2439.490 2796.110 2440.670 ;
        RECT 2794.930 2261.090 2796.110 2262.270 ;
        RECT 2794.930 2259.490 2796.110 2260.670 ;
        RECT 2794.930 2081.090 2796.110 2082.270 ;
        RECT 2794.930 2079.490 2796.110 2080.670 ;
        RECT 2794.930 1901.090 2796.110 1902.270 ;
        RECT 2794.930 1899.490 2796.110 1900.670 ;
        RECT 2794.930 1721.090 2796.110 1722.270 ;
        RECT 2794.930 1719.490 2796.110 1720.670 ;
        RECT 2794.930 1541.090 2796.110 1542.270 ;
        RECT 2794.930 1539.490 2796.110 1540.670 ;
        RECT 2794.930 1361.090 2796.110 1362.270 ;
        RECT 2794.930 1359.490 2796.110 1360.670 ;
        RECT 2794.930 1181.090 2796.110 1182.270 ;
        RECT 2794.930 1179.490 2796.110 1180.670 ;
        RECT 2794.930 1001.090 2796.110 1002.270 ;
        RECT 2794.930 999.490 2796.110 1000.670 ;
        RECT 2794.930 821.090 2796.110 822.270 ;
        RECT 2794.930 819.490 2796.110 820.670 ;
        RECT 2794.930 641.090 2796.110 642.270 ;
        RECT 2794.930 639.490 2796.110 640.670 ;
        RECT 2794.930 461.090 2796.110 462.270 ;
        RECT 2794.930 459.490 2796.110 460.670 ;
        RECT 2794.930 281.090 2796.110 282.270 ;
        RECT 2794.930 279.490 2796.110 280.670 ;
        RECT 2794.930 101.090 2796.110 102.270 ;
        RECT 2794.930 99.490 2796.110 100.670 ;
        RECT 2794.930 -7.510 2796.110 -6.330 ;
        RECT 2794.930 -9.110 2796.110 -7.930 ;
        RECT 2932.110 3527.610 2933.290 3528.790 ;
        RECT 2932.110 3526.010 2933.290 3527.190 ;
        RECT 2932.110 3341.090 2933.290 3342.270 ;
        RECT 2932.110 3339.490 2933.290 3340.670 ;
        RECT 2932.110 3161.090 2933.290 3162.270 ;
        RECT 2932.110 3159.490 2933.290 3160.670 ;
        RECT 2932.110 2981.090 2933.290 2982.270 ;
        RECT 2932.110 2979.490 2933.290 2980.670 ;
        RECT 2932.110 2801.090 2933.290 2802.270 ;
        RECT 2932.110 2799.490 2933.290 2800.670 ;
        RECT 2932.110 2621.090 2933.290 2622.270 ;
        RECT 2932.110 2619.490 2933.290 2620.670 ;
        RECT 2932.110 2441.090 2933.290 2442.270 ;
        RECT 2932.110 2439.490 2933.290 2440.670 ;
        RECT 2932.110 2261.090 2933.290 2262.270 ;
        RECT 2932.110 2259.490 2933.290 2260.670 ;
        RECT 2932.110 2081.090 2933.290 2082.270 ;
        RECT 2932.110 2079.490 2933.290 2080.670 ;
        RECT 2932.110 1901.090 2933.290 1902.270 ;
        RECT 2932.110 1899.490 2933.290 1900.670 ;
        RECT 2932.110 1721.090 2933.290 1722.270 ;
        RECT 2932.110 1719.490 2933.290 1720.670 ;
        RECT 2932.110 1541.090 2933.290 1542.270 ;
        RECT 2932.110 1539.490 2933.290 1540.670 ;
        RECT 2932.110 1361.090 2933.290 1362.270 ;
        RECT 2932.110 1359.490 2933.290 1360.670 ;
        RECT 2932.110 1181.090 2933.290 1182.270 ;
        RECT 2932.110 1179.490 2933.290 1180.670 ;
        RECT 2932.110 1001.090 2933.290 1002.270 ;
        RECT 2932.110 999.490 2933.290 1000.670 ;
        RECT 2932.110 821.090 2933.290 822.270 ;
        RECT 2932.110 819.490 2933.290 820.670 ;
        RECT 2932.110 641.090 2933.290 642.270 ;
        RECT 2932.110 639.490 2933.290 640.670 ;
        RECT 2932.110 461.090 2933.290 462.270 ;
        RECT 2932.110 459.490 2933.290 460.670 ;
        RECT 2932.110 281.090 2933.290 282.270 ;
        RECT 2932.110 279.490 2933.290 280.670 ;
        RECT 2932.110 101.090 2933.290 102.270 ;
        RECT 2932.110 99.490 2933.290 100.670 ;
        RECT 2932.110 -7.510 2933.290 -6.330 ;
        RECT 2932.110 -9.110 2933.290 -7.930 ;
      LAYER met5 ;
        RECT -14.580 3528.900 -11.580 3528.910 ;
        RECT 94.020 3528.900 97.020 3528.910 ;
        RECT 274.020 3528.900 277.020 3528.910 ;
        RECT 454.020 3528.900 457.020 3528.910 ;
        RECT 634.020 3528.900 637.020 3528.910 ;
        RECT 814.020 3528.900 817.020 3528.910 ;
        RECT 994.020 3528.900 997.020 3528.910 ;
        RECT 1174.020 3528.900 1177.020 3528.910 ;
        RECT 1354.020 3528.900 1357.020 3528.910 ;
        RECT 1534.020 3528.900 1537.020 3528.910 ;
        RECT 1714.020 3528.900 1717.020 3528.910 ;
        RECT 1894.020 3528.900 1897.020 3528.910 ;
        RECT 2074.020 3528.900 2077.020 3528.910 ;
        RECT 2254.020 3528.900 2257.020 3528.910 ;
        RECT 2434.020 3528.900 2437.020 3528.910 ;
        RECT 2614.020 3528.900 2617.020 3528.910 ;
        RECT 2794.020 3528.900 2797.020 3528.910 ;
        RECT 2931.200 3528.900 2934.200 3528.910 ;
        RECT -14.580 3525.900 2934.200 3528.900 ;
        RECT -14.580 3525.890 -11.580 3525.900 ;
        RECT 94.020 3525.890 97.020 3525.900 ;
        RECT 274.020 3525.890 277.020 3525.900 ;
        RECT 454.020 3525.890 457.020 3525.900 ;
        RECT 634.020 3525.890 637.020 3525.900 ;
        RECT 814.020 3525.890 817.020 3525.900 ;
        RECT 994.020 3525.890 997.020 3525.900 ;
        RECT 1174.020 3525.890 1177.020 3525.900 ;
        RECT 1354.020 3525.890 1357.020 3525.900 ;
        RECT 1534.020 3525.890 1537.020 3525.900 ;
        RECT 1714.020 3525.890 1717.020 3525.900 ;
        RECT 1894.020 3525.890 1897.020 3525.900 ;
        RECT 2074.020 3525.890 2077.020 3525.900 ;
        RECT 2254.020 3525.890 2257.020 3525.900 ;
        RECT 2434.020 3525.890 2437.020 3525.900 ;
        RECT 2614.020 3525.890 2617.020 3525.900 ;
        RECT 2794.020 3525.890 2797.020 3525.900 ;
        RECT 2931.200 3525.890 2934.200 3525.900 ;
        RECT -14.580 3342.380 -11.580 3342.390 ;
        RECT 94.020 3342.380 97.020 3342.390 ;
        RECT 274.020 3342.380 277.020 3342.390 ;
        RECT 454.020 3342.380 457.020 3342.390 ;
        RECT 634.020 3342.380 637.020 3342.390 ;
        RECT 814.020 3342.380 817.020 3342.390 ;
        RECT 994.020 3342.380 997.020 3342.390 ;
        RECT 1174.020 3342.380 1177.020 3342.390 ;
        RECT 1354.020 3342.380 1357.020 3342.390 ;
        RECT 1534.020 3342.380 1537.020 3342.390 ;
        RECT 1714.020 3342.380 1717.020 3342.390 ;
        RECT 1894.020 3342.380 1897.020 3342.390 ;
        RECT 2074.020 3342.380 2077.020 3342.390 ;
        RECT 2254.020 3342.380 2257.020 3342.390 ;
        RECT 2434.020 3342.380 2437.020 3342.390 ;
        RECT 2614.020 3342.380 2617.020 3342.390 ;
        RECT 2794.020 3342.380 2797.020 3342.390 ;
        RECT 2931.200 3342.380 2934.200 3342.390 ;
        RECT -14.580 3339.380 2934.200 3342.380 ;
        RECT -14.580 3339.370 -11.580 3339.380 ;
        RECT 94.020 3339.370 97.020 3339.380 ;
        RECT 274.020 3339.370 277.020 3339.380 ;
        RECT 454.020 3339.370 457.020 3339.380 ;
        RECT 634.020 3339.370 637.020 3339.380 ;
        RECT 814.020 3339.370 817.020 3339.380 ;
        RECT 994.020 3339.370 997.020 3339.380 ;
        RECT 1174.020 3339.370 1177.020 3339.380 ;
        RECT 1354.020 3339.370 1357.020 3339.380 ;
        RECT 1534.020 3339.370 1537.020 3339.380 ;
        RECT 1714.020 3339.370 1717.020 3339.380 ;
        RECT 1894.020 3339.370 1897.020 3339.380 ;
        RECT 2074.020 3339.370 2077.020 3339.380 ;
        RECT 2254.020 3339.370 2257.020 3339.380 ;
        RECT 2434.020 3339.370 2437.020 3339.380 ;
        RECT 2614.020 3339.370 2617.020 3339.380 ;
        RECT 2794.020 3339.370 2797.020 3339.380 ;
        RECT 2931.200 3339.370 2934.200 3339.380 ;
        RECT -14.580 3162.380 -11.580 3162.390 ;
        RECT 94.020 3162.380 97.020 3162.390 ;
        RECT 274.020 3162.380 277.020 3162.390 ;
        RECT 454.020 3162.380 457.020 3162.390 ;
        RECT 634.020 3162.380 637.020 3162.390 ;
        RECT 814.020 3162.380 817.020 3162.390 ;
        RECT 994.020 3162.380 997.020 3162.390 ;
        RECT 1174.020 3162.380 1177.020 3162.390 ;
        RECT 1354.020 3162.380 1357.020 3162.390 ;
        RECT 1534.020 3162.380 1537.020 3162.390 ;
        RECT 1714.020 3162.380 1717.020 3162.390 ;
        RECT 1894.020 3162.380 1897.020 3162.390 ;
        RECT 2074.020 3162.380 2077.020 3162.390 ;
        RECT 2254.020 3162.380 2257.020 3162.390 ;
        RECT 2434.020 3162.380 2437.020 3162.390 ;
        RECT 2614.020 3162.380 2617.020 3162.390 ;
        RECT 2794.020 3162.380 2797.020 3162.390 ;
        RECT 2931.200 3162.380 2934.200 3162.390 ;
        RECT -14.580 3159.380 2934.200 3162.380 ;
        RECT -14.580 3159.370 -11.580 3159.380 ;
        RECT 94.020 3159.370 97.020 3159.380 ;
        RECT 274.020 3159.370 277.020 3159.380 ;
        RECT 454.020 3159.370 457.020 3159.380 ;
        RECT 634.020 3159.370 637.020 3159.380 ;
        RECT 814.020 3159.370 817.020 3159.380 ;
        RECT 994.020 3159.370 997.020 3159.380 ;
        RECT 1174.020 3159.370 1177.020 3159.380 ;
        RECT 1354.020 3159.370 1357.020 3159.380 ;
        RECT 1534.020 3159.370 1537.020 3159.380 ;
        RECT 1714.020 3159.370 1717.020 3159.380 ;
        RECT 1894.020 3159.370 1897.020 3159.380 ;
        RECT 2074.020 3159.370 2077.020 3159.380 ;
        RECT 2254.020 3159.370 2257.020 3159.380 ;
        RECT 2434.020 3159.370 2437.020 3159.380 ;
        RECT 2614.020 3159.370 2617.020 3159.380 ;
        RECT 2794.020 3159.370 2797.020 3159.380 ;
        RECT 2931.200 3159.370 2934.200 3159.380 ;
        RECT -14.580 2982.380 -11.580 2982.390 ;
        RECT 94.020 2982.380 97.020 2982.390 ;
        RECT 274.020 2982.380 277.020 2982.390 ;
        RECT 454.020 2982.380 457.020 2982.390 ;
        RECT 634.020 2982.380 637.020 2982.390 ;
        RECT 814.020 2982.380 817.020 2982.390 ;
        RECT 994.020 2982.380 997.020 2982.390 ;
        RECT 1174.020 2982.380 1177.020 2982.390 ;
        RECT 1354.020 2982.380 1357.020 2982.390 ;
        RECT 1534.020 2982.380 1537.020 2982.390 ;
        RECT 1714.020 2982.380 1717.020 2982.390 ;
        RECT 1894.020 2982.380 1897.020 2982.390 ;
        RECT 2074.020 2982.380 2077.020 2982.390 ;
        RECT 2254.020 2982.380 2257.020 2982.390 ;
        RECT 2434.020 2982.380 2437.020 2982.390 ;
        RECT 2614.020 2982.380 2617.020 2982.390 ;
        RECT 2794.020 2982.380 2797.020 2982.390 ;
        RECT 2931.200 2982.380 2934.200 2982.390 ;
        RECT -14.580 2979.380 2934.200 2982.380 ;
        RECT -14.580 2979.370 -11.580 2979.380 ;
        RECT 94.020 2979.370 97.020 2979.380 ;
        RECT 274.020 2979.370 277.020 2979.380 ;
        RECT 454.020 2979.370 457.020 2979.380 ;
        RECT 634.020 2979.370 637.020 2979.380 ;
        RECT 814.020 2979.370 817.020 2979.380 ;
        RECT 994.020 2979.370 997.020 2979.380 ;
        RECT 1174.020 2979.370 1177.020 2979.380 ;
        RECT 1354.020 2979.370 1357.020 2979.380 ;
        RECT 1534.020 2979.370 1537.020 2979.380 ;
        RECT 1714.020 2979.370 1717.020 2979.380 ;
        RECT 1894.020 2979.370 1897.020 2979.380 ;
        RECT 2074.020 2979.370 2077.020 2979.380 ;
        RECT 2254.020 2979.370 2257.020 2979.380 ;
        RECT 2434.020 2979.370 2437.020 2979.380 ;
        RECT 2614.020 2979.370 2617.020 2979.380 ;
        RECT 2794.020 2979.370 2797.020 2979.380 ;
        RECT 2931.200 2979.370 2934.200 2979.380 ;
        RECT -14.580 2802.380 -11.580 2802.390 ;
        RECT 94.020 2802.380 97.020 2802.390 ;
        RECT 274.020 2802.380 277.020 2802.390 ;
        RECT 454.020 2802.380 457.020 2802.390 ;
        RECT 634.020 2802.380 637.020 2802.390 ;
        RECT 814.020 2802.380 817.020 2802.390 ;
        RECT 994.020 2802.380 997.020 2802.390 ;
        RECT 1174.020 2802.380 1177.020 2802.390 ;
        RECT 1354.020 2802.380 1357.020 2802.390 ;
        RECT 1534.020 2802.380 1537.020 2802.390 ;
        RECT 1714.020 2802.380 1717.020 2802.390 ;
        RECT 1894.020 2802.380 1897.020 2802.390 ;
        RECT 2074.020 2802.380 2077.020 2802.390 ;
        RECT 2254.020 2802.380 2257.020 2802.390 ;
        RECT 2434.020 2802.380 2437.020 2802.390 ;
        RECT 2614.020 2802.380 2617.020 2802.390 ;
        RECT 2794.020 2802.380 2797.020 2802.390 ;
        RECT 2931.200 2802.380 2934.200 2802.390 ;
        RECT -14.580 2799.380 2934.200 2802.380 ;
        RECT -14.580 2799.370 -11.580 2799.380 ;
        RECT 94.020 2799.370 97.020 2799.380 ;
        RECT 274.020 2799.370 277.020 2799.380 ;
        RECT 454.020 2799.370 457.020 2799.380 ;
        RECT 634.020 2799.370 637.020 2799.380 ;
        RECT 814.020 2799.370 817.020 2799.380 ;
        RECT 994.020 2799.370 997.020 2799.380 ;
        RECT 1174.020 2799.370 1177.020 2799.380 ;
        RECT 1354.020 2799.370 1357.020 2799.380 ;
        RECT 1534.020 2799.370 1537.020 2799.380 ;
        RECT 1714.020 2799.370 1717.020 2799.380 ;
        RECT 1894.020 2799.370 1897.020 2799.380 ;
        RECT 2074.020 2799.370 2077.020 2799.380 ;
        RECT 2254.020 2799.370 2257.020 2799.380 ;
        RECT 2434.020 2799.370 2437.020 2799.380 ;
        RECT 2614.020 2799.370 2617.020 2799.380 ;
        RECT 2794.020 2799.370 2797.020 2799.380 ;
        RECT 2931.200 2799.370 2934.200 2799.380 ;
        RECT -14.580 2622.380 -11.580 2622.390 ;
        RECT 94.020 2622.380 97.020 2622.390 ;
        RECT 274.020 2622.380 277.020 2622.390 ;
        RECT 454.020 2622.380 457.020 2622.390 ;
        RECT 634.020 2622.380 637.020 2622.390 ;
        RECT 814.020 2622.380 817.020 2622.390 ;
        RECT 994.020 2622.380 997.020 2622.390 ;
        RECT 1174.020 2622.380 1177.020 2622.390 ;
        RECT 1354.020 2622.380 1357.020 2622.390 ;
        RECT 1534.020 2622.380 1537.020 2622.390 ;
        RECT 1714.020 2622.380 1717.020 2622.390 ;
        RECT 1894.020 2622.380 1897.020 2622.390 ;
        RECT 2074.020 2622.380 2077.020 2622.390 ;
        RECT 2254.020 2622.380 2257.020 2622.390 ;
        RECT 2434.020 2622.380 2437.020 2622.390 ;
        RECT 2614.020 2622.380 2617.020 2622.390 ;
        RECT 2794.020 2622.380 2797.020 2622.390 ;
        RECT 2931.200 2622.380 2934.200 2622.390 ;
        RECT -14.580 2619.380 2934.200 2622.380 ;
        RECT -14.580 2619.370 -11.580 2619.380 ;
        RECT 94.020 2619.370 97.020 2619.380 ;
        RECT 274.020 2619.370 277.020 2619.380 ;
        RECT 454.020 2619.370 457.020 2619.380 ;
        RECT 634.020 2619.370 637.020 2619.380 ;
        RECT 814.020 2619.370 817.020 2619.380 ;
        RECT 994.020 2619.370 997.020 2619.380 ;
        RECT 1174.020 2619.370 1177.020 2619.380 ;
        RECT 1354.020 2619.370 1357.020 2619.380 ;
        RECT 1534.020 2619.370 1537.020 2619.380 ;
        RECT 1714.020 2619.370 1717.020 2619.380 ;
        RECT 1894.020 2619.370 1897.020 2619.380 ;
        RECT 2074.020 2619.370 2077.020 2619.380 ;
        RECT 2254.020 2619.370 2257.020 2619.380 ;
        RECT 2434.020 2619.370 2437.020 2619.380 ;
        RECT 2614.020 2619.370 2617.020 2619.380 ;
        RECT 2794.020 2619.370 2797.020 2619.380 ;
        RECT 2931.200 2619.370 2934.200 2619.380 ;
        RECT -14.580 2442.380 -11.580 2442.390 ;
        RECT 94.020 2442.380 97.020 2442.390 ;
        RECT 274.020 2442.380 277.020 2442.390 ;
        RECT 454.020 2442.380 457.020 2442.390 ;
        RECT 634.020 2442.380 637.020 2442.390 ;
        RECT 814.020 2442.380 817.020 2442.390 ;
        RECT 994.020 2442.380 997.020 2442.390 ;
        RECT 1174.020 2442.380 1177.020 2442.390 ;
        RECT 1354.020 2442.380 1357.020 2442.390 ;
        RECT 1534.020 2442.380 1537.020 2442.390 ;
        RECT 1714.020 2442.380 1717.020 2442.390 ;
        RECT 1894.020 2442.380 1897.020 2442.390 ;
        RECT 2074.020 2442.380 2077.020 2442.390 ;
        RECT 2254.020 2442.380 2257.020 2442.390 ;
        RECT 2434.020 2442.380 2437.020 2442.390 ;
        RECT 2614.020 2442.380 2617.020 2442.390 ;
        RECT 2794.020 2442.380 2797.020 2442.390 ;
        RECT 2931.200 2442.380 2934.200 2442.390 ;
        RECT -14.580 2439.380 2934.200 2442.380 ;
        RECT -14.580 2439.370 -11.580 2439.380 ;
        RECT 94.020 2439.370 97.020 2439.380 ;
        RECT 274.020 2439.370 277.020 2439.380 ;
        RECT 454.020 2439.370 457.020 2439.380 ;
        RECT 634.020 2439.370 637.020 2439.380 ;
        RECT 814.020 2439.370 817.020 2439.380 ;
        RECT 994.020 2439.370 997.020 2439.380 ;
        RECT 1174.020 2439.370 1177.020 2439.380 ;
        RECT 1354.020 2439.370 1357.020 2439.380 ;
        RECT 1534.020 2439.370 1537.020 2439.380 ;
        RECT 1714.020 2439.370 1717.020 2439.380 ;
        RECT 1894.020 2439.370 1897.020 2439.380 ;
        RECT 2074.020 2439.370 2077.020 2439.380 ;
        RECT 2254.020 2439.370 2257.020 2439.380 ;
        RECT 2434.020 2439.370 2437.020 2439.380 ;
        RECT 2614.020 2439.370 2617.020 2439.380 ;
        RECT 2794.020 2439.370 2797.020 2439.380 ;
        RECT 2931.200 2439.370 2934.200 2439.380 ;
        RECT -14.580 2262.380 -11.580 2262.390 ;
        RECT 94.020 2262.380 97.020 2262.390 ;
        RECT 274.020 2262.380 277.020 2262.390 ;
        RECT 454.020 2262.380 457.020 2262.390 ;
        RECT 634.020 2262.380 637.020 2262.390 ;
        RECT 814.020 2262.380 817.020 2262.390 ;
        RECT 994.020 2262.380 997.020 2262.390 ;
        RECT 1174.020 2262.380 1177.020 2262.390 ;
        RECT 1354.020 2262.380 1357.020 2262.390 ;
        RECT 1534.020 2262.380 1537.020 2262.390 ;
        RECT 1714.020 2262.380 1717.020 2262.390 ;
        RECT 1894.020 2262.380 1897.020 2262.390 ;
        RECT 2074.020 2262.380 2077.020 2262.390 ;
        RECT 2254.020 2262.380 2257.020 2262.390 ;
        RECT 2434.020 2262.380 2437.020 2262.390 ;
        RECT 2614.020 2262.380 2617.020 2262.390 ;
        RECT 2794.020 2262.380 2797.020 2262.390 ;
        RECT 2931.200 2262.380 2934.200 2262.390 ;
        RECT -14.580 2259.380 2934.200 2262.380 ;
        RECT -14.580 2259.370 -11.580 2259.380 ;
        RECT 94.020 2259.370 97.020 2259.380 ;
        RECT 274.020 2259.370 277.020 2259.380 ;
        RECT 454.020 2259.370 457.020 2259.380 ;
        RECT 634.020 2259.370 637.020 2259.380 ;
        RECT 814.020 2259.370 817.020 2259.380 ;
        RECT 994.020 2259.370 997.020 2259.380 ;
        RECT 1174.020 2259.370 1177.020 2259.380 ;
        RECT 1354.020 2259.370 1357.020 2259.380 ;
        RECT 1534.020 2259.370 1537.020 2259.380 ;
        RECT 1714.020 2259.370 1717.020 2259.380 ;
        RECT 1894.020 2259.370 1897.020 2259.380 ;
        RECT 2074.020 2259.370 2077.020 2259.380 ;
        RECT 2254.020 2259.370 2257.020 2259.380 ;
        RECT 2434.020 2259.370 2437.020 2259.380 ;
        RECT 2614.020 2259.370 2617.020 2259.380 ;
        RECT 2794.020 2259.370 2797.020 2259.380 ;
        RECT 2931.200 2259.370 2934.200 2259.380 ;
        RECT -14.580 2082.380 -11.580 2082.390 ;
        RECT 94.020 2082.380 97.020 2082.390 ;
        RECT 274.020 2082.380 277.020 2082.390 ;
        RECT 454.020 2082.380 457.020 2082.390 ;
        RECT 634.020 2082.380 637.020 2082.390 ;
        RECT 814.020 2082.380 817.020 2082.390 ;
        RECT 994.020 2082.380 997.020 2082.390 ;
        RECT 1174.020 2082.380 1177.020 2082.390 ;
        RECT 1354.020 2082.380 1357.020 2082.390 ;
        RECT 1534.020 2082.380 1537.020 2082.390 ;
        RECT 1714.020 2082.380 1717.020 2082.390 ;
        RECT 1894.020 2082.380 1897.020 2082.390 ;
        RECT 2074.020 2082.380 2077.020 2082.390 ;
        RECT 2254.020 2082.380 2257.020 2082.390 ;
        RECT 2434.020 2082.380 2437.020 2082.390 ;
        RECT 2614.020 2082.380 2617.020 2082.390 ;
        RECT 2794.020 2082.380 2797.020 2082.390 ;
        RECT 2931.200 2082.380 2934.200 2082.390 ;
        RECT -14.580 2079.380 2934.200 2082.380 ;
        RECT -14.580 2079.370 -11.580 2079.380 ;
        RECT 94.020 2079.370 97.020 2079.380 ;
        RECT 274.020 2079.370 277.020 2079.380 ;
        RECT 454.020 2079.370 457.020 2079.380 ;
        RECT 634.020 2079.370 637.020 2079.380 ;
        RECT 814.020 2079.370 817.020 2079.380 ;
        RECT 994.020 2079.370 997.020 2079.380 ;
        RECT 1174.020 2079.370 1177.020 2079.380 ;
        RECT 1354.020 2079.370 1357.020 2079.380 ;
        RECT 1534.020 2079.370 1537.020 2079.380 ;
        RECT 1714.020 2079.370 1717.020 2079.380 ;
        RECT 1894.020 2079.370 1897.020 2079.380 ;
        RECT 2074.020 2079.370 2077.020 2079.380 ;
        RECT 2254.020 2079.370 2257.020 2079.380 ;
        RECT 2434.020 2079.370 2437.020 2079.380 ;
        RECT 2614.020 2079.370 2617.020 2079.380 ;
        RECT 2794.020 2079.370 2797.020 2079.380 ;
        RECT 2931.200 2079.370 2934.200 2079.380 ;
        RECT -14.580 1902.380 -11.580 1902.390 ;
        RECT 94.020 1902.380 97.020 1902.390 ;
        RECT 274.020 1902.380 277.020 1902.390 ;
        RECT 454.020 1902.380 457.020 1902.390 ;
        RECT 634.020 1902.380 637.020 1902.390 ;
        RECT 814.020 1902.380 817.020 1902.390 ;
        RECT 994.020 1902.380 997.020 1902.390 ;
        RECT 1174.020 1902.380 1177.020 1902.390 ;
        RECT 1354.020 1902.380 1357.020 1902.390 ;
        RECT 1534.020 1902.380 1537.020 1902.390 ;
        RECT 1714.020 1902.380 1717.020 1902.390 ;
        RECT 1894.020 1902.380 1897.020 1902.390 ;
        RECT 2074.020 1902.380 2077.020 1902.390 ;
        RECT 2254.020 1902.380 2257.020 1902.390 ;
        RECT 2434.020 1902.380 2437.020 1902.390 ;
        RECT 2614.020 1902.380 2617.020 1902.390 ;
        RECT 2794.020 1902.380 2797.020 1902.390 ;
        RECT 2931.200 1902.380 2934.200 1902.390 ;
        RECT -14.580 1899.380 2934.200 1902.380 ;
        RECT -14.580 1899.370 -11.580 1899.380 ;
        RECT 94.020 1899.370 97.020 1899.380 ;
        RECT 274.020 1899.370 277.020 1899.380 ;
        RECT 454.020 1899.370 457.020 1899.380 ;
        RECT 634.020 1899.370 637.020 1899.380 ;
        RECT 814.020 1899.370 817.020 1899.380 ;
        RECT 994.020 1899.370 997.020 1899.380 ;
        RECT 1174.020 1899.370 1177.020 1899.380 ;
        RECT 1354.020 1899.370 1357.020 1899.380 ;
        RECT 1534.020 1899.370 1537.020 1899.380 ;
        RECT 1714.020 1899.370 1717.020 1899.380 ;
        RECT 1894.020 1899.370 1897.020 1899.380 ;
        RECT 2074.020 1899.370 2077.020 1899.380 ;
        RECT 2254.020 1899.370 2257.020 1899.380 ;
        RECT 2434.020 1899.370 2437.020 1899.380 ;
        RECT 2614.020 1899.370 2617.020 1899.380 ;
        RECT 2794.020 1899.370 2797.020 1899.380 ;
        RECT 2931.200 1899.370 2934.200 1899.380 ;
        RECT -14.580 1722.380 -11.580 1722.390 ;
        RECT 94.020 1722.380 97.020 1722.390 ;
        RECT 274.020 1722.380 277.020 1722.390 ;
        RECT 454.020 1722.380 457.020 1722.390 ;
        RECT 634.020 1722.380 637.020 1722.390 ;
        RECT 814.020 1722.380 817.020 1722.390 ;
        RECT 994.020 1722.380 997.020 1722.390 ;
        RECT 1174.020 1722.380 1177.020 1722.390 ;
        RECT 1354.020 1722.380 1357.020 1722.390 ;
        RECT 1534.020 1722.380 1537.020 1722.390 ;
        RECT 1714.020 1722.380 1717.020 1722.390 ;
        RECT 1894.020 1722.380 1897.020 1722.390 ;
        RECT 2074.020 1722.380 2077.020 1722.390 ;
        RECT 2254.020 1722.380 2257.020 1722.390 ;
        RECT 2434.020 1722.380 2437.020 1722.390 ;
        RECT 2614.020 1722.380 2617.020 1722.390 ;
        RECT 2794.020 1722.380 2797.020 1722.390 ;
        RECT 2931.200 1722.380 2934.200 1722.390 ;
        RECT -14.580 1719.380 2934.200 1722.380 ;
        RECT -14.580 1719.370 -11.580 1719.380 ;
        RECT 94.020 1719.370 97.020 1719.380 ;
        RECT 274.020 1719.370 277.020 1719.380 ;
        RECT 454.020 1719.370 457.020 1719.380 ;
        RECT 634.020 1719.370 637.020 1719.380 ;
        RECT 814.020 1719.370 817.020 1719.380 ;
        RECT 994.020 1719.370 997.020 1719.380 ;
        RECT 1174.020 1719.370 1177.020 1719.380 ;
        RECT 1354.020 1719.370 1357.020 1719.380 ;
        RECT 1534.020 1719.370 1537.020 1719.380 ;
        RECT 1714.020 1719.370 1717.020 1719.380 ;
        RECT 1894.020 1719.370 1897.020 1719.380 ;
        RECT 2074.020 1719.370 2077.020 1719.380 ;
        RECT 2254.020 1719.370 2257.020 1719.380 ;
        RECT 2434.020 1719.370 2437.020 1719.380 ;
        RECT 2614.020 1719.370 2617.020 1719.380 ;
        RECT 2794.020 1719.370 2797.020 1719.380 ;
        RECT 2931.200 1719.370 2934.200 1719.380 ;
        RECT -14.580 1542.380 -11.580 1542.390 ;
        RECT 94.020 1542.380 97.020 1542.390 ;
        RECT 274.020 1542.380 277.020 1542.390 ;
        RECT 454.020 1542.380 457.020 1542.390 ;
        RECT 634.020 1542.380 637.020 1542.390 ;
        RECT 814.020 1542.380 817.020 1542.390 ;
        RECT 994.020 1542.380 997.020 1542.390 ;
        RECT 1174.020 1542.380 1177.020 1542.390 ;
        RECT 1354.020 1542.380 1357.020 1542.390 ;
        RECT 1534.020 1542.380 1537.020 1542.390 ;
        RECT 1714.020 1542.380 1717.020 1542.390 ;
        RECT 1894.020 1542.380 1897.020 1542.390 ;
        RECT 2074.020 1542.380 2077.020 1542.390 ;
        RECT 2254.020 1542.380 2257.020 1542.390 ;
        RECT 2434.020 1542.380 2437.020 1542.390 ;
        RECT 2614.020 1542.380 2617.020 1542.390 ;
        RECT 2794.020 1542.380 2797.020 1542.390 ;
        RECT 2931.200 1542.380 2934.200 1542.390 ;
        RECT -14.580 1539.380 2934.200 1542.380 ;
        RECT -14.580 1539.370 -11.580 1539.380 ;
        RECT 94.020 1539.370 97.020 1539.380 ;
        RECT 274.020 1539.370 277.020 1539.380 ;
        RECT 454.020 1539.370 457.020 1539.380 ;
        RECT 634.020 1539.370 637.020 1539.380 ;
        RECT 814.020 1539.370 817.020 1539.380 ;
        RECT 994.020 1539.370 997.020 1539.380 ;
        RECT 1174.020 1539.370 1177.020 1539.380 ;
        RECT 1354.020 1539.370 1357.020 1539.380 ;
        RECT 1534.020 1539.370 1537.020 1539.380 ;
        RECT 1714.020 1539.370 1717.020 1539.380 ;
        RECT 1894.020 1539.370 1897.020 1539.380 ;
        RECT 2074.020 1539.370 2077.020 1539.380 ;
        RECT 2254.020 1539.370 2257.020 1539.380 ;
        RECT 2434.020 1539.370 2437.020 1539.380 ;
        RECT 2614.020 1539.370 2617.020 1539.380 ;
        RECT 2794.020 1539.370 2797.020 1539.380 ;
        RECT 2931.200 1539.370 2934.200 1539.380 ;
        RECT -14.580 1362.380 -11.580 1362.390 ;
        RECT 94.020 1362.380 97.020 1362.390 ;
        RECT 274.020 1362.380 277.020 1362.390 ;
        RECT 454.020 1362.380 457.020 1362.390 ;
        RECT 634.020 1362.380 637.020 1362.390 ;
        RECT 814.020 1362.380 817.020 1362.390 ;
        RECT 994.020 1362.380 997.020 1362.390 ;
        RECT 1174.020 1362.380 1177.020 1362.390 ;
        RECT 1354.020 1362.380 1357.020 1362.390 ;
        RECT 1534.020 1362.380 1537.020 1362.390 ;
        RECT 1714.020 1362.380 1717.020 1362.390 ;
        RECT 1894.020 1362.380 1897.020 1362.390 ;
        RECT 2074.020 1362.380 2077.020 1362.390 ;
        RECT 2254.020 1362.380 2257.020 1362.390 ;
        RECT 2434.020 1362.380 2437.020 1362.390 ;
        RECT 2614.020 1362.380 2617.020 1362.390 ;
        RECT 2794.020 1362.380 2797.020 1362.390 ;
        RECT 2931.200 1362.380 2934.200 1362.390 ;
        RECT -14.580 1359.380 2934.200 1362.380 ;
        RECT -14.580 1359.370 -11.580 1359.380 ;
        RECT 94.020 1359.370 97.020 1359.380 ;
        RECT 274.020 1359.370 277.020 1359.380 ;
        RECT 454.020 1359.370 457.020 1359.380 ;
        RECT 634.020 1359.370 637.020 1359.380 ;
        RECT 814.020 1359.370 817.020 1359.380 ;
        RECT 994.020 1359.370 997.020 1359.380 ;
        RECT 1174.020 1359.370 1177.020 1359.380 ;
        RECT 1354.020 1359.370 1357.020 1359.380 ;
        RECT 1534.020 1359.370 1537.020 1359.380 ;
        RECT 1714.020 1359.370 1717.020 1359.380 ;
        RECT 1894.020 1359.370 1897.020 1359.380 ;
        RECT 2074.020 1359.370 2077.020 1359.380 ;
        RECT 2254.020 1359.370 2257.020 1359.380 ;
        RECT 2434.020 1359.370 2437.020 1359.380 ;
        RECT 2614.020 1359.370 2617.020 1359.380 ;
        RECT 2794.020 1359.370 2797.020 1359.380 ;
        RECT 2931.200 1359.370 2934.200 1359.380 ;
        RECT -14.580 1182.380 -11.580 1182.390 ;
        RECT 94.020 1182.380 97.020 1182.390 ;
        RECT 274.020 1182.380 277.020 1182.390 ;
        RECT 454.020 1182.380 457.020 1182.390 ;
        RECT 634.020 1182.380 637.020 1182.390 ;
        RECT 814.020 1182.380 817.020 1182.390 ;
        RECT 994.020 1182.380 997.020 1182.390 ;
        RECT 1174.020 1182.380 1177.020 1182.390 ;
        RECT 1354.020 1182.380 1357.020 1182.390 ;
        RECT 1534.020 1182.380 1537.020 1182.390 ;
        RECT 1714.020 1182.380 1717.020 1182.390 ;
        RECT 1894.020 1182.380 1897.020 1182.390 ;
        RECT 2074.020 1182.380 2077.020 1182.390 ;
        RECT 2254.020 1182.380 2257.020 1182.390 ;
        RECT 2434.020 1182.380 2437.020 1182.390 ;
        RECT 2614.020 1182.380 2617.020 1182.390 ;
        RECT 2794.020 1182.380 2797.020 1182.390 ;
        RECT 2931.200 1182.380 2934.200 1182.390 ;
        RECT -14.580 1179.380 2934.200 1182.380 ;
        RECT -14.580 1179.370 -11.580 1179.380 ;
        RECT 94.020 1179.370 97.020 1179.380 ;
        RECT 274.020 1179.370 277.020 1179.380 ;
        RECT 454.020 1179.370 457.020 1179.380 ;
        RECT 634.020 1179.370 637.020 1179.380 ;
        RECT 814.020 1179.370 817.020 1179.380 ;
        RECT 994.020 1179.370 997.020 1179.380 ;
        RECT 1174.020 1179.370 1177.020 1179.380 ;
        RECT 1354.020 1179.370 1357.020 1179.380 ;
        RECT 1534.020 1179.370 1537.020 1179.380 ;
        RECT 1714.020 1179.370 1717.020 1179.380 ;
        RECT 1894.020 1179.370 1897.020 1179.380 ;
        RECT 2074.020 1179.370 2077.020 1179.380 ;
        RECT 2254.020 1179.370 2257.020 1179.380 ;
        RECT 2434.020 1179.370 2437.020 1179.380 ;
        RECT 2614.020 1179.370 2617.020 1179.380 ;
        RECT 2794.020 1179.370 2797.020 1179.380 ;
        RECT 2931.200 1179.370 2934.200 1179.380 ;
        RECT -14.580 1002.380 -11.580 1002.390 ;
        RECT 94.020 1002.380 97.020 1002.390 ;
        RECT 274.020 1002.380 277.020 1002.390 ;
        RECT 454.020 1002.380 457.020 1002.390 ;
        RECT 634.020 1002.380 637.020 1002.390 ;
        RECT 814.020 1002.380 817.020 1002.390 ;
        RECT 994.020 1002.380 997.020 1002.390 ;
        RECT 1174.020 1002.380 1177.020 1002.390 ;
        RECT 1354.020 1002.380 1357.020 1002.390 ;
        RECT 1534.020 1002.380 1537.020 1002.390 ;
        RECT 1714.020 1002.380 1717.020 1002.390 ;
        RECT 1894.020 1002.380 1897.020 1002.390 ;
        RECT 2074.020 1002.380 2077.020 1002.390 ;
        RECT 2254.020 1002.380 2257.020 1002.390 ;
        RECT 2434.020 1002.380 2437.020 1002.390 ;
        RECT 2614.020 1002.380 2617.020 1002.390 ;
        RECT 2794.020 1002.380 2797.020 1002.390 ;
        RECT 2931.200 1002.380 2934.200 1002.390 ;
        RECT -14.580 999.380 2934.200 1002.380 ;
        RECT -14.580 999.370 -11.580 999.380 ;
        RECT 94.020 999.370 97.020 999.380 ;
        RECT 274.020 999.370 277.020 999.380 ;
        RECT 454.020 999.370 457.020 999.380 ;
        RECT 634.020 999.370 637.020 999.380 ;
        RECT 814.020 999.370 817.020 999.380 ;
        RECT 994.020 999.370 997.020 999.380 ;
        RECT 1174.020 999.370 1177.020 999.380 ;
        RECT 1354.020 999.370 1357.020 999.380 ;
        RECT 1534.020 999.370 1537.020 999.380 ;
        RECT 1714.020 999.370 1717.020 999.380 ;
        RECT 1894.020 999.370 1897.020 999.380 ;
        RECT 2074.020 999.370 2077.020 999.380 ;
        RECT 2254.020 999.370 2257.020 999.380 ;
        RECT 2434.020 999.370 2437.020 999.380 ;
        RECT 2614.020 999.370 2617.020 999.380 ;
        RECT 2794.020 999.370 2797.020 999.380 ;
        RECT 2931.200 999.370 2934.200 999.380 ;
        RECT -14.580 822.380 -11.580 822.390 ;
        RECT 94.020 822.380 97.020 822.390 ;
        RECT 274.020 822.380 277.020 822.390 ;
        RECT 454.020 822.380 457.020 822.390 ;
        RECT 634.020 822.380 637.020 822.390 ;
        RECT 814.020 822.380 817.020 822.390 ;
        RECT 994.020 822.380 997.020 822.390 ;
        RECT 1174.020 822.380 1177.020 822.390 ;
        RECT 1354.020 822.380 1357.020 822.390 ;
        RECT 1534.020 822.380 1537.020 822.390 ;
        RECT 1714.020 822.380 1717.020 822.390 ;
        RECT 1894.020 822.380 1897.020 822.390 ;
        RECT 2074.020 822.380 2077.020 822.390 ;
        RECT 2254.020 822.380 2257.020 822.390 ;
        RECT 2434.020 822.380 2437.020 822.390 ;
        RECT 2614.020 822.380 2617.020 822.390 ;
        RECT 2794.020 822.380 2797.020 822.390 ;
        RECT 2931.200 822.380 2934.200 822.390 ;
        RECT -14.580 819.380 2934.200 822.380 ;
        RECT -14.580 819.370 -11.580 819.380 ;
        RECT 94.020 819.370 97.020 819.380 ;
        RECT 274.020 819.370 277.020 819.380 ;
        RECT 454.020 819.370 457.020 819.380 ;
        RECT 634.020 819.370 637.020 819.380 ;
        RECT 814.020 819.370 817.020 819.380 ;
        RECT 994.020 819.370 997.020 819.380 ;
        RECT 1174.020 819.370 1177.020 819.380 ;
        RECT 1354.020 819.370 1357.020 819.380 ;
        RECT 1534.020 819.370 1537.020 819.380 ;
        RECT 1714.020 819.370 1717.020 819.380 ;
        RECT 1894.020 819.370 1897.020 819.380 ;
        RECT 2074.020 819.370 2077.020 819.380 ;
        RECT 2254.020 819.370 2257.020 819.380 ;
        RECT 2434.020 819.370 2437.020 819.380 ;
        RECT 2614.020 819.370 2617.020 819.380 ;
        RECT 2794.020 819.370 2797.020 819.380 ;
        RECT 2931.200 819.370 2934.200 819.380 ;
        RECT -14.580 642.380 -11.580 642.390 ;
        RECT 94.020 642.380 97.020 642.390 ;
        RECT 274.020 642.380 277.020 642.390 ;
        RECT 454.020 642.380 457.020 642.390 ;
        RECT 634.020 642.380 637.020 642.390 ;
        RECT 814.020 642.380 817.020 642.390 ;
        RECT 994.020 642.380 997.020 642.390 ;
        RECT 1174.020 642.380 1177.020 642.390 ;
        RECT 1354.020 642.380 1357.020 642.390 ;
        RECT 1534.020 642.380 1537.020 642.390 ;
        RECT 1714.020 642.380 1717.020 642.390 ;
        RECT 1894.020 642.380 1897.020 642.390 ;
        RECT 2074.020 642.380 2077.020 642.390 ;
        RECT 2254.020 642.380 2257.020 642.390 ;
        RECT 2434.020 642.380 2437.020 642.390 ;
        RECT 2614.020 642.380 2617.020 642.390 ;
        RECT 2794.020 642.380 2797.020 642.390 ;
        RECT 2931.200 642.380 2934.200 642.390 ;
        RECT -14.580 639.380 2934.200 642.380 ;
        RECT -14.580 639.370 -11.580 639.380 ;
        RECT 94.020 639.370 97.020 639.380 ;
        RECT 274.020 639.370 277.020 639.380 ;
        RECT 454.020 639.370 457.020 639.380 ;
        RECT 634.020 639.370 637.020 639.380 ;
        RECT 814.020 639.370 817.020 639.380 ;
        RECT 994.020 639.370 997.020 639.380 ;
        RECT 1174.020 639.370 1177.020 639.380 ;
        RECT 1354.020 639.370 1357.020 639.380 ;
        RECT 1534.020 639.370 1537.020 639.380 ;
        RECT 1714.020 639.370 1717.020 639.380 ;
        RECT 1894.020 639.370 1897.020 639.380 ;
        RECT 2074.020 639.370 2077.020 639.380 ;
        RECT 2254.020 639.370 2257.020 639.380 ;
        RECT 2434.020 639.370 2437.020 639.380 ;
        RECT 2614.020 639.370 2617.020 639.380 ;
        RECT 2794.020 639.370 2797.020 639.380 ;
        RECT 2931.200 639.370 2934.200 639.380 ;
        RECT -14.580 462.380 -11.580 462.390 ;
        RECT 94.020 462.380 97.020 462.390 ;
        RECT 274.020 462.380 277.020 462.390 ;
        RECT 454.020 462.380 457.020 462.390 ;
        RECT 634.020 462.380 637.020 462.390 ;
        RECT 814.020 462.380 817.020 462.390 ;
        RECT 994.020 462.380 997.020 462.390 ;
        RECT 1174.020 462.380 1177.020 462.390 ;
        RECT 1354.020 462.380 1357.020 462.390 ;
        RECT 1534.020 462.380 1537.020 462.390 ;
        RECT 1714.020 462.380 1717.020 462.390 ;
        RECT 1894.020 462.380 1897.020 462.390 ;
        RECT 2074.020 462.380 2077.020 462.390 ;
        RECT 2254.020 462.380 2257.020 462.390 ;
        RECT 2434.020 462.380 2437.020 462.390 ;
        RECT 2614.020 462.380 2617.020 462.390 ;
        RECT 2794.020 462.380 2797.020 462.390 ;
        RECT 2931.200 462.380 2934.200 462.390 ;
        RECT -14.580 459.380 2934.200 462.380 ;
        RECT -14.580 459.370 -11.580 459.380 ;
        RECT 94.020 459.370 97.020 459.380 ;
        RECT 274.020 459.370 277.020 459.380 ;
        RECT 454.020 459.370 457.020 459.380 ;
        RECT 634.020 459.370 637.020 459.380 ;
        RECT 814.020 459.370 817.020 459.380 ;
        RECT 994.020 459.370 997.020 459.380 ;
        RECT 1174.020 459.370 1177.020 459.380 ;
        RECT 1354.020 459.370 1357.020 459.380 ;
        RECT 1534.020 459.370 1537.020 459.380 ;
        RECT 1714.020 459.370 1717.020 459.380 ;
        RECT 1894.020 459.370 1897.020 459.380 ;
        RECT 2074.020 459.370 2077.020 459.380 ;
        RECT 2254.020 459.370 2257.020 459.380 ;
        RECT 2434.020 459.370 2437.020 459.380 ;
        RECT 2614.020 459.370 2617.020 459.380 ;
        RECT 2794.020 459.370 2797.020 459.380 ;
        RECT 2931.200 459.370 2934.200 459.380 ;
        RECT -14.580 282.380 -11.580 282.390 ;
        RECT 94.020 282.380 97.020 282.390 ;
        RECT 274.020 282.380 277.020 282.390 ;
        RECT 454.020 282.380 457.020 282.390 ;
        RECT 634.020 282.380 637.020 282.390 ;
        RECT 814.020 282.380 817.020 282.390 ;
        RECT 994.020 282.380 997.020 282.390 ;
        RECT 1174.020 282.380 1177.020 282.390 ;
        RECT 1354.020 282.380 1357.020 282.390 ;
        RECT 1534.020 282.380 1537.020 282.390 ;
        RECT 1714.020 282.380 1717.020 282.390 ;
        RECT 1894.020 282.380 1897.020 282.390 ;
        RECT 2074.020 282.380 2077.020 282.390 ;
        RECT 2254.020 282.380 2257.020 282.390 ;
        RECT 2434.020 282.380 2437.020 282.390 ;
        RECT 2614.020 282.380 2617.020 282.390 ;
        RECT 2794.020 282.380 2797.020 282.390 ;
        RECT 2931.200 282.380 2934.200 282.390 ;
        RECT -14.580 279.380 2934.200 282.380 ;
        RECT -14.580 279.370 -11.580 279.380 ;
        RECT 94.020 279.370 97.020 279.380 ;
        RECT 274.020 279.370 277.020 279.380 ;
        RECT 454.020 279.370 457.020 279.380 ;
        RECT 634.020 279.370 637.020 279.380 ;
        RECT 814.020 279.370 817.020 279.380 ;
        RECT 994.020 279.370 997.020 279.380 ;
        RECT 1174.020 279.370 1177.020 279.380 ;
        RECT 1354.020 279.370 1357.020 279.380 ;
        RECT 1534.020 279.370 1537.020 279.380 ;
        RECT 1714.020 279.370 1717.020 279.380 ;
        RECT 1894.020 279.370 1897.020 279.380 ;
        RECT 2074.020 279.370 2077.020 279.380 ;
        RECT 2254.020 279.370 2257.020 279.380 ;
        RECT 2434.020 279.370 2437.020 279.380 ;
        RECT 2614.020 279.370 2617.020 279.380 ;
        RECT 2794.020 279.370 2797.020 279.380 ;
        RECT 2931.200 279.370 2934.200 279.380 ;
        RECT -14.580 102.380 -11.580 102.390 ;
        RECT 94.020 102.380 97.020 102.390 ;
        RECT 274.020 102.380 277.020 102.390 ;
        RECT 454.020 102.380 457.020 102.390 ;
        RECT 634.020 102.380 637.020 102.390 ;
        RECT 814.020 102.380 817.020 102.390 ;
        RECT 994.020 102.380 997.020 102.390 ;
        RECT 1174.020 102.380 1177.020 102.390 ;
        RECT 1354.020 102.380 1357.020 102.390 ;
        RECT 1534.020 102.380 1537.020 102.390 ;
        RECT 1714.020 102.380 1717.020 102.390 ;
        RECT 1894.020 102.380 1897.020 102.390 ;
        RECT 2074.020 102.380 2077.020 102.390 ;
        RECT 2254.020 102.380 2257.020 102.390 ;
        RECT 2434.020 102.380 2437.020 102.390 ;
        RECT 2614.020 102.380 2617.020 102.390 ;
        RECT 2794.020 102.380 2797.020 102.390 ;
        RECT 2931.200 102.380 2934.200 102.390 ;
        RECT -14.580 99.380 2934.200 102.380 ;
        RECT -14.580 99.370 -11.580 99.380 ;
        RECT 94.020 99.370 97.020 99.380 ;
        RECT 274.020 99.370 277.020 99.380 ;
        RECT 454.020 99.370 457.020 99.380 ;
        RECT 634.020 99.370 637.020 99.380 ;
        RECT 814.020 99.370 817.020 99.380 ;
        RECT 994.020 99.370 997.020 99.380 ;
        RECT 1174.020 99.370 1177.020 99.380 ;
        RECT 1354.020 99.370 1357.020 99.380 ;
        RECT 1534.020 99.370 1537.020 99.380 ;
        RECT 1714.020 99.370 1717.020 99.380 ;
        RECT 1894.020 99.370 1897.020 99.380 ;
        RECT 2074.020 99.370 2077.020 99.380 ;
        RECT 2254.020 99.370 2257.020 99.380 ;
        RECT 2434.020 99.370 2437.020 99.380 ;
        RECT 2614.020 99.370 2617.020 99.380 ;
        RECT 2794.020 99.370 2797.020 99.380 ;
        RECT 2931.200 99.370 2934.200 99.380 ;
        RECT -14.580 -6.220 -11.580 -6.210 ;
        RECT 94.020 -6.220 97.020 -6.210 ;
        RECT 274.020 -6.220 277.020 -6.210 ;
        RECT 454.020 -6.220 457.020 -6.210 ;
        RECT 634.020 -6.220 637.020 -6.210 ;
        RECT 814.020 -6.220 817.020 -6.210 ;
        RECT 994.020 -6.220 997.020 -6.210 ;
        RECT 1174.020 -6.220 1177.020 -6.210 ;
        RECT 1354.020 -6.220 1357.020 -6.210 ;
        RECT 1534.020 -6.220 1537.020 -6.210 ;
        RECT 1714.020 -6.220 1717.020 -6.210 ;
        RECT 1894.020 -6.220 1897.020 -6.210 ;
        RECT 2074.020 -6.220 2077.020 -6.210 ;
        RECT 2254.020 -6.220 2257.020 -6.210 ;
        RECT 2434.020 -6.220 2437.020 -6.210 ;
        RECT 2614.020 -6.220 2617.020 -6.210 ;
        RECT 2794.020 -6.220 2797.020 -6.210 ;
        RECT 2931.200 -6.220 2934.200 -6.210 ;
        RECT -14.580 -9.220 2934.200 -6.220 ;
        RECT -14.580 -9.230 -11.580 -9.220 ;
        RECT 94.020 -9.230 97.020 -9.220 ;
        RECT 274.020 -9.230 277.020 -9.220 ;
        RECT 454.020 -9.230 457.020 -9.220 ;
        RECT 634.020 -9.230 637.020 -9.220 ;
        RECT 814.020 -9.230 817.020 -9.220 ;
        RECT 994.020 -9.230 997.020 -9.220 ;
        RECT 1174.020 -9.230 1177.020 -9.220 ;
        RECT 1354.020 -9.230 1357.020 -9.220 ;
        RECT 1534.020 -9.230 1537.020 -9.220 ;
        RECT 1714.020 -9.230 1717.020 -9.220 ;
        RECT 1894.020 -9.230 1897.020 -9.220 ;
        RECT 2074.020 -9.230 2077.020 -9.220 ;
        RECT 2254.020 -9.230 2257.020 -9.220 ;
        RECT 2434.020 -9.230 2437.020 -9.220 ;
        RECT 2614.020 -9.230 2617.020 -9.220 ;
        RECT 2794.020 -9.230 2797.020 -9.220 ;
        RECT 2931.200 -9.230 2934.200 -9.220 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -19.180 -13.820 -16.180 3533.500 ;
        RECT 22.020 -18.420 25.020 3538.100 ;
        RECT 202.020 -18.420 205.020 3538.100 ;
        RECT 382.020 -18.420 385.020 3538.100 ;
        RECT 562.020 -18.420 565.020 3538.100 ;
        RECT 742.020 -18.420 745.020 3538.100 ;
        RECT 922.020 -18.420 925.020 3538.100 ;
        RECT 1102.020 -18.420 1105.020 3538.100 ;
        RECT 1282.020 -18.420 1285.020 3538.100 ;
        RECT 1462.020 -18.420 1465.020 3538.100 ;
        RECT 1642.020 -18.420 1645.020 3538.100 ;
        RECT 1822.020 -18.420 1825.020 3538.100 ;
        RECT 2002.020 -18.420 2005.020 3538.100 ;
        RECT 2182.020 -18.420 2185.020 3538.100 ;
        RECT 2362.020 -18.420 2365.020 3538.100 ;
        RECT 2542.020 -18.420 2545.020 3538.100 ;
        RECT 2722.020 -18.420 2725.020 3538.100 ;
        RECT 2902.020 -18.420 2905.020 3538.100 ;
        RECT 2935.800 -13.820 2938.800 3533.500 ;
      LAYER via4 ;
        RECT -18.270 3532.210 -17.090 3533.390 ;
        RECT -18.270 3530.610 -17.090 3531.790 ;
        RECT -18.270 3449.090 -17.090 3450.270 ;
        RECT -18.270 3447.490 -17.090 3448.670 ;
        RECT -18.270 3269.090 -17.090 3270.270 ;
        RECT -18.270 3267.490 -17.090 3268.670 ;
        RECT -18.270 3089.090 -17.090 3090.270 ;
        RECT -18.270 3087.490 -17.090 3088.670 ;
        RECT -18.270 2909.090 -17.090 2910.270 ;
        RECT -18.270 2907.490 -17.090 2908.670 ;
        RECT -18.270 2729.090 -17.090 2730.270 ;
        RECT -18.270 2727.490 -17.090 2728.670 ;
        RECT -18.270 2549.090 -17.090 2550.270 ;
        RECT -18.270 2547.490 -17.090 2548.670 ;
        RECT -18.270 2369.090 -17.090 2370.270 ;
        RECT -18.270 2367.490 -17.090 2368.670 ;
        RECT -18.270 2189.090 -17.090 2190.270 ;
        RECT -18.270 2187.490 -17.090 2188.670 ;
        RECT -18.270 2009.090 -17.090 2010.270 ;
        RECT -18.270 2007.490 -17.090 2008.670 ;
        RECT -18.270 1829.090 -17.090 1830.270 ;
        RECT -18.270 1827.490 -17.090 1828.670 ;
        RECT -18.270 1649.090 -17.090 1650.270 ;
        RECT -18.270 1647.490 -17.090 1648.670 ;
        RECT -18.270 1469.090 -17.090 1470.270 ;
        RECT -18.270 1467.490 -17.090 1468.670 ;
        RECT -18.270 1289.090 -17.090 1290.270 ;
        RECT -18.270 1287.490 -17.090 1288.670 ;
        RECT -18.270 1109.090 -17.090 1110.270 ;
        RECT -18.270 1107.490 -17.090 1108.670 ;
        RECT -18.270 929.090 -17.090 930.270 ;
        RECT -18.270 927.490 -17.090 928.670 ;
        RECT -18.270 749.090 -17.090 750.270 ;
        RECT -18.270 747.490 -17.090 748.670 ;
        RECT -18.270 569.090 -17.090 570.270 ;
        RECT -18.270 567.490 -17.090 568.670 ;
        RECT -18.270 389.090 -17.090 390.270 ;
        RECT -18.270 387.490 -17.090 388.670 ;
        RECT -18.270 209.090 -17.090 210.270 ;
        RECT -18.270 207.490 -17.090 208.670 ;
        RECT -18.270 29.090 -17.090 30.270 ;
        RECT -18.270 27.490 -17.090 28.670 ;
        RECT -18.270 -12.110 -17.090 -10.930 ;
        RECT -18.270 -13.710 -17.090 -12.530 ;
        RECT 22.930 3532.210 24.110 3533.390 ;
        RECT 22.930 3530.610 24.110 3531.790 ;
        RECT 22.930 3449.090 24.110 3450.270 ;
        RECT 22.930 3447.490 24.110 3448.670 ;
        RECT 22.930 3269.090 24.110 3270.270 ;
        RECT 22.930 3267.490 24.110 3268.670 ;
        RECT 22.930 3089.090 24.110 3090.270 ;
        RECT 22.930 3087.490 24.110 3088.670 ;
        RECT 22.930 2909.090 24.110 2910.270 ;
        RECT 22.930 2907.490 24.110 2908.670 ;
        RECT 22.930 2729.090 24.110 2730.270 ;
        RECT 22.930 2727.490 24.110 2728.670 ;
        RECT 22.930 2549.090 24.110 2550.270 ;
        RECT 22.930 2547.490 24.110 2548.670 ;
        RECT 22.930 2369.090 24.110 2370.270 ;
        RECT 22.930 2367.490 24.110 2368.670 ;
        RECT 22.930 2189.090 24.110 2190.270 ;
        RECT 22.930 2187.490 24.110 2188.670 ;
        RECT 22.930 2009.090 24.110 2010.270 ;
        RECT 22.930 2007.490 24.110 2008.670 ;
        RECT 22.930 1829.090 24.110 1830.270 ;
        RECT 22.930 1827.490 24.110 1828.670 ;
        RECT 22.930 1649.090 24.110 1650.270 ;
        RECT 22.930 1647.490 24.110 1648.670 ;
        RECT 22.930 1469.090 24.110 1470.270 ;
        RECT 22.930 1467.490 24.110 1468.670 ;
        RECT 22.930 1289.090 24.110 1290.270 ;
        RECT 22.930 1287.490 24.110 1288.670 ;
        RECT 22.930 1109.090 24.110 1110.270 ;
        RECT 22.930 1107.490 24.110 1108.670 ;
        RECT 22.930 929.090 24.110 930.270 ;
        RECT 22.930 927.490 24.110 928.670 ;
        RECT 22.930 749.090 24.110 750.270 ;
        RECT 22.930 747.490 24.110 748.670 ;
        RECT 22.930 569.090 24.110 570.270 ;
        RECT 22.930 567.490 24.110 568.670 ;
        RECT 22.930 389.090 24.110 390.270 ;
        RECT 22.930 387.490 24.110 388.670 ;
        RECT 22.930 209.090 24.110 210.270 ;
        RECT 22.930 207.490 24.110 208.670 ;
        RECT 22.930 29.090 24.110 30.270 ;
        RECT 22.930 27.490 24.110 28.670 ;
        RECT 22.930 -12.110 24.110 -10.930 ;
        RECT 22.930 -13.710 24.110 -12.530 ;
        RECT 202.930 3532.210 204.110 3533.390 ;
        RECT 202.930 3530.610 204.110 3531.790 ;
        RECT 202.930 3449.090 204.110 3450.270 ;
        RECT 202.930 3447.490 204.110 3448.670 ;
        RECT 202.930 3269.090 204.110 3270.270 ;
        RECT 202.930 3267.490 204.110 3268.670 ;
        RECT 202.930 3089.090 204.110 3090.270 ;
        RECT 202.930 3087.490 204.110 3088.670 ;
        RECT 202.930 2909.090 204.110 2910.270 ;
        RECT 202.930 2907.490 204.110 2908.670 ;
        RECT 202.930 2729.090 204.110 2730.270 ;
        RECT 202.930 2727.490 204.110 2728.670 ;
        RECT 202.930 2549.090 204.110 2550.270 ;
        RECT 202.930 2547.490 204.110 2548.670 ;
        RECT 202.930 2369.090 204.110 2370.270 ;
        RECT 202.930 2367.490 204.110 2368.670 ;
        RECT 202.930 2189.090 204.110 2190.270 ;
        RECT 202.930 2187.490 204.110 2188.670 ;
        RECT 202.930 2009.090 204.110 2010.270 ;
        RECT 202.930 2007.490 204.110 2008.670 ;
        RECT 202.930 1829.090 204.110 1830.270 ;
        RECT 202.930 1827.490 204.110 1828.670 ;
        RECT 202.930 1649.090 204.110 1650.270 ;
        RECT 202.930 1647.490 204.110 1648.670 ;
        RECT 202.930 1469.090 204.110 1470.270 ;
        RECT 202.930 1467.490 204.110 1468.670 ;
        RECT 202.930 1289.090 204.110 1290.270 ;
        RECT 202.930 1287.490 204.110 1288.670 ;
        RECT 202.930 1109.090 204.110 1110.270 ;
        RECT 202.930 1107.490 204.110 1108.670 ;
        RECT 202.930 929.090 204.110 930.270 ;
        RECT 202.930 927.490 204.110 928.670 ;
        RECT 202.930 749.090 204.110 750.270 ;
        RECT 202.930 747.490 204.110 748.670 ;
        RECT 202.930 569.090 204.110 570.270 ;
        RECT 202.930 567.490 204.110 568.670 ;
        RECT 202.930 389.090 204.110 390.270 ;
        RECT 202.930 387.490 204.110 388.670 ;
        RECT 202.930 209.090 204.110 210.270 ;
        RECT 202.930 207.490 204.110 208.670 ;
        RECT 202.930 29.090 204.110 30.270 ;
        RECT 202.930 27.490 204.110 28.670 ;
        RECT 202.930 -12.110 204.110 -10.930 ;
        RECT 202.930 -13.710 204.110 -12.530 ;
        RECT 382.930 3532.210 384.110 3533.390 ;
        RECT 382.930 3530.610 384.110 3531.790 ;
        RECT 382.930 3449.090 384.110 3450.270 ;
        RECT 382.930 3447.490 384.110 3448.670 ;
        RECT 382.930 3269.090 384.110 3270.270 ;
        RECT 382.930 3267.490 384.110 3268.670 ;
        RECT 382.930 3089.090 384.110 3090.270 ;
        RECT 382.930 3087.490 384.110 3088.670 ;
        RECT 382.930 2909.090 384.110 2910.270 ;
        RECT 382.930 2907.490 384.110 2908.670 ;
        RECT 382.930 2729.090 384.110 2730.270 ;
        RECT 382.930 2727.490 384.110 2728.670 ;
        RECT 382.930 2549.090 384.110 2550.270 ;
        RECT 382.930 2547.490 384.110 2548.670 ;
        RECT 382.930 2369.090 384.110 2370.270 ;
        RECT 382.930 2367.490 384.110 2368.670 ;
        RECT 382.930 2189.090 384.110 2190.270 ;
        RECT 382.930 2187.490 384.110 2188.670 ;
        RECT 382.930 2009.090 384.110 2010.270 ;
        RECT 382.930 2007.490 384.110 2008.670 ;
        RECT 382.930 1829.090 384.110 1830.270 ;
        RECT 382.930 1827.490 384.110 1828.670 ;
        RECT 382.930 1649.090 384.110 1650.270 ;
        RECT 382.930 1647.490 384.110 1648.670 ;
        RECT 382.930 1469.090 384.110 1470.270 ;
        RECT 382.930 1467.490 384.110 1468.670 ;
        RECT 382.930 1289.090 384.110 1290.270 ;
        RECT 382.930 1287.490 384.110 1288.670 ;
        RECT 382.930 1109.090 384.110 1110.270 ;
        RECT 382.930 1107.490 384.110 1108.670 ;
        RECT 382.930 929.090 384.110 930.270 ;
        RECT 382.930 927.490 384.110 928.670 ;
        RECT 382.930 749.090 384.110 750.270 ;
        RECT 382.930 747.490 384.110 748.670 ;
        RECT 382.930 569.090 384.110 570.270 ;
        RECT 382.930 567.490 384.110 568.670 ;
        RECT 382.930 389.090 384.110 390.270 ;
        RECT 382.930 387.490 384.110 388.670 ;
        RECT 382.930 209.090 384.110 210.270 ;
        RECT 382.930 207.490 384.110 208.670 ;
        RECT 382.930 29.090 384.110 30.270 ;
        RECT 382.930 27.490 384.110 28.670 ;
        RECT 382.930 -12.110 384.110 -10.930 ;
        RECT 382.930 -13.710 384.110 -12.530 ;
        RECT 562.930 3532.210 564.110 3533.390 ;
        RECT 562.930 3530.610 564.110 3531.790 ;
        RECT 562.930 3449.090 564.110 3450.270 ;
        RECT 562.930 3447.490 564.110 3448.670 ;
        RECT 562.930 3269.090 564.110 3270.270 ;
        RECT 562.930 3267.490 564.110 3268.670 ;
        RECT 562.930 3089.090 564.110 3090.270 ;
        RECT 562.930 3087.490 564.110 3088.670 ;
        RECT 562.930 2909.090 564.110 2910.270 ;
        RECT 562.930 2907.490 564.110 2908.670 ;
        RECT 562.930 2729.090 564.110 2730.270 ;
        RECT 562.930 2727.490 564.110 2728.670 ;
        RECT 562.930 2549.090 564.110 2550.270 ;
        RECT 562.930 2547.490 564.110 2548.670 ;
        RECT 562.930 2369.090 564.110 2370.270 ;
        RECT 562.930 2367.490 564.110 2368.670 ;
        RECT 562.930 2189.090 564.110 2190.270 ;
        RECT 562.930 2187.490 564.110 2188.670 ;
        RECT 562.930 2009.090 564.110 2010.270 ;
        RECT 562.930 2007.490 564.110 2008.670 ;
        RECT 562.930 1829.090 564.110 1830.270 ;
        RECT 562.930 1827.490 564.110 1828.670 ;
        RECT 562.930 1649.090 564.110 1650.270 ;
        RECT 562.930 1647.490 564.110 1648.670 ;
        RECT 562.930 1469.090 564.110 1470.270 ;
        RECT 562.930 1467.490 564.110 1468.670 ;
        RECT 562.930 1289.090 564.110 1290.270 ;
        RECT 562.930 1287.490 564.110 1288.670 ;
        RECT 562.930 1109.090 564.110 1110.270 ;
        RECT 562.930 1107.490 564.110 1108.670 ;
        RECT 562.930 929.090 564.110 930.270 ;
        RECT 562.930 927.490 564.110 928.670 ;
        RECT 562.930 749.090 564.110 750.270 ;
        RECT 562.930 747.490 564.110 748.670 ;
        RECT 562.930 569.090 564.110 570.270 ;
        RECT 562.930 567.490 564.110 568.670 ;
        RECT 562.930 389.090 564.110 390.270 ;
        RECT 562.930 387.490 564.110 388.670 ;
        RECT 562.930 209.090 564.110 210.270 ;
        RECT 562.930 207.490 564.110 208.670 ;
        RECT 562.930 29.090 564.110 30.270 ;
        RECT 562.930 27.490 564.110 28.670 ;
        RECT 562.930 -12.110 564.110 -10.930 ;
        RECT 562.930 -13.710 564.110 -12.530 ;
        RECT 742.930 3532.210 744.110 3533.390 ;
        RECT 742.930 3530.610 744.110 3531.790 ;
        RECT 742.930 3449.090 744.110 3450.270 ;
        RECT 742.930 3447.490 744.110 3448.670 ;
        RECT 742.930 3269.090 744.110 3270.270 ;
        RECT 742.930 3267.490 744.110 3268.670 ;
        RECT 742.930 3089.090 744.110 3090.270 ;
        RECT 742.930 3087.490 744.110 3088.670 ;
        RECT 742.930 2909.090 744.110 2910.270 ;
        RECT 742.930 2907.490 744.110 2908.670 ;
        RECT 742.930 2729.090 744.110 2730.270 ;
        RECT 742.930 2727.490 744.110 2728.670 ;
        RECT 742.930 2549.090 744.110 2550.270 ;
        RECT 742.930 2547.490 744.110 2548.670 ;
        RECT 742.930 2369.090 744.110 2370.270 ;
        RECT 742.930 2367.490 744.110 2368.670 ;
        RECT 742.930 2189.090 744.110 2190.270 ;
        RECT 742.930 2187.490 744.110 2188.670 ;
        RECT 742.930 2009.090 744.110 2010.270 ;
        RECT 742.930 2007.490 744.110 2008.670 ;
        RECT 742.930 1829.090 744.110 1830.270 ;
        RECT 742.930 1827.490 744.110 1828.670 ;
        RECT 742.930 1649.090 744.110 1650.270 ;
        RECT 742.930 1647.490 744.110 1648.670 ;
        RECT 742.930 1469.090 744.110 1470.270 ;
        RECT 742.930 1467.490 744.110 1468.670 ;
        RECT 742.930 1289.090 744.110 1290.270 ;
        RECT 742.930 1287.490 744.110 1288.670 ;
        RECT 742.930 1109.090 744.110 1110.270 ;
        RECT 742.930 1107.490 744.110 1108.670 ;
        RECT 742.930 929.090 744.110 930.270 ;
        RECT 742.930 927.490 744.110 928.670 ;
        RECT 742.930 749.090 744.110 750.270 ;
        RECT 742.930 747.490 744.110 748.670 ;
        RECT 742.930 569.090 744.110 570.270 ;
        RECT 742.930 567.490 744.110 568.670 ;
        RECT 742.930 389.090 744.110 390.270 ;
        RECT 742.930 387.490 744.110 388.670 ;
        RECT 742.930 209.090 744.110 210.270 ;
        RECT 742.930 207.490 744.110 208.670 ;
        RECT 742.930 29.090 744.110 30.270 ;
        RECT 742.930 27.490 744.110 28.670 ;
        RECT 742.930 -12.110 744.110 -10.930 ;
        RECT 742.930 -13.710 744.110 -12.530 ;
        RECT 922.930 3532.210 924.110 3533.390 ;
        RECT 922.930 3530.610 924.110 3531.790 ;
        RECT 922.930 3449.090 924.110 3450.270 ;
        RECT 922.930 3447.490 924.110 3448.670 ;
        RECT 922.930 3269.090 924.110 3270.270 ;
        RECT 922.930 3267.490 924.110 3268.670 ;
        RECT 922.930 3089.090 924.110 3090.270 ;
        RECT 922.930 3087.490 924.110 3088.670 ;
        RECT 922.930 2909.090 924.110 2910.270 ;
        RECT 922.930 2907.490 924.110 2908.670 ;
        RECT 922.930 2729.090 924.110 2730.270 ;
        RECT 922.930 2727.490 924.110 2728.670 ;
        RECT 922.930 2549.090 924.110 2550.270 ;
        RECT 922.930 2547.490 924.110 2548.670 ;
        RECT 922.930 2369.090 924.110 2370.270 ;
        RECT 922.930 2367.490 924.110 2368.670 ;
        RECT 922.930 2189.090 924.110 2190.270 ;
        RECT 922.930 2187.490 924.110 2188.670 ;
        RECT 922.930 2009.090 924.110 2010.270 ;
        RECT 922.930 2007.490 924.110 2008.670 ;
        RECT 922.930 1829.090 924.110 1830.270 ;
        RECT 922.930 1827.490 924.110 1828.670 ;
        RECT 922.930 1649.090 924.110 1650.270 ;
        RECT 922.930 1647.490 924.110 1648.670 ;
        RECT 922.930 1469.090 924.110 1470.270 ;
        RECT 922.930 1467.490 924.110 1468.670 ;
        RECT 922.930 1289.090 924.110 1290.270 ;
        RECT 922.930 1287.490 924.110 1288.670 ;
        RECT 922.930 1109.090 924.110 1110.270 ;
        RECT 922.930 1107.490 924.110 1108.670 ;
        RECT 922.930 929.090 924.110 930.270 ;
        RECT 922.930 927.490 924.110 928.670 ;
        RECT 922.930 749.090 924.110 750.270 ;
        RECT 922.930 747.490 924.110 748.670 ;
        RECT 922.930 569.090 924.110 570.270 ;
        RECT 922.930 567.490 924.110 568.670 ;
        RECT 922.930 389.090 924.110 390.270 ;
        RECT 922.930 387.490 924.110 388.670 ;
        RECT 922.930 209.090 924.110 210.270 ;
        RECT 922.930 207.490 924.110 208.670 ;
        RECT 922.930 29.090 924.110 30.270 ;
        RECT 922.930 27.490 924.110 28.670 ;
        RECT 922.930 -12.110 924.110 -10.930 ;
        RECT 922.930 -13.710 924.110 -12.530 ;
        RECT 1102.930 3532.210 1104.110 3533.390 ;
        RECT 1102.930 3530.610 1104.110 3531.790 ;
        RECT 1102.930 3449.090 1104.110 3450.270 ;
        RECT 1102.930 3447.490 1104.110 3448.670 ;
        RECT 1102.930 3269.090 1104.110 3270.270 ;
        RECT 1102.930 3267.490 1104.110 3268.670 ;
        RECT 1102.930 3089.090 1104.110 3090.270 ;
        RECT 1102.930 3087.490 1104.110 3088.670 ;
        RECT 1102.930 2909.090 1104.110 2910.270 ;
        RECT 1102.930 2907.490 1104.110 2908.670 ;
        RECT 1102.930 2729.090 1104.110 2730.270 ;
        RECT 1102.930 2727.490 1104.110 2728.670 ;
        RECT 1102.930 2549.090 1104.110 2550.270 ;
        RECT 1102.930 2547.490 1104.110 2548.670 ;
        RECT 1102.930 2369.090 1104.110 2370.270 ;
        RECT 1102.930 2367.490 1104.110 2368.670 ;
        RECT 1102.930 2189.090 1104.110 2190.270 ;
        RECT 1102.930 2187.490 1104.110 2188.670 ;
        RECT 1102.930 2009.090 1104.110 2010.270 ;
        RECT 1102.930 2007.490 1104.110 2008.670 ;
        RECT 1102.930 1829.090 1104.110 1830.270 ;
        RECT 1102.930 1827.490 1104.110 1828.670 ;
        RECT 1102.930 1649.090 1104.110 1650.270 ;
        RECT 1102.930 1647.490 1104.110 1648.670 ;
        RECT 1102.930 1469.090 1104.110 1470.270 ;
        RECT 1102.930 1467.490 1104.110 1468.670 ;
        RECT 1102.930 1289.090 1104.110 1290.270 ;
        RECT 1102.930 1287.490 1104.110 1288.670 ;
        RECT 1102.930 1109.090 1104.110 1110.270 ;
        RECT 1102.930 1107.490 1104.110 1108.670 ;
        RECT 1102.930 929.090 1104.110 930.270 ;
        RECT 1102.930 927.490 1104.110 928.670 ;
        RECT 1102.930 749.090 1104.110 750.270 ;
        RECT 1102.930 747.490 1104.110 748.670 ;
        RECT 1102.930 569.090 1104.110 570.270 ;
        RECT 1102.930 567.490 1104.110 568.670 ;
        RECT 1102.930 389.090 1104.110 390.270 ;
        RECT 1102.930 387.490 1104.110 388.670 ;
        RECT 1102.930 209.090 1104.110 210.270 ;
        RECT 1102.930 207.490 1104.110 208.670 ;
        RECT 1102.930 29.090 1104.110 30.270 ;
        RECT 1102.930 27.490 1104.110 28.670 ;
        RECT 1102.930 -12.110 1104.110 -10.930 ;
        RECT 1102.930 -13.710 1104.110 -12.530 ;
        RECT 1282.930 3532.210 1284.110 3533.390 ;
        RECT 1282.930 3530.610 1284.110 3531.790 ;
        RECT 1282.930 3449.090 1284.110 3450.270 ;
        RECT 1282.930 3447.490 1284.110 3448.670 ;
        RECT 1282.930 3269.090 1284.110 3270.270 ;
        RECT 1282.930 3267.490 1284.110 3268.670 ;
        RECT 1282.930 3089.090 1284.110 3090.270 ;
        RECT 1282.930 3087.490 1284.110 3088.670 ;
        RECT 1282.930 2909.090 1284.110 2910.270 ;
        RECT 1282.930 2907.490 1284.110 2908.670 ;
        RECT 1282.930 2729.090 1284.110 2730.270 ;
        RECT 1282.930 2727.490 1284.110 2728.670 ;
        RECT 1282.930 2549.090 1284.110 2550.270 ;
        RECT 1282.930 2547.490 1284.110 2548.670 ;
        RECT 1282.930 2369.090 1284.110 2370.270 ;
        RECT 1282.930 2367.490 1284.110 2368.670 ;
        RECT 1282.930 2189.090 1284.110 2190.270 ;
        RECT 1282.930 2187.490 1284.110 2188.670 ;
        RECT 1282.930 2009.090 1284.110 2010.270 ;
        RECT 1282.930 2007.490 1284.110 2008.670 ;
        RECT 1282.930 1829.090 1284.110 1830.270 ;
        RECT 1282.930 1827.490 1284.110 1828.670 ;
        RECT 1282.930 1649.090 1284.110 1650.270 ;
        RECT 1282.930 1647.490 1284.110 1648.670 ;
        RECT 1282.930 1469.090 1284.110 1470.270 ;
        RECT 1282.930 1467.490 1284.110 1468.670 ;
        RECT 1282.930 1289.090 1284.110 1290.270 ;
        RECT 1282.930 1287.490 1284.110 1288.670 ;
        RECT 1282.930 1109.090 1284.110 1110.270 ;
        RECT 1282.930 1107.490 1284.110 1108.670 ;
        RECT 1282.930 929.090 1284.110 930.270 ;
        RECT 1282.930 927.490 1284.110 928.670 ;
        RECT 1282.930 749.090 1284.110 750.270 ;
        RECT 1282.930 747.490 1284.110 748.670 ;
        RECT 1282.930 569.090 1284.110 570.270 ;
        RECT 1282.930 567.490 1284.110 568.670 ;
        RECT 1282.930 389.090 1284.110 390.270 ;
        RECT 1282.930 387.490 1284.110 388.670 ;
        RECT 1282.930 209.090 1284.110 210.270 ;
        RECT 1282.930 207.490 1284.110 208.670 ;
        RECT 1282.930 29.090 1284.110 30.270 ;
        RECT 1282.930 27.490 1284.110 28.670 ;
        RECT 1282.930 -12.110 1284.110 -10.930 ;
        RECT 1282.930 -13.710 1284.110 -12.530 ;
        RECT 1462.930 3532.210 1464.110 3533.390 ;
        RECT 1462.930 3530.610 1464.110 3531.790 ;
        RECT 1462.930 3449.090 1464.110 3450.270 ;
        RECT 1462.930 3447.490 1464.110 3448.670 ;
        RECT 1462.930 3269.090 1464.110 3270.270 ;
        RECT 1462.930 3267.490 1464.110 3268.670 ;
        RECT 1462.930 3089.090 1464.110 3090.270 ;
        RECT 1462.930 3087.490 1464.110 3088.670 ;
        RECT 1462.930 2909.090 1464.110 2910.270 ;
        RECT 1462.930 2907.490 1464.110 2908.670 ;
        RECT 1462.930 2729.090 1464.110 2730.270 ;
        RECT 1462.930 2727.490 1464.110 2728.670 ;
        RECT 1462.930 2549.090 1464.110 2550.270 ;
        RECT 1462.930 2547.490 1464.110 2548.670 ;
        RECT 1462.930 2369.090 1464.110 2370.270 ;
        RECT 1462.930 2367.490 1464.110 2368.670 ;
        RECT 1462.930 2189.090 1464.110 2190.270 ;
        RECT 1462.930 2187.490 1464.110 2188.670 ;
        RECT 1462.930 2009.090 1464.110 2010.270 ;
        RECT 1462.930 2007.490 1464.110 2008.670 ;
        RECT 1462.930 1829.090 1464.110 1830.270 ;
        RECT 1462.930 1827.490 1464.110 1828.670 ;
        RECT 1462.930 1649.090 1464.110 1650.270 ;
        RECT 1462.930 1647.490 1464.110 1648.670 ;
        RECT 1462.930 1469.090 1464.110 1470.270 ;
        RECT 1462.930 1467.490 1464.110 1468.670 ;
        RECT 1462.930 1289.090 1464.110 1290.270 ;
        RECT 1462.930 1287.490 1464.110 1288.670 ;
        RECT 1462.930 1109.090 1464.110 1110.270 ;
        RECT 1462.930 1107.490 1464.110 1108.670 ;
        RECT 1462.930 929.090 1464.110 930.270 ;
        RECT 1462.930 927.490 1464.110 928.670 ;
        RECT 1462.930 749.090 1464.110 750.270 ;
        RECT 1462.930 747.490 1464.110 748.670 ;
        RECT 1462.930 569.090 1464.110 570.270 ;
        RECT 1462.930 567.490 1464.110 568.670 ;
        RECT 1462.930 389.090 1464.110 390.270 ;
        RECT 1462.930 387.490 1464.110 388.670 ;
        RECT 1462.930 209.090 1464.110 210.270 ;
        RECT 1462.930 207.490 1464.110 208.670 ;
        RECT 1462.930 29.090 1464.110 30.270 ;
        RECT 1462.930 27.490 1464.110 28.670 ;
        RECT 1462.930 -12.110 1464.110 -10.930 ;
        RECT 1462.930 -13.710 1464.110 -12.530 ;
        RECT 1642.930 3532.210 1644.110 3533.390 ;
        RECT 1642.930 3530.610 1644.110 3531.790 ;
        RECT 1642.930 3449.090 1644.110 3450.270 ;
        RECT 1642.930 3447.490 1644.110 3448.670 ;
        RECT 1642.930 3269.090 1644.110 3270.270 ;
        RECT 1642.930 3267.490 1644.110 3268.670 ;
        RECT 1642.930 3089.090 1644.110 3090.270 ;
        RECT 1642.930 3087.490 1644.110 3088.670 ;
        RECT 1642.930 2909.090 1644.110 2910.270 ;
        RECT 1642.930 2907.490 1644.110 2908.670 ;
        RECT 1642.930 2729.090 1644.110 2730.270 ;
        RECT 1642.930 2727.490 1644.110 2728.670 ;
        RECT 1642.930 2549.090 1644.110 2550.270 ;
        RECT 1642.930 2547.490 1644.110 2548.670 ;
        RECT 1642.930 2369.090 1644.110 2370.270 ;
        RECT 1642.930 2367.490 1644.110 2368.670 ;
        RECT 1642.930 2189.090 1644.110 2190.270 ;
        RECT 1642.930 2187.490 1644.110 2188.670 ;
        RECT 1642.930 2009.090 1644.110 2010.270 ;
        RECT 1642.930 2007.490 1644.110 2008.670 ;
        RECT 1642.930 1829.090 1644.110 1830.270 ;
        RECT 1642.930 1827.490 1644.110 1828.670 ;
        RECT 1642.930 1649.090 1644.110 1650.270 ;
        RECT 1642.930 1647.490 1644.110 1648.670 ;
        RECT 1642.930 1469.090 1644.110 1470.270 ;
        RECT 1642.930 1467.490 1644.110 1468.670 ;
        RECT 1642.930 1289.090 1644.110 1290.270 ;
        RECT 1642.930 1287.490 1644.110 1288.670 ;
        RECT 1642.930 1109.090 1644.110 1110.270 ;
        RECT 1642.930 1107.490 1644.110 1108.670 ;
        RECT 1642.930 929.090 1644.110 930.270 ;
        RECT 1642.930 927.490 1644.110 928.670 ;
        RECT 1642.930 749.090 1644.110 750.270 ;
        RECT 1642.930 747.490 1644.110 748.670 ;
        RECT 1642.930 569.090 1644.110 570.270 ;
        RECT 1642.930 567.490 1644.110 568.670 ;
        RECT 1642.930 389.090 1644.110 390.270 ;
        RECT 1642.930 387.490 1644.110 388.670 ;
        RECT 1642.930 209.090 1644.110 210.270 ;
        RECT 1642.930 207.490 1644.110 208.670 ;
        RECT 1642.930 29.090 1644.110 30.270 ;
        RECT 1642.930 27.490 1644.110 28.670 ;
        RECT 1642.930 -12.110 1644.110 -10.930 ;
        RECT 1642.930 -13.710 1644.110 -12.530 ;
        RECT 1822.930 3532.210 1824.110 3533.390 ;
        RECT 1822.930 3530.610 1824.110 3531.790 ;
        RECT 1822.930 3449.090 1824.110 3450.270 ;
        RECT 1822.930 3447.490 1824.110 3448.670 ;
        RECT 1822.930 3269.090 1824.110 3270.270 ;
        RECT 1822.930 3267.490 1824.110 3268.670 ;
        RECT 1822.930 3089.090 1824.110 3090.270 ;
        RECT 1822.930 3087.490 1824.110 3088.670 ;
        RECT 1822.930 2909.090 1824.110 2910.270 ;
        RECT 1822.930 2907.490 1824.110 2908.670 ;
        RECT 1822.930 2729.090 1824.110 2730.270 ;
        RECT 1822.930 2727.490 1824.110 2728.670 ;
        RECT 1822.930 2549.090 1824.110 2550.270 ;
        RECT 1822.930 2547.490 1824.110 2548.670 ;
        RECT 1822.930 2369.090 1824.110 2370.270 ;
        RECT 1822.930 2367.490 1824.110 2368.670 ;
        RECT 1822.930 2189.090 1824.110 2190.270 ;
        RECT 1822.930 2187.490 1824.110 2188.670 ;
        RECT 1822.930 2009.090 1824.110 2010.270 ;
        RECT 1822.930 2007.490 1824.110 2008.670 ;
        RECT 1822.930 1829.090 1824.110 1830.270 ;
        RECT 1822.930 1827.490 1824.110 1828.670 ;
        RECT 1822.930 1649.090 1824.110 1650.270 ;
        RECT 1822.930 1647.490 1824.110 1648.670 ;
        RECT 1822.930 1469.090 1824.110 1470.270 ;
        RECT 1822.930 1467.490 1824.110 1468.670 ;
        RECT 1822.930 1289.090 1824.110 1290.270 ;
        RECT 1822.930 1287.490 1824.110 1288.670 ;
        RECT 1822.930 1109.090 1824.110 1110.270 ;
        RECT 1822.930 1107.490 1824.110 1108.670 ;
        RECT 1822.930 929.090 1824.110 930.270 ;
        RECT 1822.930 927.490 1824.110 928.670 ;
        RECT 1822.930 749.090 1824.110 750.270 ;
        RECT 1822.930 747.490 1824.110 748.670 ;
        RECT 1822.930 569.090 1824.110 570.270 ;
        RECT 1822.930 567.490 1824.110 568.670 ;
        RECT 1822.930 389.090 1824.110 390.270 ;
        RECT 1822.930 387.490 1824.110 388.670 ;
        RECT 1822.930 209.090 1824.110 210.270 ;
        RECT 1822.930 207.490 1824.110 208.670 ;
        RECT 1822.930 29.090 1824.110 30.270 ;
        RECT 1822.930 27.490 1824.110 28.670 ;
        RECT 1822.930 -12.110 1824.110 -10.930 ;
        RECT 1822.930 -13.710 1824.110 -12.530 ;
        RECT 2002.930 3532.210 2004.110 3533.390 ;
        RECT 2002.930 3530.610 2004.110 3531.790 ;
        RECT 2002.930 3449.090 2004.110 3450.270 ;
        RECT 2002.930 3447.490 2004.110 3448.670 ;
        RECT 2002.930 3269.090 2004.110 3270.270 ;
        RECT 2002.930 3267.490 2004.110 3268.670 ;
        RECT 2002.930 3089.090 2004.110 3090.270 ;
        RECT 2002.930 3087.490 2004.110 3088.670 ;
        RECT 2002.930 2909.090 2004.110 2910.270 ;
        RECT 2002.930 2907.490 2004.110 2908.670 ;
        RECT 2002.930 2729.090 2004.110 2730.270 ;
        RECT 2002.930 2727.490 2004.110 2728.670 ;
        RECT 2002.930 2549.090 2004.110 2550.270 ;
        RECT 2002.930 2547.490 2004.110 2548.670 ;
        RECT 2002.930 2369.090 2004.110 2370.270 ;
        RECT 2002.930 2367.490 2004.110 2368.670 ;
        RECT 2002.930 2189.090 2004.110 2190.270 ;
        RECT 2002.930 2187.490 2004.110 2188.670 ;
        RECT 2002.930 2009.090 2004.110 2010.270 ;
        RECT 2002.930 2007.490 2004.110 2008.670 ;
        RECT 2002.930 1829.090 2004.110 1830.270 ;
        RECT 2002.930 1827.490 2004.110 1828.670 ;
        RECT 2002.930 1649.090 2004.110 1650.270 ;
        RECT 2002.930 1647.490 2004.110 1648.670 ;
        RECT 2002.930 1469.090 2004.110 1470.270 ;
        RECT 2002.930 1467.490 2004.110 1468.670 ;
        RECT 2002.930 1289.090 2004.110 1290.270 ;
        RECT 2002.930 1287.490 2004.110 1288.670 ;
        RECT 2002.930 1109.090 2004.110 1110.270 ;
        RECT 2002.930 1107.490 2004.110 1108.670 ;
        RECT 2002.930 929.090 2004.110 930.270 ;
        RECT 2002.930 927.490 2004.110 928.670 ;
        RECT 2002.930 749.090 2004.110 750.270 ;
        RECT 2002.930 747.490 2004.110 748.670 ;
        RECT 2002.930 569.090 2004.110 570.270 ;
        RECT 2002.930 567.490 2004.110 568.670 ;
        RECT 2002.930 389.090 2004.110 390.270 ;
        RECT 2002.930 387.490 2004.110 388.670 ;
        RECT 2002.930 209.090 2004.110 210.270 ;
        RECT 2002.930 207.490 2004.110 208.670 ;
        RECT 2002.930 29.090 2004.110 30.270 ;
        RECT 2002.930 27.490 2004.110 28.670 ;
        RECT 2002.930 -12.110 2004.110 -10.930 ;
        RECT 2002.930 -13.710 2004.110 -12.530 ;
        RECT 2182.930 3532.210 2184.110 3533.390 ;
        RECT 2182.930 3530.610 2184.110 3531.790 ;
        RECT 2182.930 3449.090 2184.110 3450.270 ;
        RECT 2182.930 3447.490 2184.110 3448.670 ;
        RECT 2182.930 3269.090 2184.110 3270.270 ;
        RECT 2182.930 3267.490 2184.110 3268.670 ;
        RECT 2182.930 3089.090 2184.110 3090.270 ;
        RECT 2182.930 3087.490 2184.110 3088.670 ;
        RECT 2182.930 2909.090 2184.110 2910.270 ;
        RECT 2182.930 2907.490 2184.110 2908.670 ;
        RECT 2182.930 2729.090 2184.110 2730.270 ;
        RECT 2182.930 2727.490 2184.110 2728.670 ;
        RECT 2182.930 2549.090 2184.110 2550.270 ;
        RECT 2182.930 2547.490 2184.110 2548.670 ;
        RECT 2182.930 2369.090 2184.110 2370.270 ;
        RECT 2182.930 2367.490 2184.110 2368.670 ;
        RECT 2182.930 2189.090 2184.110 2190.270 ;
        RECT 2182.930 2187.490 2184.110 2188.670 ;
        RECT 2182.930 2009.090 2184.110 2010.270 ;
        RECT 2182.930 2007.490 2184.110 2008.670 ;
        RECT 2182.930 1829.090 2184.110 1830.270 ;
        RECT 2182.930 1827.490 2184.110 1828.670 ;
        RECT 2182.930 1649.090 2184.110 1650.270 ;
        RECT 2182.930 1647.490 2184.110 1648.670 ;
        RECT 2182.930 1469.090 2184.110 1470.270 ;
        RECT 2182.930 1467.490 2184.110 1468.670 ;
        RECT 2182.930 1289.090 2184.110 1290.270 ;
        RECT 2182.930 1287.490 2184.110 1288.670 ;
        RECT 2182.930 1109.090 2184.110 1110.270 ;
        RECT 2182.930 1107.490 2184.110 1108.670 ;
        RECT 2182.930 929.090 2184.110 930.270 ;
        RECT 2182.930 927.490 2184.110 928.670 ;
        RECT 2182.930 749.090 2184.110 750.270 ;
        RECT 2182.930 747.490 2184.110 748.670 ;
        RECT 2182.930 569.090 2184.110 570.270 ;
        RECT 2182.930 567.490 2184.110 568.670 ;
        RECT 2182.930 389.090 2184.110 390.270 ;
        RECT 2182.930 387.490 2184.110 388.670 ;
        RECT 2182.930 209.090 2184.110 210.270 ;
        RECT 2182.930 207.490 2184.110 208.670 ;
        RECT 2182.930 29.090 2184.110 30.270 ;
        RECT 2182.930 27.490 2184.110 28.670 ;
        RECT 2182.930 -12.110 2184.110 -10.930 ;
        RECT 2182.930 -13.710 2184.110 -12.530 ;
        RECT 2362.930 3532.210 2364.110 3533.390 ;
        RECT 2362.930 3530.610 2364.110 3531.790 ;
        RECT 2362.930 3449.090 2364.110 3450.270 ;
        RECT 2362.930 3447.490 2364.110 3448.670 ;
        RECT 2362.930 3269.090 2364.110 3270.270 ;
        RECT 2362.930 3267.490 2364.110 3268.670 ;
        RECT 2362.930 3089.090 2364.110 3090.270 ;
        RECT 2362.930 3087.490 2364.110 3088.670 ;
        RECT 2362.930 2909.090 2364.110 2910.270 ;
        RECT 2362.930 2907.490 2364.110 2908.670 ;
        RECT 2362.930 2729.090 2364.110 2730.270 ;
        RECT 2362.930 2727.490 2364.110 2728.670 ;
        RECT 2362.930 2549.090 2364.110 2550.270 ;
        RECT 2362.930 2547.490 2364.110 2548.670 ;
        RECT 2362.930 2369.090 2364.110 2370.270 ;
        RECT 2362.930 2367.490 2364.110 2368.670 ;
        RECT 2362.930 2189.090 2364.110 2190.270 ;
        RECT 2362.930 2187.490 2364.110 2188.670 ;
        RECT 2362.930 2009.090 2364.110 2010.270 ;
        RECT 2362.930 2007.490 2364.110 2008.670 ;
        RECT 2362.930 1829.090 2364.110 1830.270 ;
        RECT 2362.930 1827.490 2364.110 1828.670 ;
        RECT 2362.930 1649.090 2364.110 1650.270 ;
        RECT 2362.930 1647.490 2364.110 1648.670 ;
        RECT 2362.930 1469.090 2364.110 1470.270 ;
        RECT 2362.930 1467.490 2364.110 1468.670 ;
        RECT 2362.930 1289.090 2364.110 1290.270 ;
        RECT 2362.930 1287.490 2364.110 1288.670 ;
        RECT 2362.930 1109.090 2364.110 1110.270 ;
        RECT 2362.930 1107.490 2364.110 1108.670 ;
        RECT 2362.930 929.090 2364.110 930.270 ;
        RECT 2362.930 927.490 2364.110 928.670 ;
        RECT 2362.930 749.090 2364.110 750.270 ;
        RECT 2362.930 747.490 2364.110 748.670 ;
        RECT 2362.930 569.090 2364.110 570.270 ;
        RECT 2362.930 567.490 2364.110 568.670 ;
        RECT 2362.930 389.090 2364.110 390.270 ;
        RECT 2362.930 387.490 2364.110 388.670 ;
        RECT 2362.930 209.090 2364.110 210.270 ;
        RECT 2362.930 207.490 2364.110 208.670 ;
        RECT 2362.930 29.090 2364.110 30.270 ;
        RECT 2362.930 27.490 2364.110 28.670 ;
        RECT 2362.930 -12.110 2364.110 -10.930 ;
        RECT 2362.930 -13.710 2364.110 -12.530 ;
        RECT 2542.930 3532.210 2544.110 3533.390 ;
        RECT 2542.930 3530.610 2544.110 3531.790 ;
        RECT 2542.930 3449.090 2544.110 3450.270 ;
        RECT 2542.930 3447.490 2544.110 3448.670 ;
        RECT 2542.930 3269.090 2544.110 3270.270 ;
        RECT 2542.930 3267.490 2544.110 3268.670 ;
        RECT 2542.930 3089.090 2544.110 3090.270 ;
        RECT 2542.930 3087.490 2544.110 3088.670 ;
        RECT 2542.930 2909.090 2544.110 2910.270 ;
        RECT 2542.930 2907.490 2544.110 2908.670 ;
        RECT 2542.930 2729.090 2544.110 2730.270 ;
        RECT 2542.930 2727.490 2544.110 2728.670 ;
        RECT 2542.930 2549.090 2544.110 2550.270 ;
        RECT 2542.930 2547.490 2544.110 2548.670 ;
        RECT 2542.930 2369.090 2544.110 2370.270 ;
        RECT 2542.930 2367.490 2544.110 2368.670 ;
        RECT 2542.930 2189.090 2544.110 2190.270 ;
        RECT 2542.930 2187.490 2544.110 2188.670 ;
        RECT 2542.930 2009.090 2544.110 2010.270 ;
        RECT 2542.930 2007.490 2544.110 2008.670 ;
        RECT 2542.930 1829.090 2544.110 1830.270 ;
        RECT 2542.930 1827.490 2544.110 1828.670 ;
        RECT 2542.930 1649.090 2544.110 1650.270 ;
        RECT 2542.930 1647.490 2544.110 1648.670 ;
        RECT 2542.930 1469.090 2544.110 1470.270 ;
        RECT 2542.930 1467.490 2544.110 1468.670 ;
        RECT 2542.930 1289.090 2544.110 1290.270 ;
        RECT 2542.930 1287.490 2544.110 1288.670 ;
        RECT 2542.930 1109.090 2544.110 1110.270 ;
        RECT 2542.930 1107.490 2544.110 1108.670 ;
        RECT 2542.930 929.090 2544.110 930.270 ;
        RECT 2542.930 927.490 2544.110 928.670 ;
        RECT 2542.930 749.090 2544.110 750.270 ;
        RECT 2542.930 747.490 2544.110 748.670 ;
        RECT 2542.930 569.090 2544.110 570.270 ;
        RECT 2542.930 567.490 2544.110 568.670 ;
        RECT 2542.930 389.090 2544.110 390.270 ;
        RECT 2542.930 387.490 2544.110 388.670 ;
        RECT 2542.930 209.090 2544.110 210.270 ;
        RECT 2542.930 207.490 2544.110 208.670 ;
        RECT 2542.930 29.090 2544.110 30.270 ;
        RECT 2542.930 27.490 2544.110 28.670 ;
        RECT 2542.930 -12.110 2544.110 -10.930 ;
        RECT 2542.930 -13.710 2544.110 -12.530 ;
        RECT 2722.930 3532.210 2724.110 3533.390 ;
        RECT 2722.930 3530.610 2724.110 3531.790 ;
        RECT 2722.930 3449.090 2724.110 3450.270 ;
        RECT 2722.930 3447.490 2724.110 3448.670 ;
        RECT 2722.930 3269.090 2724.110 3270.270 ;
        RECT 2722.930 3267.490 2724.110 3268.670 ;
        RECT 2722.930 3089.090 2724.110 3090.270 ;
        RECT 2722.930 3087.490 2724.110 3088.670 ;
        RECT 2722.930 2909.090 2724.110 2910.270 ;
        RECT 2722.930 2907.490 2724.110 2908.670 ;
        RECT 2722.930 2729.090 2724.110 2730.270 ;
        RECT 2722.930 2727.490 2724.110 2728.670 ;
        RECT 2722.930 2549.090 2724.110 2550.270 ;
        RECT 2722.930 2547.490 2724.110 2548.670 ;
        RECT 2722.930 2369.090 2724.110 2370.270 ;
        RECT 2722.930 2367.490 2724.110 2368.670 ;
        RECT 2722.930 2189.090 2724.110 2190.270 ;
        RECT 2722.930 2187.490 2724.110 2188.670 ;
        RECT 2722.930 2009.090 2724.110 2010.270 ;
        RECT 2722.930 2007.490 2724.110 2008.670 ;
        RECT 2722.930 1829.090 2724.110 1830.270 ;
        RECT 2722.930 1827.490 2724.110 1828.670 ;
        RECT 2722.930 1649.090 2724.110 1650.270 ;
        RECT 2722.930 1647.490 2724.110 1648.670 ;
        RECT 2722.930 1469.090 2724.110 1470.270 ;
        RECT 2722.930 1467.490 2724.110 1468.670 ;
        RECT 2722.930 1289.090 2724.110 1290.270 ;
        RECT 2722.930 1287.490 2724.110 1288.670 ;
        RECT 2722.930 1109.090 2724.110 1110.270 ;
        RECT 2722.930 1107.490 2724.110 1108.670 ;
        RECT 2722.930 929.090 2724.110 930.270 ;
        RECT 2722.930 927.490 2724.110 928.670 ;
        RECT 2722.930 749.090 2724.110 750.270 ;
        RECT 2722.930 747.490 2724.110 748.670 ;
        RECT 2722.930 569.090 2724.110 570.270 ;
        RECT 2722.930 567.490 2724.110 568.670 ;
        RECT 2722.930 389.090 2724.110 390.270 ;
        RECT 2722.930 387.490 2724.110 388.670 ;
        RECT 2722.930 209.090 2724.110 210.270 ;
        RECT 2722.930 207.490 2724.110 208.670 ;
        RECT 2722.930 29.090 2724.110 30.270 ;
        RECT 2722.930 27.490 2724.110 28.670 ;
        RECT 2722.930 -12.110 2724.110 -10.930 ;
        RECT 2722.930 -13.710 2724.110 -12.530 ;
        RECT 2902.930 3532.210 2904.110 3533.390 ;
        RECT 2902.930 3530.610 2904.110 3531.790 ;
        RECT 2902.930 3449.090 2904.110 3450.270 ;
        RECT 2902.930 3447.490 2904.110 3448.670 ;
        RECT 2902.930 3269.090 2904.110 3270.270 ;
        RECT 2902.930 3267.490 2904.110 3268.670 ;
        RECT 2902.930 3089.090 2904.110 3090.270 ;
        RECT 2902.930 3087.490 2904.110 3088.670 ;
        RECT 2902.930 2909.090 2904.110 2910.270 ;
        RECT 2902.930 2907.490 2904.110 2908.670 ;
        RECT 2902.930 2729.090 2904.110 2730.270 ;
        RECT 2902.930 2727.490 2904.110 2728.670 ;
        RECT 2902.930 2549.090 2904.110 2550.270 ;
        RECT 2902.930 2547.490 2904.110 2548.670 ;
        RECT 2902.930 2369.090 2904.110 2370.270 ;
        RECT 2902.930 2367.490 2904.110 2368.670 ;
        RECT 2902.930 2189.090 2904.110 2190.270 ;
        RECT 2902.930 2187.490 2904.110 2188.670 ;
        RECT 2902.930 2009.090 2904.110 2010.270 ;
        RECT 2902.930 2007.490 2904.110 2008.670 ;
        RECT 2902.930 1829.090 2904.110 1830.270 ;
        RECT 2902.930 1827.490 2904.110 1828.670 ;
        RECT 2902.930 1649.090 2904.110 1650.270 ;
        RECT 2902.930 1647.490 2904.110 1648.670 ;
        RECT 2902.930 1469.090 2904.110 1470.270 ;
        RECT 2902.930 1467.490 2904.110 1468.670 ;
        RECT 2902.930 1289.090 2904.110 1290.270 ;
        RECT 2902.930 1287.490 2904.110 1288.670 ;
        RECT 2902.930 1109.090 2904.110 1110.270 ;
        RECT 2902.930 1107.490 2904.110 1108.670 ;
        RECT 2902.930 929.090 2904.110 930.270 ;
        RECT 2902.930 927.490 2904.110 928.670 ;
        RECT 2902.930 749.090 2904.110 750.270 ;
        RECT 2902.930 747.490 2904.110 748.670 ;
        RECT 2902.930 569.090 2904.110 570.270 ;
        RECT 2902.930 567.490 2904.110 568.670 ;
        RECT 2902.930 389.090 2904.110 390.270 ;
        RECT 2902.930 387.490 2904.110 388.670 ;
        RECT 2902.930 209.090 2904.110 210.270 ;
        RECT 2902.930 207.490 2904.110 208.670 ;
        RECT 2902.930 29.090 2904.110 30.270 ;
        RECT 2902.930 27.490 2904.110 28.670 ;
        RECT 2902.930 -12.110 2904.110 -10.930 ;
        RECT 2902.930 -13.710 2904.110 -12.530 ;
        RECT 2936.710 3532.210 2937.890 3533.390 ;
        RECT 2936.710 3530.610 2937.890 3531.790 ;
        RECT 2936.710 3449.090 2937.890 3450.270 ;
        RECT 2936.710 3447.490 2937.890 3448.670 ;
        RECT 2936.710 3269.090 2937.890 3270.270 ;
        RECT 2936.710 3267.490 2937.890 3268.670 ;
        RECT 2936.710 3089.090 2937.890 3090.270 ;
        RECT 2936.710 3087.490 2937.890 3088.670 ;
        RECT 2936.710 2909.090 2937.890 2910.270 ;
        RECT 2936.710 2907.490 2937.890 2908.670 ;
        RECT 2936.710 2729.090 2937.890 2730.270 ;
        RECT 2936.710 2727.490 2937.890 2728.670 ;
        RECT 2936.710 2549.090 2937.890 2550.270 ;
        RECT 2936.710 2547.490 2937.890 2548.670 ;
        RECT 2936.710 2369.090 2937.890 2370.270 ;
        RECT 2936.710 2367.490 2937.890 2368.670 ;
        RECT 2936.710 2189.090 2937.890 2190.270 ;
        RECT 2936.710 2187.490 2937.890 2188.670 ;
        RECT 2936.710 2009.090 2937.890 2010.270 ;
        RECT 2936.710 2007.490 2937.890 2008.670 ;
        RECT 2936.710 1829.090 2937.890 1830.270 ;
        RECT 2936.710 1827.490 2937.890 1828.670 ;
        RECT 2936.710 1649.090 2937.890 1650.270 ;
        RECT 2936.710 1647.490 2937.890 1648.670 ;
        RECT 2936.710 1469.090 2937.890 1470.270 ;
        RECT 2936.710 1467.490 2937.890 1468.670 ;
        RECT 2936.710 1289.090 2937.890 1290.270 ;
        RECT 2936.710 1287.490 2937.890 1288.670 ;
        RECT 2936.710 1109.090 2937.890 1110.270 ;
        RECT 2936.710 1107.490 2937.890 1108.670 ;
        RECT 2936.710 929.090 2937.890 930.270 ;
        RECT 2936.710 927.490 2937.890 928.670 ;
        RECT 2936.710 749.090 2937.890 750.270 ;
        RECT 2936.710 747.490 2937.890 748.670 ;
        RECT 2936.710 569.090 2937.890 570.270 ;
        RECT 2936.710 567.490 2937.890 568.670 ;
        RECT 2936.710 389.090 2937.890 390.270 ;
        RECT 2936.710 387.490 2937.890 388.670 ;
        RECT 2936.710 209.090 2937.890 210.270 ;
        RECT 2936.710 207.490 2937.890 208.670 ;
        RECT 2936.710 29.090 2937.890 30.270 ;
        RECT 2936.710 27.490 2937.890 28.670 ;
        RECT 2936.710 -12.110 2937.890 -10.930 ;
        RECT 2936.710 -13.710 2937.890 -12.530 ;
      LAYER met5 ;
        RECT -19.180 3533.500 -16.180 3533.510 ;
        RECT 22.020 3533.500 25.020 3533.510 ;
        RECT 202.020 3533.500 205.020 3533.510 ;
        RECT 382.020 3533.500 385.020 3533.510 ;
        RECT 562.020 3533.500 565.020 3533.510 ;
        RECT 742.020 3533.500 745.020 3533.510 ;
        RECT 922.020 3533.500 925.020 3533.510 ;
        RECT 1102.020 3533.500 1105.020 3533.510 ;
        RECT 1282.020 3533.500 1285.020 3533.510 ;
        RECT 1462.020 3533.500 1465.020 3533.510 ;
        RECT 1642.020 3533.500 1645.020 3533.510 ;
        RECT 1822.020 3533.500 1825.020 3533.510 ;
        RECT 2002.020 3533.500 2005.020 3533.510 ;
        RECT 2182.020 3533.500 2185.020 3533.510 ;
        RECT 2362.020 3533.500 2365.020 3533.510 ;
        RECT 2542.020 3533.500 2545.020 3533.510 ;
        RECT 2722.020 3533.500 2725.020 3533.510 ;
        RECT 2902.020 3533.500 2905.020 3533.510 ;
        RECT 2935.800 3533.500 2938.800 3533.510 ;
        RECT -19.180 3530.500 2938.800 3533.500 ;
        RECT -19.180 3530.490 -16.180 3530.500 ;
        RECT 22.020 3530.490 25.020 3530.500 ;
        RECT 202.020 3530.490 205.020 3530.500 ;
        RECT 382.020 3530.490 385.020 3530.500 ;
        RECT 562.020 3530.490 565.020 3530.500 ;
        RECT 742.020 3530.490 745.020 3530.500 ;
        RECT 922.020 3530.490 925.020 3530.500 ;
        RECT 1102.020 3530.490 1105.020 3530.500 ;
        RECT 1282.020 3530.490 1285.020 3530.500 ;
        RECT 1462.020 3530.490 1465.020 3530.500 ;
        RECT 1642.020 3530.490 1645.020 3530.500 ;
        RECT 1822.020 3530.490 1825.020 3530.500 ;
        RECT 2002.020 3530.490 2005.020 3530.500 ;
        RECT 2182.020 3530.490 2185.020 3530.500 ;
        RECT 2362.020 3530.490 2365.020 3530.500 ;
        RECT 2542.020 3530.490 2545.020 3530.500 ;
        RECT 2722.020 3530.490 2725.020 3530.500 ;
        RECT 2902.020 3530.490 2905.020 3530.500 ;
        RECT 2935.800 3530.490 2938.800 3530.500 ;
        RECT -19.180 3450.380 -16.180 3450.390 ;
        RECT 22.020 3450.380 25.020 3450.390 ;
        RECT 202.020 3450.380 205.020 3450.390 ;
        RECT 382.020 3450.380 385.020 3450.390 ;
        RECT 562.020 3450.380 565.020 3450.390 ;
        RECT 742.020 3450.380 745.020 3450.390 ;
        RECT 922.020 3450.380 925.020 3450.390 ;
        RECT 1102.020 3450.380 1105.020 3450.390 ;
        RECT 1282.020 3450.380 1285.020 3450.390 ;
        RECT 1462.020 3450.380 1465.020 3450.390 ;
        RECT 1642.020 3450.380 1645.020 3450.390 ;
        RECT 1822.020 3450.380 1825.020 3450.390 ;
        RECT 2002.020 3450.380 2005.020 3450.390 ;
        RECT 2182.020 3450.380 2185.020 3450.390 ;
        RECT 2362.020 3450.380 2365.020 3450.390 ;
        RECT 2542.020 3450.380 2545.020 3450.390 ;
        RECT 2722.020 3450.380 2725.020 3450.390 ;
        RECT 2902.020 3450.380 2905.020 3450.390 ;
        RECT 2935.800 3450.380 2938.800 3450.390 ;
        RECT -23.780 3447.380 2943.400 3450.380 ;
        RECT -19.180 3447.370 -16.180 3447.380 ;
        RECT 22.020 3447.370 25.020 3447.380 ;
        RECT 202.020 3447.370 205.020 3447.380 ;
        RECT 382.020 3447.370 385.020 3447.380 ;
        RECT 562.020 3447.370 565.020 3447.380 ;
        RECT 742.020 3447.370 745.020 3447.380 ;
        RECT 922.020 3447.370 925.020 3447.380 ;
        RECT 1102.020 3447.370 1105.020 3447.380 ;
        RECT 1282.020 3447.370 1285.020 3447.380 ;
        RECT 1462.020 3447.370 1465.020 3447.380 ;
        RECT 1642.020 3447.370 1645.020 3447.380 ;
        RECT 1822.020 3447.370 1825.020 3447.380 ;
        RECT 2002.020 3447.370 2005.020 3447.380 ;
        RECT 2182.020 3447.370 2185.020 3447.380 ;
        RECT 2362.020 3447.370 2365.020 3447.380 ;
        RECT 2542.020 3447.370 2545.020 3447.380 ;
        RECT 2722.020 3447.370 2725.020 3447.380 ;
        RECT 2902.020 3447.370 2905.020 3447.380 ;
        RECT 2935.800 3447.370 2938.800 3447.380 ;
        RECT -19.180 3270.380 -16.180 3270.390 ;
        RECT 22.020 3270.380 25.020 3270.390 ;
        RECT 202.020 3270.380 205.020 3270.390 ;
        RECT 382.020 3270.380 385.020 3270.390 ;
        RECT 562.020 3270.380 565.020 3270.390 ;
        RECT 742.020 3270.380 745.020 3270.390 ;
        RECT 922.020 3270.380 925.020 3270.390 ;
        RECT 1102.020 3270.380 1105.020 3270.390 ;
        RECT 1282.020 3270.380 1285.020 3270.390 ;
        RECT 1462.020 3270.380 1465.020 3270.390 ;
        RECT 1642.020 3270.380 1645.020 3270.390 ;
        RECT 1822.020 3270.380 1825.020 3270.390 ;
        RECT 2002.020 3270.380 2005.020 3270.390 ;
        RECT 2182.020 3270.380 2185.020 3270.390 ;
        RECT 2362.020 3270.380 2365.020 3270.390 ;
        RECT 2542.020 3270.380 2545.020 3270.390 ;
        RECT 2722.020 3270.380 2725.020 3270.390 ;
        RECT 2902.020 3270.380 2905.020 3270.390 ;
        RECT 2935.800 3270.380 2938.800 3270.390 ;
        RECT -23.780 3267.380 2943.400 3270.380 ;
        RECT -19.180 3267.370 -16.180 3267.380 ;
        RECT 22.020 3267.370 25.020 3267.380 ;
        RECT 202.020 3267.370 205.020 3267.380 ;
        RECT 382.020 3267.370 385.020 3267.380 ;
        RECT 562.020 3267.370 565.020 3267.380 ;
        RECT 742.020 3267.370 745.020 3267.380 ;
        RECT 922.020 3267.370 925.020 3267.380 ;
        RECT 1102.020 3267.370 1105.020 3267.380 ;
        RECT 1282.020 3267.370 1285.020 3267.380 ;
        RECT 1462.020 3267.370 1465.020 3267.380 ;
        RECT 1642.020 3267.370 1645.020 3267.380 ;
        RECT 1822.020 3267.370 1825.020 3267.380 ;
        RECT 2002.020 3267.370 2005.020 3267.380 ;
        RECT 2182.020 3267.370 2185.020 3267.380 ;
        RECT 2362.020 3267.370 2365.020 3267.380 ;
        RECT 2542.020 3267.370 2545.020 3267.380 ;
        RECT 2722.020 3267.370 2725.020 3267.380 ;
        RECT 2902.020 3267.370 2905.020 3267.380 ;
        RECT 2935.800 3267.370 2938.800 3267.380 ;
        RECT -19.180 3090.380 -16.180 3090.390 ;
        RECT 22.020 3090.380 25.020 3090.390 ;
        RECT 202.020 3090.380 205.020 3090.390 ;
        RECT 382.020 3090.380 385.020 3090.390 ;
        RECT 562.020 3090.380 565.020 3090.390 ;
        RECT 742.020 3090.380 745.020 3090.390 ;
        RECT 922.020 3090.380 925.020 3090.390 ;
        RECT 1102.020 3090.380 1105.020 3090.390 ;
        RECT 1282.020 3090.380 1285.020 3090.390 ;
        RECT 1462.020 3090.380 1465.020 3090.390 ;
        RECT 1642.020 3090.380 1645.020 3090.390 ;
        RECT 1822.020 3090.380 1825.020 3090.390 ;
        RECT 2002.020 3090.380 2005.020 3090.390 ;
        RECT 2182.020 3090.380 2185.020 3090.390 ;
        RECT 2362.020 3090.380 2365.020 3090.390 ;
        RECT 2542.020 3090.380 2545.020 3090.390 ;
        RECT 2722.020 3090.380 2725.020 3090.390 ;
        RECT 2902.020 3090.380 2905.020 3090.390 ;
        RECT 2935.800 3090.380 2938.800 3090.390 ;
        RECT -23.780 3087.380 2943.400 3090.380 ;
        RECT -19.180 3087.370 -16.180 3087.380 ;
        RECT 22.020 3087.370 25.020 3087.380 ;
        RECT 202.020 3087.370 205.020 3087.380 ;
        RECT 382.020 3087.370 385.020 3087.380 ;
        RECT 562.020 3087.370 565.020 3087.380 ;
        RECT 742.020 3087.370 745.020 3087.380 ;
        RECT 922.020 3087.370 925.020 3087.380 ;
        RECT 1102.020 3087.370 1105.020 3087.380 ;
        RECT 1282.020 3087.370 1285.020 3087.380 ;
        RECT 1462.020 3087.370 1465.020 3087.380 ;
        RECT 1642.020 3087.370 1645.020 3087.380 ;
        RECT 1822.020 3087.370 1825.020 3087.380 ;
        RECT 2002.020 3087.370 2005.020 3087.380 ;
        RECT 2182.020 3087.370 2185.020 3087.380 ;
        RECT 2362.020 3087.370 2365.020 3087.380 ;
        RECT 2542.020 3087.370 2545.020 3087.380 ;
        RECT 2722.020 3087.370 2725.020 3087.380 ;
        RECT 2902.020 3087.370 2905.020 3087.380 ;
        RECT 2935.800 3087.370 2938.800 3087.380 ;
        RECT -19.180 2910.380 -16.180 2910.390 ;
        RECT 22.020 2910.380 25.020 2910.390 ;
        RECT 202.020 2910.380 205.020 2910.390 ;
        RECT 382.020 2910.380 385.020 2910.390 ;
        RECT 562.020 2910.380 565.020 2910.390 ;
        RECT 742.020 2910.380 745.020 2910.390 ;
        RECT 922.020 2910.380 925.020 2910.390 ;
        RECT 1102.020 2910.380 1105.020 2910.390 ;
        RECT 1282.020 2910.380 1285.020 2910.390 ;
        RECT 1462.020 2910.380 1465.020 2910.390 ;
        RECT 1642.020 2910.380 1645.020 2910.390 ;
        RECT 1822.020 2910.380 1825.020 2910.390 ;
        RECT 2002.020 2910.380 2005.020 2910.390 ;
        RECT 2182.020 2910.380 2185.020 2910.390 ;
        RECT 2362.020 2910.380 2365.020 2910.390 ;
        RECT 2542.020 2910.380 2545.020 2910.390 ;
        RECT 2722.020 2910.380 2725.020 2910.390 ;
        RECT 2902.020 2910.380 2905.020 2910.390 ;
        RECT 2935.800 2910.380 2938.800 2910.390 ;
        RECT -23.780 2907.380 2943.400 2910.380 ;
        RECT -19.180 2907.370 -16.180 2907.380 ;
        RECT 22.020 2907.370 25.020 2907.380 ;
        RECT 202.020 2907.370 205.020 2907.380 ;
        RECT 382.020 2907.370 385.020 2907.380 ;
        RECT 562.020 2907.370 565.020 2907.380 ;
        RECT 742.020 2907.370 745.020 2907.380 ;
        RECT 922.020 2907.370 925.020 2907.380 ;
        RECT 1102.020 2907.370 1105.020 2907.380 ;
        RECT 1282.020 2907.370 1285.020 2907.380 ;
        RECT 1462.020 2907.370 1465.020 2907.380 ;
        RECT 1642.020 2907.370 1645.020 2907.380 ;
        RECT 1822.020 2907.370 1825.020 2907.380 ;
        RECT 2002.020 2907.370 2005.020 2907.380 ;
        RECT 2182.020 2907.370 2185.020 2907.380 ;
        RECT 2362.020 2907.370 2365.020 2907.380 ;
        RECT 2542.020 2907.370 2545.020 2907.380 ;
        RECT 2722.020 2907.370 2725.020 2907.380 ;
        RECT 2902.020 2907.370 2905.020 2907.380 ;
        RECT 2935.800 2907.370 2938.800 2907.380 ;
        RECT -19.180 2730.380 -16.180 2730.390 ;
        RECT 22.020 2730.380 25.020 2730.390 ;
        RECT 202.020 2730.380 205.020 2730.390 ;
        RECT 382.020 2730.380 385.020 2730.390 ;
        RECT 562.020 2730.380 565.020 2730.390 ;
        RECT 742.020 2730.380 745.020 2730.390 ;
        RECT 922.020 2730.380 925.020 2730.390 ;
        RECT 1102.020 2730.380 1105.020 2730.390 ;
        RECT 1282.020 2730.380 1285.020 2730.390 ;
        RECT 1462.020 2730.380 1465.020 2730.390 ;
        RECT 1642.020 2730.380 1645.020 2730.390 ;
        RECT 1822.020 2730.380 1825.020 2730.390 ;
        RECT 2002.020 2730.380 2005.020 2730.390 ;
        RECT 2182.020 2730.380 2185.020 2730.390 ;
        RECT 2362.020 2730.380 2365.020 2730.390 ;
        RECT 2542.020 2730.380 2545.020 2730.390 ;
        RECT 2722.020 2730.380 2725.020 2730.390 ;
        RECT 2902.020 2730.380 2905.020 2730.390 ;
        RECT 2935.800 2730.380 2938.800 2730.390 ;
        RECT -23.780 2727.380 2943.400 2730.380 ;
        RECT -19.180 2727.370 -16.180 2727.380 ;
        RECT 22.020 2727.370 25.020 2727.380 ;
        RECT 202.020 2727.370 205.020 2727.380 ;
        RECT 382.020 2727.370 385.020 2727.380 ;
        RECT 562.020 2727.370 565.020 2727.380 ;
        RECT 742.020 2727.370 745.020 2727.380 ;
        RECT 922.020 2727.370 925.020 2727.380 ;
        RECT 1102.020 2727.370 1105.020 2727.380 ;
        RECT 1282.020 2727.370 1285.020 2727.380 ;
        RECT 1462.020 2727.370 1465.020 2727.380 ;
        RECT 1642.020 2727.370 1645.020 2727.380 ;
        RECT 1822.020 2727.370 1825.020 2727.380 ;
        RECT 2002.020 2727.370 2005.020 2727.380 ;
        RECT 2182.020 2727.370 2185.020 2727.380 ;
        RECT 2362.020 2727.370 2365.020 2727.380 ;
        RECT 2542.020 2727.370 2545.020 2727.380 ;
        RECT 2722.020 2727.370 2725.020 2727.380 ;
        RECT 2902.020 2727.370 2905.020 2727.380 ;
        RECT 2935.800 2727.370 2938.800 2727.380 ;
        RECT -19.180 2550.380 -16.180 2550.390 ;
        RECT 22.020 2550.380 25.020 2550.390 ;
        RECT 202.020 2550.380 205.020 2550.390 ;
        RECT 382.020 2550.380 385.020 2550.390 ;
        RECT 562.020 2550.380 565.020 2550.390 ;
        RECT 742.020 2550.380 745.020 2550.390 ;
        RECT 922.020 2550.380 925.020 2550.390 ;
        RECT 1102.020 2550.380 1105.020 2550.390 ;
        RECT 1282.020 2550.380 1285.020 2550.390 ;
        RECT 1462.020 2550.380 1465.020 2550.390 ;
        RECT 1642.020 2550.380 1645.020 2550.390 ;
        RECT 1822.020 2550.380 1825.020 2550.390 ;
        RECT 2002.020 2550.380 2005.020 2550.390 ;
        RECT 2182.020 2550.380 2185.020 2550.390 ;
        RECT 2362.020 2550.380 2365.020 2550.390 ;
        RECT 2542.020 2550.380 2545.020 2550.390 ;
        RECT 2722.020 2550.380 2725.020 2550.390 ;
        RECT 2902.020 2550.380 2905.020 2550.390 ;
        RECT 2935.800 2550.380 2938.800 2550.390 ;
        RECT -23.780 2547.380 2943.400 2550.380 ;
        RECT -19.180 2547.370 -16.180 2547.380 ;
        RECT 22.020 2547.370 25.020 2547.380 ;
        RECT 202.020 2547.370 205.020 2547.380 ;
        RECT 382.020 2547.370 385.020 2547.380 ;
        RECT 562.020 2547.370 565.020 2547.380 ;
        RECT 742.020 2547.370 745.020 2547.380 ;
        RECT 922.020 2547.370 925.020 2547.380 ;
        RECT 1102.020 2547.370 1105.020 2547.380 ;
        RECT 1282.020 2547.370 1285.020 2547.380 ;
        RECT 1462.020 2547.370 1465.020 2547.380 ;
        RECT 1642.020 2547.370 1645.020 2547.380 ;
        RECT 1822.020 2547.370 1825.020 2547.380 ;
        RECT 2002.020 2547.370 2005.020 2547.380 ;
        RECT 2182.020 2547.370 2185.020 2547.380 ;
        RECT 2362.020 2547.370 2365.020 2547.380 ;
        RECT 2542.020 2547.370 2545.020 2547.380 ;
        RECT 2722.020 2547.370 2725.020 2547.380 ;
        RECT 2902.020 2547.370 2905.020 2547.380 ;
        RECT 2935.800 2547.370 2938.800 2547.380 ;
        RECT -19.180 2370.380 -16.180 2370.390 ;
        RECT 22.020 2370.380 25.020 2370.390 ;
        RECT 202.020 2370.380 205.020 2370.390 ;
        RECT 382.020 2370.380 385.020 2370.390 ;
        RECT 562.020 2370.380 565.020 2370.390 ;
        RECT 742.020 2370.380 745.020 2370.390 ;
        RECT 922.020 2370.380 925.020 2370.390 ;
        RECT 1102.020 2370.380 1105.020 2370.390 ;
        RECT 1282.020 2370.380 1285.020 2370.390 ;
        RECT 1462.020 2370.380 1465.020 2370.390 ;
        RECT 1642.020 2370.380 1645.020 2370.390 ;
        RECT 1822.020 2370.380 1825.020 2370.390 ;
        RECT 2002.020 2370.380 2005.020 2370.390 ;
        RECT 2182.020 2370.380 2185.020 2370.390 ;
        RECT 2362.020 2370.380 2365.020 2370.390 ;
        RECT 2542.020 2370.380 2545.020 2370.390 ;
        RECT 2722.020 2370.380 2725.020 2370.390 ;
        RECT 2902.020 2370.380 2905.020 2370.390 ;
        RECT 2935.800 2370.380 2938.800 2370.390 ;
        RECT -23.780 2367.380 2943.400 2370.380 ;
        RECT -19.180 2367.370 -16.180 2367.380 ;
        RECT 22.020 2367.370 25.020 2367.380 ;
        RECT 202.020 2367.370 205.020 2367.380 ;
        RECT 382.020 2367.370 385.020 2367.380 ;
        RECT 562.020 2367.370 565.020 2367.380 ;
        RECT 742.020 2367.370 745.020 2367.380 ;
        RECT 922.020 2367.370 925.020 2367.380 ;
        RECT 1102.020 2367.370 1105.020 2367.380 ;
        RECT 1282.020 2367.370 1285.020 2367.380 ;
        RECT 1462.020 2367.370 1465.020 2367.380 ;
        RECT 1642.020 2367.370 1645.020 2367.380 ;
        RECT 1822.020 2367.370 1825.020 2367.380 ;
        RECT 2002.020 2367.370 2005.020 2367.380 ;
        RECT 2182.020 2367.370 2185.020 2367.380 ;
        RECT 2362.020 2367.370 2365.020 2367.380 ;
        RECT 2542.020 2367.370 2545.020 2367.380 ;
        RECT 2722.020 2367.370 2725.020 2367.380 ;
        RECT 2902.020 2367.370 2905.020 2367.380 ;
        RECT 2935.800 2367.370 2938.800 2367.380 ;
        RECT -19.180 2190.380 -16.180 2190.390 ;
        RECT 22.020 2190.380 25.020 2190.390 ;
        RECT 202.020 2190.380 205.020 2190.390 ;
        RECT 382.020 2190.380 385.020 2190.390 ;
        RECT 562.020 2190.380 565.020 2190.390 ;
        RECT 742.020 2190.380 745.020 2190.390 ;
        RECT 922.020 2190.380 925.020 2190.390 ;
        RECT 1102.020 2190.380 1105.020 2190.390 ;
        RECT 1282.020 2190.380 1285.020 2190.390 ;
        RECT 1462.020 2190.380 1465.020 2190.390 ;
        RECT 1642.020 2190.380 1645.020 2190.390 ;
        RECT 1822.020 2190.380 1825.020 2190.390 ;
        RECT 2002.020 2190.380 2005.020 2190.390 ;
        RECT 2182.020 2190.380 2185.020 2190.390 ;
        RECT 2362.020 2190.380 2365.020 2190.390 ;
        RECT 2542.020 2190.380 2545.020 2190.390 ;
        RECT 2722.020 2190.380 2725.020 2190.390 ;
        RECT 2902.020 2190.380 2905.020 2190.390 ;
        RECT 2935.800 2190.380 2938.800 2190.390 ;
        RECT -23.780 2187.380 2943.400 2190.380 ;
        RECT -19.180 2187.370 -16.180 2187.380 ;
        RECT 22.020 2187.370 25.020 2187.380 ;
        RECT 202.020 2187.370 205.020 2187.380 ;
        RECT 382.020 2187.370 385.020 2187.380 ;
        RECT 562.020 2187.370 565.020 2187.380 ;
        RECT 742.020 2187.370 745.020 2187.380 ;
        RECT 922.020 2187.370 925.020 2187.380 ;
        RECT 1102.020 2187.370 1105.020 2187.380 ;
        RECT 1282.020 2187.370 1285.020 2187.380 ;
        RECT 1462.020 2187.370 1465.020 2187.380 ;
        RECT 1642.020 2187.370 1645.020 2187.380 ;
        RECT 1822.020 2187.370 1825.020 2187.380 ;
        RECT 2002.020 2187.370 2005.020 2187.380 ;
        RECT 2182.020 2187.370 2185.020 2187.380 ;
        RECT 2362.020 2187.370 2365.020 2187.380 ;
        RECT 2542.020 2187.370 2545.020 2187.380 ;
        RECT 2722.020 2187.370 2725.020 2187.380 ;
        RECT 2902.020 2187.370 2905.020 2187.380 ;
        RECT 2935.800 2187.370 2938.800 2187.380 ;
        RECT -19.180 2010.380 -16.180 2010.390 ;
        RECT 22.020 2010.380 25.020 2010.390 ;
        RECT 202.020 2010.380 205.020 2010.390 ;
        RECT 382.020 2010.380 385.020 2010.390 ;
        RECT 562.020 2010.380 565.020 2010.390 ;
        RECT 742.020 2010.380 745.020 2010.390 ;
        RECT 922.020 2010.380 925.020 2010.390 ;
        RECT 1102.020 2010.380 1105.020 2010.390 ;
        RECT 1282.020 2010.380 1285.020 2010.390 ;
        RECT 1462.020 2010.380 1465.020 2010.390 ;
        RECT 1642.020 2010.380 1645.020 2010.390 ;
        RECT 1822.020 2010.380 1825.020 2010.390 ;
        RECT 2002.020 2010.380 2005.020 2010.390 ;
        RECT 2182.020 2010.380 2185.020 2010.390 ;
        RECT 2362.020 2010.380 2365.020 2010.390 ;
        RECT 2542.020 2010.380 2545.020 2010.390 ;
        RECT 2722.020 2010.380 2725.020 2010.390 ;
        RECT 2902.020 2010.380 2905.020 2010.390 ;
        RECT 2935.800 2010.380 2938.800 2010.390 ;
        RECT -23.780 2007.380 2943.400 2010.380 ;
        RECT -19.180 2007.370 -16.180 2007.380 ;
        RECT 22.020 2007.370 25.020 2007.380 ;
        RECT 202.020 2007.370 205.020 2007.380 ;
        RECT 382.020 2007.370 385.020 2007.380 ;
        RECT 562.020 2007.370 565.020 2007.380 ;
        RECT 742.020 2007.370 745.020 2007.380 ;
        RECT 922.020 2007.370 925.020 2007.380 ;
        RECT 1102.020 2007.370 1105.020 2007.380 ;
        RECT 1282.020 2007.370 1285.020 2007.380 ;
        RECT 1462.020 2007.370 1465.020 2007.380 ;
        RECT 1642.020 2007.370 1645.020 2007.380 ;
        RECT 1822.020 2007.370 1825.020 2007.380 ;
        RECT 2002.020 2007.370 2005.020 2007.380 ;
        RECT 2182.020 2007.370 2185.020 2007.380 ;
        RECT 2362.020 2007.370 2365.020 2007.380 ;
        RECT 2542.020 2007.370 2545.020 2007.380 ;
        RECT 2722.020 2007.370 2725.020 2007.380 ;
        RECT 2902.020 2007.370 2905.020 2007.380 ;
        RECT 2935.800 2007.370 2938.800 2007.380 ;
        RECT -19.180 1830.380 -16.180 1830.390 ;
        RECT 22.020 1830.380 25.020 1830.390 ;
        RECT 202.020 1830.380 205.020 1830.390 ;
        RECT 382.020 1830.380 385.020 1830.390 ;
        RECT 562.020 1830.380 565.020 1830.390 ;
        RECT 742.020 1830.380 745.020 1830.390 ;
        RECT 922.020 1830.380 925.020 1830.390 ;
        RECT 1102.020 1830.380 1105.020 1830.390 ;
        RECT 1282.020 1830.380 1285.020 1830.390 ;
        RECT 1462.020 1830.380 1465.020 1830.390 ;
        RECT 1642.020 1830.380 1645.020 1830.390 ;
        RECT 1822.020 1830.380 1825.020 1830.390 ;
        RECT 2002.020 1830.380 2005.020 1830.390 ;
        RECT 2182.020 1830.380 2185.020 1830.390 ;
        RECT 2362.020 1830.380 2365.020 1830.390 ;
        RECT 2542.020 1830.380 2545.020 1830.390 ;
        RECT 2722.020 1830.380 2725.020 1830.390 ;
        RECT 2902.020 1830.380 2905.020 1830.390 ;
        RECT 2935.800 1830.380 2938.800 1830.390 ;
        RECT -23.780 1827.380 2943.400 1830.380 ;
        RECT -19.180 1827.370 -16.180 1827.380 ;
        RECT 22.020 1827.370 25.020 1827.380 ;
        RECT 202.020 1827.370 205.020 1827.380 ;
        RECT 382.020 1827.370 385.020 1827.380 ;
        RECT 562.020 1827.370 565.020 1827.380 ;
        RECT 742.020 1827.370 745.020 1827.380 ;
        RECT 922.020 1827.370 925.020 1827.380 ;
        RECT 1102.020 1827.370 1105.020 1827.380 ;
        RECT 1282.020 1827.370 1285.020 1827.380 ;
        RECT 1462.020 1827.370 1465.020 1827.380 ;
        RECT 1642.020 1827.370 1645.020 1827.380 ;
        RECT 1822.020 1827.370 1825.020 1827.380 ;
        RECT 2002.020 1827.370 2005.020 1827.380 ;
        RECT 2182.020 1827.370 2185.020 1827.380 ;
        RECT 2362.020 1827.370 2365.020 1827.380 ;
        RECT 2542.020 1827.370 2545.020 1827.380 ;
        RECT 2722.020 1827.370 2725.020 1827.380 ;
        RECT 2902.020 1827.370 2905.020 1827.380 ;
        RECT 2935.800 1827.370 2938.800 1827.380 ;
        RECT -19.180 1650.380 -16.180 1650.390 ;
        RECT 22.020 1650.380 25.020 1650.390 ;
        RECT 202.020 1650.380 205.020 1650.390 ;
        RECT 382.020 1650.380 385.020 1650.390 ;
        RECT 562.020 1650.380 565.020 1650.390 ;
        RECT 742.020 1650.380 745.020 1650.390 ;
        RECT 922.020 1650.380 925.020 1650.390 ;
        RECT 1102.020 1650.380 1105.020 1650.390 ;
        RECT 1282.020 1650.380 1285.020 1650.390 ;
        RECT 1462.020 1650.380 1465.020 1650.390 ;
        RECT 1642.020 1650.380 1645.020 1650.390 ;
        RECT 1822.020 1650.380 1825.020 1650.390 ;
        RECT 2002.020 1650.380 2005.020 1650.390 ;
        RECT 2182.020 1650.380 2185.020 1650.390 ;
        RECT 2362.020 1650.380 2365.020 1650.390 ;
        RECT 2542.020 1650.380 2545.020 1650.390 ;
        RECT 2722.020 1650.380 2725.020 1650.390 ;
        RECT 2902.020 1650.380 2905.020 1650.390 ;
        RECT 2935.800 1650.380 2938.800 1650.390 ;
        RECT -23.780 1647.380 2943.400 1650.380 ;
        RECT -19.180 1647.370 -16.180 1647.380 ;
        RECT 22.020 1647.370 25.020 1647.380 ;
        RECT 202.020 1647.370 205.020 1647.380 ;
        RECT 382.020 1647.370 385.020 1647.380 ;
        RECT 562.020 1647.370 565.020 1647.380 ;
        RECT 742.020 1647.370 745.020 1647.380 ;
        RECT 922.020 1647.370 925.020 1647.380 ;
        RECT 1102.020 1647.370 1105.020 1647.380 ;
        RECT 1282.020 1647.370 1285.020 1647.380 ;
        RECT 1462.020 1647.370 1465.020 1647.380 ;
        RECT 1642.020 1647.370 1645.020 1647.380 ;
        RECT 1822.020 1647.370 1825.020 1647.380 ;
        RECT 2002.020 1647.370 2005.020 1647.380 ;
        RECT 2182.020 1647.370 2185.020 1647.380 ;
        RECT 2362.020 1647.370 2365.020 1647.380 ;
        RECT 2542.020 1647.370 2545.020 1647.380 ;
        RECT 2722.020 1647.370 2725.020 1647.380 ;
        RECT 2902.020 1647.370 2905.020 1647.380 ;
        RECT 2935.800 1647.370 2938.800 1647.380 ;
        RECT -19.180 1470.380 -16.180 1470.390 ;
        RECT 22.020 1470.380 25.020 1470.390 ;
        RECT 202.020 1470.380 205.020 1470.390 ;
        RECT 382.020 1470.380 385.020 1470.390 ;
        RECT 562.020 1470.380 565.020 1470.390 ;
        RECT 742.020 1470.380 745.020 1470.390 ;
        RECT 922.020 1470.380 925.020 1470.390 ;
        RECT 1102.020 1470.380 1105.020 1470.390 ;
        RECT 1282.020 1470.380 1285.020 1470.390 ;
        RECT 1462.020 1470.380 1465.020 1470.390 ;
        RECT 1642.020 1470.380 1645.020 1470.390 ;
        RECT 1822.020 1470.380 1825.020 1470.390 ;
        RECT 2002.020 1470.380 2005.020 1470.390 ;
        RECT 2182.020 1470.380 2185.020 1470.390 ;
        RECT 2362.020 1470.380 2365.020 1470.390 ;
        RECT 2542.020 1470.380 2545.020 1470.390 ;
        RECT 2722.020 1470.380 2725.020 1470.390 ;
        RECT 2902.020 1470.380 2905.020 1470.390 ;
        RECT 2935.800 1470.380 2938.800 1470.390 ;
        RECT -23.780 1467.380 2943.400 1470.380 ;
        RECT -19.180 1467.370 -16.180 1467.380 ;
        RECT 22.020 1467.370 25.020 1467.380 ;
        RECT 202.020 1467.370 205.020 1467.380 ;
        RECT 382.020 1467.370 385.020 1467.380 ;
        RECT 562.020 1467.370 565.020 1467.380 ;
        RECT 742.020 1467.370 745.020 1467.380 ;
        RECT 922.020 1467.370 925.020 1467.380 ;
        RECT 1102.020 1467.370 1105.020 1467.380 ;
        RECT 1282.020 1467.370 1285.020 1467.380 ;
        RECT 1462.020 1467.370 1465.020 1467.380 ;
        RECT 1642.020 1467.370 1645.020 1467.380 ;
        RECT 1822.020 1467.370 1825.020 1467.380 ;
        RECT 2002.020 1467.370 2005.020 1467.380 ;
        RECT 2182.020 1467.370 2185.020 1467.380 ;
        RECT 2362.020 1467.370 2365.020 1467.380 ;
        RECT 2542.020 1467.370 2545.020 1467.380 ;
        RECT 2722.020 1467.370 2725.020 1467.380 ;
        RECT 2902.020 1467.370 2905.020 1467.380 ;
        RECT 2935.800 1467.370 2938.800 1467.380 ;
        RECT -19.180 1290.380 -16.180 1290.390 ;
        RECT 22.020 1290.380 25.020 1290.390 ;
        RECT 202.020 1290.380 205.020 1290.390 ;
        RECT 382.020 1290.380 385.020 1290.390 ;
        RECT 562.020 1290.380 565.020 1290.390 ;
        RECT 742.020 1290.380 745.020 1290.390 ;
        RECT 922.020 1290.380 925.020 1290.390 ;
        RECT 1102.020 1290.380 1105.020 1290.390 ;
        RECT 1282.020 1290.380 1285.020 1290.390 ;
        RECT 1462.020 1290.380 1465.020 1290.390 ;
        RECT 1642.020 1290.380 1645.020 1290.390 ;
        RECT 1822.020 1290.380 1825.020 1290.390 ;
        RECT 2002.020 1290.380 2005.020 1290.390 ;
        RECT 2182.020 1290.380 2185.020 1290.390 ;
        RECT 2362.020 1290.380 2365.020 1290.390 ;
        RECT 2542.020 1290.380 2545.020 1290.390 ;
        RECT 2722.020 1290.380 2725.020 1290.390 ;
        RECT 2902.020 1290.380 2905.020 1290.390 ;
        RECT 2935.800 1290.380 2938.800 1290.390 ;
        RECT -23.780 1287.380 2943.400 1290.380 ;
        RECT -19.180 1287.370 -16.180 1287.380 ;
        RECT 22.020 1287.370 25.020 1287.380 ;
        RECT 202.020 1287.370 205.020 1287.380 ;
        RECT 382.020 1287.370 385.020 1287.380 ;
        RECT 562.020 1287.370 565.020 1287.380 ;
        RECT 742.020 1287.370 745.020 1287.380 ;
        RECT 922.020 1287.370 925.020 1287.380 ;
        RECT 1102.020 1287.370 1105.020 1287.380 ;
        RECT 1282.020 1287.370 1285.020 1287.380 ;
        RECT 1462.020 1287.370 1465.020 1287.380 ;
        RECT 1642.020 1287.370 1645.020 1287.380 ;
        RECT 1822.020 1287.370 1825.020 1287.380 ;
        RECT 2002.020 1287.370 2005.020 1287.380 ;
        RECT 2182.020 1287.370 2185.020 1287.380 ;
        RECT 2362.020 1287.370 2365.020 1287.380 ;
        RECT 2542.020 1287.370 2545.020 1287.380 ;
        RECT 2722.020 1287.370 2725.020 1287.380 ;
        RECT 2902.020 1287.370 2905.020 1287.380 ;
        RECT 2935.800 1287.370 2938.800 1287.380 ;
        RECT -19.180 1110.380 -16.180 1110.390 ;
        RECT 22.020 1110.380 25.020 1110.390 ;
        RECT 202.020 1110.380 205.020 1110.390 ;
        RECT 382.020 1110.380 385.020 1110.390 ;
        RECT 562.020 1110.380 565.020 1110.390 ;
        RECT 742.020 1110.380 745.020 1110.390 ;
        RECT 922.020 1110.380 925.020 1110.390 ;
        RECT 1102.020 1110.380 1105.020 1110.390 ;
        RECT 1282.020 1110.380 1285.020 1110.390 ;
        RECT 1462.020 1110.380 1465.020 1110.390 ;
        RECT 1642.020 1110.380 1645.020 1110.390 ;
        RECT 1822.020 1110.380 1825.020 1110.390 ;
        RECT 2002.020 1110.380 2005.020 1110.390 ;
        RECT 2182.020 1110.380 2185.020 1110.390 ;
        RECT 2362.020 1110.380 2365.020 1110.390 ;
        RECT 2542.020 1110.380 2545.020 1110.390 ;
        RECT 2722.020 1110.380 2725.020 1110.390 ;
        RECT 2902.020 1110.380 2905.020 1110.390 ;
        RECT 2935.800 1110.380 2938.800 1110.390 ;
        RECT -23.780 1107.380 2943.400 1110.380 ;
        RECT -19.180 1107.370 -16.180 1107.380 ;
        RECT 22.020 1107.370 25.020 1107.380 ;
        RECT 202.020 1107.370 205.020 1107.380 ;
        RECT 382.020 1107.370 385.020 1107.380 ;
        RECT 562.020 1107.370 565.020 1107.380 ;
        RECT 742.020 1107.370 745.020 1107.380 ;
        RECT 922.020 1107.370 925.020 1107.380 ;
        RECT 1102.020 1107.370 1105.020 1107.380 ;
        RECT 1282.020 1107.370 1285.020 1107.380 ;
        RECT 1462.020 1107.370 1465.020 1107.380 ;
        RECT 1642.020 1107.370 1645.020 1107.380 ;
        RECT 1822.020 1107.370 1825.020 1107.380 ;
        RECT 2002.020 1107.370 2005.020 1107.380 ;
        RECT 2182.020 1107.370 2185.020 1107.380 ;
        RECT 2362.020 1107.370 2365.020 1107.380 ;
        RECT 2542.020 1107.370 2545.020 1107.380 ;
        RECT 2722.020 1107.370 2725.020 1107.380 ;
        RECT 2902.020 1107.370 2905.020 1107.380 ;
        RECT 2935.800 1107.370 2938.800 1107.380 ;
        RECT -19.180 930.380 -16.180 930.390 ;
        RECT 22.020 930.380 25.020 930.390 ;
        RECT 202.020 930.380 205.020 930.390 ;
        RECT 382.020 930.380 385.020 930.390 ;
        RECT 562.020 930.380 565.020 930.390 ;
        RECT 742.020 930.380 745.020 930.390 ;
        RECT 922.020 930.380 925.020 930.390 ;
        RECT 1102.020 930.380 1105.020 930.390 ;
        RECT 1282.020 930.380 1285.020 930.390 ;
        RECT 1462.020 930.380 1465.020 930.390 ;
        RECT 1642.020 930.380 1645.020 930.390 ;
        RECT 1822.020 930.380 1825.020 930.390 ;
        RECT 2002.020 930.380 2005.020 930.390 ;
        RECT 2182.020 930.380 2185.020 930.390 ;
        RECT 2362.020 930.380 2365.020 930.390 ;
        RECT 2542.020 930.380 2545.020 930.390 ;
        RECT 2722.020 930.380 2725.020 930.390 ;
        RECT 2902.020 930.380 2905.020 930.390 ;
        RECT 2935.800 930.380 2938.800 930.390 ;
        RECT -23.780 927.380 2943.400 930.380 ;
        RECT -19.180 927.370 -16.180 927.380 ;
        RECT 22.020 927.370 25.020 927.380 ;
        RECT 202.020 927.370 205.020 927.380 ;
        RECT 382.020 927.370 385.020 927.380 ;
        RECT 562.020 927.370 565.020 927.380 ;
        RECT 742.020 927.370 745.020 927.380 ;
        RECT 922.020 927.370 925.020 927.380 ;
        RECT 1102.020 927.370 1105.020 927.380 ;
        RECT 1282.020 927.370 1285.020 927.380 ;
        RECT 1462.020 927.370 1465.020 927.380 ;
        RECT 1642.020 927.370 1645.020 927.380 ;
        RECT 1822.020 927.370 1825.020 927.380 ;
        RECT 2002.020 927.370 2005.020 927.380 ;
        RECT 2182.020 927.370 2185.020 927.380 ;
        RECT 2362.020 927.370 2365.020 927.380 ;
        RECT 2542.020 927.370 2545.020 927.380 ;
        RECT 2722.020 927.370 2725.020 927.380 ;
        RECT 2902.020 927.370 2905.020 927.380 ;
        RECT 2935.800 927.370 2938.800 927.380 ;
        RECT -19.180 750.380 -16.180 750.390 ;
        RECT 22.020 750.380 25.020 750.390 ;
        RECT 202.020 750.380 205.020 750.390 ;
        RECT 382.020 750.380 385.020 750.390 ;
        RECT 562.020 750.380 565.020 750.390 ;
        RECT 742.020 750.380 745.020 750.390 ;
        RECT 922.020 750.380 925.020 750.390 ;
        RECT 1102.020 750.380 1105.020 750.390 ;
        RECT 1282.020 750.380 1285.020 750.390 ;
        RECT 1462.020 750.380 1465.020 750.390 ;
        RECT 1642.020 750.380 1645.020 750.390 ;
        RECT 1822.020 750.380 1825.020 750.390 ;
        RECT 2002.020 750.380 2005.020 750.390 ;
        RECT 2182.020 750.380 2185.020 750.390 ;
        RECT 2362.020 750.380 2365.020 750.390 ;
        RECT 2542.020 750.380 2545.020 750.390 ;
        RECT 2722.020 750.380 2725.020 750.390 ;
        RECT 2902.020 750.380 2905.020 750.390 ;
        RECT 2935.800 750.380 2938.800 750.390 ;
        RECT -23.780 747.380 2943.400 750.380 ;
        RECT -19.180 747.370 -16.180 747.380 ;
        RECT 22.020 747.370 25.020 747.380 ;
        RECT 202.020 747.370 205.020 747.380 ;
        RECT 382.020 747.370 385.020 747.380 ;
        RECT 562.020 747.370 565.020 747.380 ;
        RECT 742.020 747.370 745.020 747.380 ;
        RECT 922.020 747.370 925.020 747.380 ;
        RECT 1102.020 747.370 1105.020 747.380 ;
        RECT 1282.020 747.370 1285.020 747.380 ;
        RECT 1462.020 747.370 1465.020 747.380 ;
        RECT 1642.020 747.370 1645.020 747.380 ;
        RECT 1822.020 747.370 1825.020 747.380 ;
        RECT 2002.020 747.370 2005.020 747.380 ;
        RECT 2182.020 747.370 2185.020 747.380 ;
        RECT 2362.020 747.370 2365.020 747.380 ;
        RECT 2542.020 747.370 2545.020 747.380 ;
        RECT 2722.020 747.370 2725.020 747.380 ;
        RECT 2902.020 747.370 2905.020 747.380 ;
        RECT 2935.800 747.370 2938.800 747.380 ;
        RECT -19.180 570.380 -16.180 570.390 ;
        RECT 22.020 570.380 25.020 570.390 ;
        RECT 202.020 570.380 205.020 570.390 ;
        RECT 382.020 570.380 385.020 570.390 ;
        RECT 562.020 570.380 565.020 570.390 ;
        RECT 742.020 570.380 745.020 570.390 ;
        RECT 922.020 570.380 925.020 570.390 ;
        RECT 1102.020 570.380 1105.020 570.390 ;
        RECT 1282.020 570.380 1285.020 570.390 ;
        RECT 1462.020 570.380 1465.020 570.390 ;
        RECT 1642.020 570.380 1645.020 570.390 ;
        RECT 1822.020 570.380 1825.020 570.390 ;
        RECT 2002.020 570.380 2005.020 570.390 ;
        RECT 2182.020 570.380 2185.020 570.390 ;
        RECT 2362.020 570.380 2365.020 570.390 ;
        RECT 2542.020 570.380 2545.020 570.390 ;
        RECT 2722.020 570.380 2725.020 570.390 ;
        RECT 2902.020 570.380 2905.020 570.390 ;
        RECT 2935.800 570.380 2938.800 570.390 ;
        RECT -23.780 567.380 2943.400 570.380 ;
        RECT -19.180 567.370 -16.180 567.380 ;
        RECT 22.020 567.370 25.020 567.380 ;
        RECT 202.020 567.370 205.020 567.380 ;
        RECT 382.020 567.370 385.020 567.380 ;
        RECT 562.020 567.370 565.020 567.380 ;
        RECT 742.020 567.370 745.020 567.380 ;
        RECT 922.020 567.370 925.020 567.380 ;
        RECT 1102.020 567.370 1105.020 567.380 ;
        RECT 1282.020 567.370 1285.020 567.380 ;
        RECT 1462.020 567.370 1465.020 567.380 ;
        RECT 1642.020 567.370 1645.020 567.380 ;
        RECT 1822.020 567.370 1825.020 567.380 ;
        RECT 2002.020 567.370 2005.020 567.380 ;
        RECT 2182.020 567.370 2185.020 567.380 ;
        RECT 2362.020 567.370 2365.020 567.380 ;
        RECT 2542.020 567.370 2545.020 567.380 ;
        RECT 2722.020 567.370 2725.020 567.380 ;
        RECT 2902.020 567.370 2905.020 567.380 ;
        RECT 2935.800 567.370 2938.800 567.380 ;
        RECT -19.180 390.380 -16.180 390.390 ;
        RECT 22.020 390.380 25.020 390.390 ;
        RECT 202.020 390.380 205.020 390.390 ;
        RECT 382.020 390.380 385.020 390.390 ;
        RECT 562.020 390.380 565.020 390.390 ;
        RECT 742.020 390.380 745.020 390.390 ;
        RECT 922.020 390.380 925.020 390.390 ;
        RECT 1102.020 390.380 1105.020 390.390 ;
        RECT 1282.020 390.380 1285.020 390.390 ;
        RECT 1462.020 390.380 1465.020 390.390 ;
        RECT 1642.020 390.380 1645.020 390.390 ;
        RECT 1822.020 390.380 1825.020 390.390 ;
        RECT 2002.020 390.380 2005.020 390.390 ;
        RECT 2182.020 390.380 2185.020 390.390 ;
        RECT 2362.020 390.380 2365.020 390.390 ;
        RECT 2542.020 390.380 2545.020 390.390 ;
        RECT 2722.020 390.380 2725.020 390.390 ;
        RECT 2902.020 390.380 2905.020 390.390 ;
        RECT 2935.800 390.380 2938.800 390.390 ;
        RECT -23.780 387.380 2943.400 390.380 ;
        RECT -19.180 387.370 -16.180 387.380 ;
        RECT 22.020 387.370 25.020 387.380 ;
        RECT 202.020 387.370 205.020 387.380 ;
        RECT 382.020 387.370 385.020 387.380 ;
        RECT 562.020 387.370 565.020 387.380 ;
        RECT 742.020 387.370 745.020 387.380 ;
        RECT 922.020 387.370 925.020 387.380 ;
        RECT 1102.020 387.370 1105.020 387.380 ;
        RECT 1282.020 387.370 1285.020 387.380 ;
        RECT 1462.020 387.370 1465.020 387.380 ;
        RECT 1642.020 387.370 1645.020 387.380 ;
        RECT 1822.020 387.370 1825.020 387.380 ;
        RECT 2002.020 387.370 2005.020 387.380 ;
        RECT 2182.020 387.370 2185.020 387.380 ;
        RECT 2362.020 387.370 2365.020 387.380 ;
        RECT 2542.020 387.370 2545.020 387.380 ;
        RECT 2722.020 387.370 2725.020 387.380 ;
        RECT 2902.020 387.370 2905.020 387.380 ;
        RECT 2935.800 387.370 2938.800 387.380 ;
        RECT -19.180 210.380 -16.180 210.390 ;
        RECT 22.020 210.380 25.020 210.390 ;
        RECT 202.020 210.380 205.020 210.390 ;
        RECT 382.020 210.380 385.020 210.390 ;
        RECT 562.020 210.380 565.020 210.390 ;
        RECT 742.020 210.380 745.020 210.390 ;
        RECT 922.020 210.380 925.020 210.390 ;
        RECT 1102.020 210.380 1105.020 210.390 ;
        RECT 1282.020 210.380 1285.020 210.390 ;
        RECT 1462.020 210.380 1465.020 210.390 ;
        RECT 1642.020 210.380 1645.020 210.390 ;
        RECT 1822.020 210.380 1825.020 210.390 ;
        RECT 2002.020 210.380 2005.020 210.390 ;
        RECT 2182.020 210.380 2185.020 210.390 ;
        RECT 2362.020 210.380 2365.020 210.390 ;
        RECT 2542.020 210.380 2545.020 210.390 ;
        RECT 2722.020 210.380 2725.020 210.390 ;
        RECT 2902.020 210.380 2905.020 210.390 ;
        RECT 2935.800 210.380 2938.800 210.390 ;
        RECT -23.780 207.380 2943.400 210.380 ;
        RECT -19.180 207.370 -16.180 207.380 ;
        RECT 22.020 207.370 25.020 207.380 ;
        RECT 202.020 207.370 205.020 207.380 ;
        RECT 382.020 207.370 385.020 207.380 ;
        RECT 562.020 207.370 565.020 207.380 ;
        RECT 742.020 207.370 745.020 207.380 ;
        RECT 922.020 207.370 925.020 207.380 ;
        RECT 1102.020 207.370 1105.020 207.380 ;
        RECT 1282.020 207.370 1285.020 207.380 ;
        RECT 1462.020 207.370 1465.020 207.380 ;
        RECT 1642.020 207.370 1645.020 207.380 ;
        RECT 1822.020 207.370 1825.020 207.380 ;
        RECT 2002.020 207.370 2005.020 207.380 ;
        RECT 2182.020 207.370 2185.020 207.380 ;
        RECT 2362.020 207.370 2365.020 207.380 ;
        RECT 2542.020 207.370 2545.020 207.380 ;
        RECT 2722.020 207.370 2725.020 207.380 ;
        RECT 2902.020 207.370 2905.020 207.380 ;
        RECT 2935.800 207.370 2938.800 207.380 ;
        RECT -19.180 30.380 -16.180 30.390 ;
        RECT 22.020 30.380 25.020 30.390 ;
        RECT 202.020 30.380 205.020 30.390 ;
        RECT 382.020 30.380 385.020 30.390 ;
        RECT 562.020 30.380 565.020 30.390 ;
        RECT 742.020 30.380 745.020 30.390 ;
        RECT 922.020 30.380 925.020 30.390 ;
        RECT 1102.020 30.380 1105.020 30.390 ;
        RECT 1282.020 30.380 1285.020 30.390 ;
        RECT 1462.020 30.380 1465.020 30.390 ;
        RECT 1642.020 30.380 1645.020 30.390 ;
        RECT 1822.020 30.380 1825.020 30.390 ;
        RECT 2002.020 30.380 2005.020 30.390 ;
        RECT 2182.020 30.380 2185.020 30.390 ;
        RECT 2362.020 30.380 2365.020 30.390 ;
        RECT 2542.020 30.380 2545.020 30.390 ;
        RECT 2722.020 30.380 2725.020 30.390 ;
        RECT 2902.020 30.380 2905.020 30.390 ;
        RECT 2935.800 30.380 2938.800 30.390 ;
        RECT -23.780 27.380 2943.400 30.380 ;
        RECT -19.180 27.370 -16.180 27.380 ;
        RECT 22.020 27.370 25.020 27.380 ;
        RECT 202.020 27.370 205.020 27.380 ;
        RECT 382.020 27.370 385.020 27.380 ;
        RECT 562.020 27.370 565.020 27.380 ;
        RECT 742.020 27.370 745.020 27.380 ;
        RECT 922.020 27.370 925.020 27.380 ;
        RECT 1102.020 27.370 1105.020 27.380 ;
        RECT 1282.020 27.370 1285.020 27.380 ;
        RECT 1462.020 27.370 1465.020 27.380 ;
        RECT 1642.020 27.370 1645.020 27.380 ;
        RECT 1822.020 27.370 1825.020 27.380 ;
        RECT 2002.020 27.370 2005.020 27.380 ;
        RECT 2182.020 27.370 2185.020 27.380 ;
        RECT 2362.020 27.370 2365.020 27.380 ;
        RECT 2542.020 27.370 2545.020 27.380 ;
        RECT 2722.020 27.370 2725.020 27.380 ;
        RECT 2902.020 27.370 2905.020 27.380 ;
        RECT 2935.800 27.370 2938.800 27.380 ;
        RECT -19.180 -10.820 -16.180 -10.810 ;
        RECT 22.020 -10.820 25.020 -10.810 ;
        RECT 202.020 -10.820 205.020 -10.810 ;
        RECT 382.020 -10.820 385.020 -10.810 ;
        RECT 562.020 -10.820 565.020 -10.810 ;
        RECT 742.020 -10.820 745.020 -10.810 ;
        RECT 922.020 -10.820 925.020 -10.810 ;
        RECT 1102.020 -10.820 1105.020 -10.810 ;
        RECT 1282.020 -10.820 1285.020 -10.810 ;
        RECT 1462.020 -10.820 1465.020 -10.810 ;
        RECT 1642.020 -10.820 1645.020 -10.810 ;
        RECT 1822.020 -10.820 1825.020 -10.810 ;
        RECT 2002.020 -10.820 2005.020 -10.810 ;
        RECT 2182.020 -10.820 2185.020 -10.810 ;
        RECT 2362.020 -10.820 2365.020 -10.810 ;
        RECT 2542.020 -10.820 2545.020 -10.810 ;
        RECT 2722.020 -10.820 2725.020 -10.810 ;
        RECT 2902.020 -10.820 2905.020 -10.810 ;
        RECT 2935.800 -10.820 2938.800 -10.810 ;
        RECT -19.180 -13.820 2938.800 -10.820 ;
        RECT -19.180 -13.830 -16.180 -13.820 ;
        RECT 22.020 -13.830 25.020 -13.820 ;
        RECT 202.020 -13.830 205.020 -13.820 ;
        RECT 382.020 -13.830 385.020 -13.820 ;
        RECT 562.020 -13.830 565.020 -13.820 ;
        RECT 742.020 -13.830 745.020 -13.820 ;
        RECT 922.020 -13.830 925.020 -13.820 ;
        RECT 1102.020 -13.830 1105.020 -13.820 ;
        RECT 1282.020 -13.830 1285.020 -13.820 ;
        RECT 1462.020 -13.830 1465.020 -13.820 ;
        RECT 1642.020 -13.830 1645.020 -13.820 ;
        RECT 1822.020 -13.830 1825.020 -13.820 ;
        RECT 2002.020 -13.830 2005.020 -13.820 ;
        RECT 2182.020 -13.830 2185.020 -13.820 ;
        RECT 2362.020 -13.830 2365.020 -13.820 ;
        RECT 2542.020 -13.830 2545.020 -13.820 ;
        RECT 2722.020 -13.830 2725.020 -13.820 ;
        RECT 2902.020 -13.830 2905.020 -13.820 ;
        RECT 2935.800 -13.830 2938.800 -13.820 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -23.780 -18.420 -20.780 3538.100 ;
        RECT 112.020 -18.420 115.020 3538.100 ;
        RECT 292.020 -18.420 295.020 3538.100 ;
        RECT 472.020 -18.420 475.020 3538.100 ;
        RECT 652.020 -18.420 655.020 3538.100 ;
        RECT 832.020 -18.420 835.020 3538.100 ;
        RECT 1012.020 -18.420 1015.020 3538.100 ;
        RECT 1192.020 -18.420 1195.020 3538.100 ;
        RECT 1372.020 -18.420 1375.020 3538.100 ;
        RECT 1552.020 -18.420 1555.020 3538.100 ;
        RECT 1732.020 -18.420 1735.020 3538.100 ;
        RECT 1912.020 -18.420 1915.020 3538.100 ;
        RECT 2092.020 -18.420 2095.020 3538.100 ;
        RECT 2272.020 -18.420 2275.020 3538.100 ;
        RECT 2452.020 -18.420 2455.020 3538.100 ;
        RECT 2632.020 -18.420 2635.020 3538.100 ;
        RECT 2812.020 -18.420 2815.020 3538.100 ;
        RECT 2940.400 -18.420 2943.400 3538.100 ;
      LAYER via4 ;
        RECT -22.870 3536.810 -21.690 3537.990 ;
        RECT -22.870 3535.210 -21.690 3536.390 ;
        RECT -22.870 3359.090 -21.690 3360.270 ;
        RECT -22.870 3357.490 -21.690 3358.670 ;
        RECT -22.870 3179.090 -21.690 3180.270 ;
        RECT -22.870 3177.490 -21.690 3178.670 ;
        RECT -22.870 2999.090 -21.690 3000.270 ;
        RECT -22.870 2997.490 -21.690 2998.670 ;
        RECT -22.870 2819.090 -21.690 2820.270 ;
        RECT -22.870 2817.490 -21.690 2818.670 ;
        RECT -22.870 2639.090 -21.690 2640.270 ;
        RECT -22.870 2637.490 -21.690 2638.670 ;
        RECT -22.870 2459.090 -21.690 2460.270 ;
        RECT -22.870 2457.490 -21.690 2458.670 ;
        RECT -22.870 2279.090 -21.690 2280.270 ;
        RECT -22.870 2277.490 -21.690 2278.670 ;
        RECT -22.870 2099.090 -21.690 2100.270 ;
        RECT -22.870 2097.490 -21.690 2098.670 ;
        RECT -22.870 1919.090 -21.690 1920.270 ;
        RECT -22.870 1917.490 -21.690 1918.670 ;
        RECT -22.870 1739.090 -21.690 1740.270 ;
        RECT -22.870 1737.490 -21.690 1738.670 ;
        RECT -22.870 1559.090 -21.690 1560.270 ;
        RECT -22.870 1557.490 -21.690 1558.670 ;
        RECT -22.870 1379.090 -21.690 1380.270 ;
        RECT -22.870 1377.490 -21.690 1378.670 ;
        RECT -22.870 1199.090 -21.690 1200.270 ;
        RECT -22.870 1197.490 -21.690 1198.670 ;
        RECT -22.870 1019.090 -21.690 1020.270 ;
        RECT -22.870 1017.490 -21.690 1018.670 ;
        RECT -22.870 839.090 -21.690 840.270 ;
        RECT -22.870 837.490 -21.690 838.670 ;
        RECT -22.870 659.090 -21.690 660.270 ;
        RECT -22.870 657.490 -21.690 658.670 ;
        RECT -22.870 479.090 -21.690 480.270 ;
        RECT -22.870 477.490 -21.690 478.670 ;
        RECT -22.870 299.090 -21.690 300.270 ;
        RECT -22.870 297.490 -21.690 298.670 ;
        RECT -22.870 119.090 -21.690 120.270 ;
        RECT -22.870 117.490 -21.690 118.670 ;
        RECT -22.870 -16.710 -21.690 -15.530 ;
        RECT -22.870 -18.310 -21.690 -17.130 ;
        RECT 112.930 3536.810 114.110 3537.990 ;
        RECT 112.930 3535.210 114.110 3536.390 ;
        RECT 112.930 3359.090 114.110 3360.270 ;
        RECT 112.930 3357.490 114.110 3358.670 ;
        RECT 112.930 3179.090 114.110 3180.270 ;
        RECT 112.930 3177.490 114.110 3178.670 ;
        RECT 112.930 2999.090 114.110 3000.270 ;
        RECT 112.930 2997.490 114.110 2998.670 ;
        RECT 112.930 2819.090 114.110 2820.270 ;
        RECT 112.930 2817.490 114.110 2818.670 ;
        RECT 112.930 2639.090 114.110 2640.270 ;
        RECT 112.930 2637.490 114.110 2638.670 ;
        RECT 112.930 2459.090 114.110 2460.270 ;
        RECT 112.930 2457.490 114.110 2458.670 ;
        RECT 112.930 2279.090 114.110 2280.270 ;
        RECT 112.930 2277.490 114.110 2278.670 ;
        RECT 112.930 2099.090 114.110 2100.270 ;
        RECT 112.930 2097.490 114.110 2098.670 ;
        RECT 112.930 1919.090 114.110 1920.270 ;
        RECT 112.930 1917.490 114.110 1918.670 ;
        RECT 112.930 1739.090 114.110 1740.270 ;
        RECT 112.930 1737.490 114.110 1738.670 ;
        RECT 112.930 1559.090 114.110 1560.270 ;
        RECT 112.930 1557.490 114.110 1558.670 ;
        RECT 112.930 1379.090 114.110 1380.270 ;
        RECT 112.930 1377.490 114.110 1378.670 ;
        RECT 112.930 1199.090 114.110 1200.270 ;
        RECT 112.930 1197.490 114.110 1198.670 ;
        RECT 112.930 1019.090 114.110 1020.270 ;
        RECT 112.930 1017.490 114.110 1018.670 ;
        RECT 112.930 839.090 114.110 840.270 ;
        RECT 112.930 837.490 114.110 838.670 ;
        RECT 112.930 659.090 114.110 660.270 ;
        RECT 112.930 657.490 114.110 658.670 ;
        RECT 112.930 479.090 114.110 480.270 ;
        RECT 112.930 477.490 114.110 478.670 ;
        RECT 112.930 299.090 114.110 300.270 ;
        RECT 112.930 297.490 114.110 298.670 ;
        RECT 112.930 119.090 114.110 120.270 ;
        RECT 112.930 117.490 114.110 118.670 ;
        RECT 112.930 -16.710 114.110 -15.530 ;
        RECT 112.930 -18.310 114.110 -17.130 ;
        RECT 292.930 3536.810 294.110 3537.990 ;
        RECT 292.930 3535.210 294.110 3536.390 ;
        RECT 292.930 3359.090 294.110 3360.270 ;
        RECT 292.930 3357.490 294.110 3358.670 ;
        RECT 292.930 3179.090 294.110 3180.270 ;
        RECT 292.930 3177.490 294.110 3178.670 ;
        RECT 292.930 2999.090 294.110 3000.270 ;
        RECT 292.930 2997.490 294.110 2998.670 ;
        RECT 292.930 2819.090 294.110 2820.270 ;
        RECT 292.930 2817.490 294.110 2818.670 ;
        RECT 292.930 2639.090 294.110 2640.270 ;
        RECT 292.930 2637.490 294.110 2638.670 ;
        RECT 292.930 2459.090 294.110 2460.270 ;
        RECT 292.930 2457.490 294.110 2458.670 ;
        RECT 292.930 2279.090 294.110 2280.270 ;
        RECT 292.930 2277.490 294.110 2278.670 ;
        RECT 292.930 2099.090 294.110 2100.270 ;
        RECT 292.930 2097.490 294.110 2098.670 ;
        RECT 292.930 1919.090 294.110 1920.270 ;
        RECT 292.930 1917.490 294.110 1918.670 ;
        RECT 292.930 1739.090 294.110 1740.270 ;
        RECT 292.930 1737.490 294.110 1738.670 ;
        RECT 292.930 1559.090 294.110 1560.270 ;
        RECT 292.930 1557.490 294.110 1558.670 ;
        RECT 292.930 1379.090 294.110 1380.270 ;
        RECT 292.930 1377.490 294.110 1378.670 ;
        RECT 292.930 1199.090 294.110 1200.270 ;
        RECT 292.930 1197.490 294.110 1198.670 ;
        RECT 292.930 1019.090 294.110 1020.270 ;
        RECT 292.930 1017.490 294.110 1018.670 ;
        RECT 292.930 839.090 294.110 840.270 ;
        RECT 292.930 837.490 294.110 838.670 ;
        RECT 292.930 659.090 294.110 660.270 ;
        RECT 292.930 657.490 294.110 658.670 ;
        RECT 292.930 479.090 294.110 480.270 ;
        RECT 292.930 477.490 294.110 478.670 ;
        RECT 292.930 299.090 294.110 300.270 ;
        RECT 292.930 297.490 294.110 298.670 ;
        RECT 292.930 119.090 294.110 120.270 ;
        RECT 292.930 117.490 294.110 118.670 ;
        RECT 292.930 -16.710 294.110 -15.530 ;
        RECT 292.930 -18.310 294.110 -17.130 ;
        RECT 472.930 3536.810 474.110 3537.990 ;
        RECT 472.930 3535.210 474.110 3536.390 ;
        RECT 472.930 3359.090 474.110 3360.270 ;
        RECT 472.930 3357.490 474.110 3358.670 ;
        RECT 472.930 3179.090 474.110 3180.270 ;
        RECT 472.930 3177.490 474.110 3178.670 ;
        RECT 472.930 2999.090 474.110 3000.270 ;
        RECT 472.930 2997.490 474.110 2998.670 ;
        RECT 472.930 2819.090 474.110 2820.270 ;
        RECT 472.930 2817.490 474.110 2818.670 ;
        RECT 472.930 2639.090 474.110 2640.270 ;
        RECT 472.930 2637.490 474.110 2638.670 ;
        RECT 472.930 2459.090 474.110 2460.270 ;
        RECT 472.930 2457.490 474.110 2458.670 ;
        RECT 472.930 2279.090 474.110 2280.270 ;
        RECT 472.930 2277.490 474.110 2278.670 ;
        RECT 472.930 2099.090 474.110 2100.270 ;
        RECT 472.930 2097.490 474.110 2098.670 ;
        RECT 472.930 1919.090 474.110 1920.270 ;
        RECT 472.930 1917.490 474.110 1918.670 ;
        RECT 472.930 1739.090 474.110 1740.270 ;
        RECT 472.930 1737.490 474.110 1738.670 ;
        RECT 472.930 1559.090 474.110 1560.270 ;
        RECT 472.930 1557.490 474.110 1558.670 ;
        RECT 472.930 1379.090 474.110 1380.270 ;
        RECT 472.930 1377.490 474.110 1378.670 ;
        RECT 472.930 1199.090 474.110 1200.270 ;
        RECT 472.930 1197.490 474.110 1198.670 ;
        RECT 472.930 1019.090 474.110 1020.270 ;
        RECT 472.930 1017.490 474.110 1018.670 ;
        RECT 472.930 839.090 474.110 840.270 ;
        RECT 472.930 837.490 474.110 838.670 ;
        RECT 472.930 659.090 474.110 660.270 ;
        RECT 472.930 657.490 474.110 658.670 ;
        RECT 472.930 479.090 474.110 480.270 ;
        RECT 472.930 477.490 474.110 478.670 ;
        RECT 472.930 299.090 474.110 300.270 ;
        RECT 472.930 297.490 474.110 298.670 ;
        RECT 472.930 119.090 474.110 120.270 ;
        RECT 472.930 117.490 474.110 118.670 ;
        RECT 472.930 -16.710 474.110 -15.530 ;
        RECT 472.930 -18.310 474.110 -17.130 ;
        RECT 652.930 3536.810 654.110 3537.990 ;
        RECT 652.930 3535.210 654.110 3536.390 ;
        RECT 652.930 3359.090 654.110 3360.270 ;
        RECT 652.930 3357.490 654.110 3358.670 ;
        RECT 652.930 3179.090 654.110 3180.270 ;
        RECT 652.930 3177.490 654.110 3178.670 ;
        RECT 652.930 2999.090 654.110 3000.270 ;
        RECT 652.930 2997.490 654.110 2998.670 ;
        RECT 652.930 2819.090 654.110 2820.270 ;
        RECT 652.930 2817.490 654.110 2818.670 ;
        RECT 652.930 2639.090 654.110 2640.270 ;
        RECT 652.930 2637.490 654.110 2638.670 ;
        RECT 652.930 2459.090 654.110 2460.270 ;
        RECT 652.930 2457.490 654.110 2458.670 ;
        RECT 652.930 2279.090 654.110 2280.270 ;
        RECT 652.930 2277.490 654.110 2278.670 ;
        RECT 652.930 2099.090 654.110 2100.270 ;
        RECT 652.930 2097.490 654.110 2098.670 ;
        RECT 652.930 1919.090 654.110 1920.270 ;
        RECT 652.930 1917.490 654.110 1918.670 ;
        RECT 652.930 1739.090 654.110 1740.270 ;
        RECT 652.930 1737.490 654.110 1738.670 ;
        RECT 652.930 1559.090 654.110 1560.270 ;
        RECT 652.930 1557.490 654.110 1558.670 ;
        RECT 652.930 1379.090 654.110 1380.270 ;
        RECT 652.930 1377.490 654.110 1378.670 ;
        RECT 652.930 1199.090 654.110 1200.270 ;
        RECT 652.930 1197.490 654.110 1198.670 ;
        RECT 652.930 1019.090 654.110 1020.270 ;
        RECT 652.930 1017.490 654.110 1018.670 ;
        RECT 652.930 839.090 654.110 840.270 ;
        RECT 652.930 837.490 654.110 838.670 ;
        RECT 652.930 659.090 654.110 660.270 ;
        RECT 652.930 657.490 654.110 658.670 ;
        RECT 652.930 479.090 654.110 480.270 ;
        RECT 652.930 477.490 654.110 478.670 ;
        RECT 652.930 299.090 654.110 300.270 ;
        RECT 652.930 297.490 654.110 298.670 ;
        RECT 652.930 119.090 654.110 120.270 ;
        RECT 652.930 117.490 654.110 118.670 ;
        RECT 652.930 -16.710 654.110 -15.530 ;
        RECT 652.930 -18.310 654.110 -17.130 ;
        RECT 832.930 3536.810 834.110 3537.990 ;
        RECT 832.930 3535.210 834.110 3536.390 ;
        RECT 832.930 3359.090 834.110 3360.270 ;
        RECT 832.930 3357.490 834.110 3358.670 ;
        RECT 832.930 3179.090 834.110 3180.270 ;
        RECT 832.930 3177.490 834.110 3178.670 ;
        RECT 832.930 2999.090 834.110 3000.270 ;
        RECT 832.930 2997.490 834.110 2998.670 ;
        RECT 832.930 2819.090 834.110 2820.270 ;
        RECT 832.930 2817.490 834.110 2818.670 ;
        RECT 832.930 2639.090 834.110 2640.270 ;
        RECT 832.930 2637.490 834.110 2638.670 ;
        RECT 832.930 2459.090 834.110 2460.270 ;
        RECT 832.930 2457.490 834.110 2458.670 ;
        RECT 832.930 2279.090 834.110 2280.270 ;
        RECT 832.930 2277.490 834.110 2278.670 ;
        RECT 832.930 2099.090 834.110 2100.270 ;
        RECT 832.930 2097.490 834.110 2098.670 ;
        RECT 832.930 1919.090 834.110 1920.270 ;
        RECT 832.930 1917.490 834.110 1918.670 ;
        RECT 832.930 1739.090 834.110 1740.270 ;
        RECT 832.930 1737.490 834.110 1738.670 ;
        RECT 832.930 1559.090 834.110 1560.270 ;
        RECT 832.930 1557.490 834.110 1558.670 ;
        RECT 832.930 1379.090 834.110 1380.270 ;
        RECT 832.930 1377.490 834.110 1378.670 ;
        RECT 832.930 1199.090 834.110 1200.270 ;
        RECT 832.930 1197.490 834.110 1198.670 ;
        RECT 832.930 1019.090 834.110 1020.270 ;
        RECT 832.930 1017.490 834.110 1018.670 ;
        RECT 832.930 839.090 834.110 840.270 ;
        RECT 832.930 837.490 834.110 838.670 ;
        RECT 832.930 659.090 834.110 660.270 ;
        RECT 832.930 657.490 834.110 658.670 ;
        RECT 832.930 479.090 834.110 480.270 ;
        RECT 832.930 477.490 834.110 478.670 ;
        RECT 832.930 299.090 834.110 300.270 ;
        RECT 832.930 297.490 834.110 298.670 ;
        RECT 832.930 119.090 834.110 120.270 ;
        RECT 832.930 117.490 834.110 118.670 ;
        RECT 832.930 -16.710 834.110 -15.530 ;
        RECT 832.930 -18.310 834.110 -17.130 ;
        RECT 1012.930 3536.810 1014.110 3537.990 ;
        RECT 1012.930 3535.210 1014.110 3536.390 ;
        RECT 1012.930 3359.090 1014.110 3360.270 ;
        RECT 1012.930 3357.490 1014.110 3358.670 ;
        RECT 1012.930 3179.090 1014.110 3180.270 ;
        RECT 1012.930 3177.490 1014.110 3178.670 ;
        RECT 1012.930 2999.090 1014.110 3000.270 ;
        RECT 1012.930 2997.490 1014.110 2998.670 ;
        RECT 1012.930 2819.090 1014.110 2820.270 ;
        RECT 1012.930 2817.490 1014.110 2818.670 ;
        RECT 1012.930 2639.090 1014.110 2640.270 ;
        RECT 1012.930 2637.490 1014.110 2638.670 ;
        RECT 1012.930 2459.090 1014.110 2460.270 ;
        RECT 1012.930 2457.490 1014.110 2458.670 ;
        RECT 1012.930 2279.090 1014.110 2280.270 ;
        RECT 1012.930 2277.490 1014.110 2278.670 ;
        RECT 1012.930 2099.090 1014.110 2100.270 ;
        RECT 1012.930 2097.490 1014.110 2098.670 ;
        RECT 1012.930 1919.090 1014.110 1920.270 ;
        RECT 1012.930 1917.490 1014.110 1918.670 ;
        RECT 1012.930 1739.090 1014.110 1740.270 ;
        RECT 1012.930 1737.490 1014.110 1738.670 ;
        RECT 1012.930 1559.090 1014.110 1560.270 ;
        RECT 1012.930 1557.490 1014.110 1558.670 ;
        RECT 1012.930 1379.090 1014.110 1380.270 ;
        RECT 1012.930 1377.490 1014.110 1378.670 ;
        RECT 1012.930 1199.090 1014.110 1200.270 ;
        RECT 1012.930 1197.490 1014.110 1198.670 ;
        RECT 1012.930 1019.090 1014.110 1020.270 ;
        RECT 1012.930 1017.490 1014.110 1018.670 ;
        RECT 1012.930 839.090 1014.110 840.270 ;
        RECT 1012.930 837.490 1014.110 838.670 ;
        RECT 1012.930 659.090 1014.110 660.270 ;
        RECT 1012.930 657.490 1014.110 658.670 ;
        RECT 1012.930 479.090 1014.110 480.270 ;
        RECT 1012.930 477.490 1014.110 478.670 ;
        RECT 1012.930 299.090 1014.110 300.270 ;
        RECT 1012.930 297.490 1014.110 298.670 ;
        RECT 1012.930 119.090 1014.110 120.270 ;
        RECT 1012.930 117.490 1014.110 118.670 ;
        RECT 1012.930 -16.710 1014.110 -15.530 ;
        RECT 1012.930 -18.310 1014.110 -17.130 ;
        RECT 1192.930 3536.810 1194.110 3537.990 ;
        RECT 1192.930 3535.210 1194.110 3536.390 ;
        RECT 1192.930 3359.090 1194.110 3360.270 ;
        RECT 1192.930 3357.490 1194.110 3358.670 ;
        RECT 1192.930 3179.090 1194.110 3180.270 ;
        RECT 1192.930 3177.490 1194.110 3178.670 ;
        RECT 1192.930 2999.090 1194.110 3000.270 ;
        RECT 1192.930 2997.490 1194.110 2998.670 ;
        RECT 1192.930 2819.090 1194.110 2820.270 ;
        RECT 1192.930 2817.490 1194.110 2818.670 ;
        RECT 1192.930 2639.090 1194.110 2640.270 ;
        RECT 1192.930 2637.490 1194.110 2638.670 ;
        RECT 1192.930 2459.090 1194.110 2460.270 ;
        RECT 1192.930 2457.490 1194.110 2458.670 ;
        RECT 1192.930 2279.090 1194.110 2280.270 ;
        RECT 1192.930 2277.490 1194.110 2278.670 ;
        RECT 1192.930 2099.090 1194.110 2100.270 ;
        RECT 1192.930 2097.490 1194.110 2098.670 ;
        RECT 1192.930 1919.090 1194.110 1920.270 ;
        RECT 1192.930 1917.490 1194.110 1918.670 ;
        RECT 1192.930 1739.090 1194.110 1740.270 ;
        RECT 1192.930 1737.490 1194.110 1738.670 ;
        RECT 1192.930 1559.090 1194.110 1560.270 ;
        RECT 1192.930 1557.490 1194.110 1558.670 ;
        RECT 1192.930 1379.090 1194.110 1380.270 ;
        RECT 1192.930 1377.490 1194.110 1378.670 ;
        RECT 1192.930 1199.090 1194.110 1200.270 ;
        RECT 1192.930 1197.490 1194.110 1198.670 ;
        RECT 1192.930 1019.090 1194.110 1020.270 ;
        RECT 1192.930 1017.490 1194.110 1018.670 ;
        RECT 1192.930 839.090 1194.110 840.270 ;
        RECT 1192.930 837.490 1194.110 838.670 ;
        RECT 1192.930 659.090 1194.110 660.270 ;
        RECT 1192.930 657.490 1194.110 658.670 ;
        RECT 1192.930 479.090 1194.110 480.270 ;
        RECT 1192.930 477.490 1194.110 478.670 ;
        RECT 1192.930 299.090 1194.110 300.270 ;
        RECT 1192.930 297.490 1194.110 298.670 ;
        RECT 1192.930 119.090 1194.110 120.270 ;
        RECT 1192.930 117.490 1194.110 118.670 ;
        RECT 1192.930 -16.710 1194.110 -15.530 ;
        RECT 1192.930 -18.310 1194.110 -17.130 ;
        RECT 1372.930 3536.810 1374.110 3537.990 ;
        RECT 1372.930 3535.210 1374.110 3536.390 ;
        RECT 1372.930 3359.090 1374.110 3360.270 ;
        RECT 1372.930 3357.490 1374.110 3358.670 ;
        RECT 1372.930 3179.090 1374.110 3180.270 ;
        RECT 1372.930 3177.490 1374.110 3178.670 ;
        RECT 1372.930 2999.090 1374.110 3000.270 ;
        RECT 1372.930 2997.490 1374.110 2998.670 ;
        RECT 1372.930 2819.090 1374.110 2820.270 ;
        RECT 1372.930 2817.490 1374.110 2818.670 ;
        RECT 1372.930 2639.090 1374.110 2640.270 ;
        RECT 1372.930 2637.490 1374.110 2638.670 ;
        RECT 1372.930 2459.090 1374.110 2460.270 ;
        RECT 1372.930 2457.490 1374.110 2458.670 ;
        RECT 1372.930 2279.090 1374.110 2280.270 ;
        RECT 1372.930 2277.490 1374.110 2278.670 ;
        RECT 1372.930 2099.090 1374.110 2100.270 ;
        RECT 1372.930 2097.490 1374.110 2098.670 ;
        RECT 1372.930 1919.090 1374.110 1920.270 ;
        RECT 1372.930 1917.490 1374.110 1918.670 ;
        RECT 1372.930 1739.090 1374.110 1740.270 ;
        RECT 1372.930 1737.490 1374.110 1738.670 ;
        RECT 1372.930 1559.090 1374.110 1560.270 ;
        RECT 1372.930 1557.490 1374.110 1558.670 ;
        RECT 1372.930 1379.090 1374.110 1380.270 ;
        RECT 1372.930 1377.490 1374.110 1378.670 ;
        RECT 1372.930 1199.090 1374.110 1200.270 ;
        RECT 1372.930 1197.490 1374.110 1198.670 ;
        RECT 1372.930 1019.090 1374.110 1020.270 ;
        RECT 1372.930 1017.490 1374.110 1018.670 ;
        RECT 1372.930 839.090 1374.110 840.270 ;
        RECT 1372.930 837.490 1374.110 838.670 ;
        RECT 1372.930 659.090 1374.110 660.270 ;
        RECT 1372.930 657.490 1374.110 658.670 ;
        RECT 1372.930 479.090 1374.110 480.270 ;
        RECT 1372.930 477.490 1374.110 478.670 ;
        RECT 1372.930 299.090 1374.110 300.270 ;
        RECT 1372.930 297.490 1374.110 298.670 ;
        RECT 1372.930 119.090 1374.110 120.270 ;
        RECT 1372.930 117.490 1374.110 118.670 ;
        RECT 1372.930 -16.710 1374.110 -15.530 ;
        RECT 1372.930 -18.310 1374.110 -17.130 ;
        RECT 1552.930 3536.810 1554.110 3537.990 ;
        RECT 1552.930 3535.210 1554.110 3536.390 ;
        RECT 1552.930 3359.090 1554.110 3360.270 ;
        RECT 1552.930 3357.490 1554.110 3358.670 ;
        RECT 1552.930 3179.090 1554.110 3180.270 ;
        RECT 1552.930 3177.490 1554.110 3178.670 ;
        RECT 1552.930 2999.090 1554.110 3000.270 ;
        RECT 1552.930 2997.490 1554.110 2998.670 ;
        RECT 1552.930 2819.090 1554.110 2820.270 ;
        RECT 1552.930 2817.490 1554.110 2818.670 ;
        RECT 1552.930 2639.090 1554.110 2640.270 ;
        RECT 1552.930 2637.490 1554.110 2638.670 ;
        RECT 1552.930 2459.090 1554.110 2460.270 ;
        RECT 1552.930 2457.490 1554.110 2458.670 ;
        RECT 1552.930 2279.090 1554.110 2280.270 ;
        RECT 1552.930 2277.490 1554.110 2278.670 ;
        RECT 1552.930 2099.090 1554.110 2100.270 ;
        RECT 1552.930 2097.490 1554.110 2098.670 ;
        RECT 1552.930 1919.090 1554.110 1920.270 ;
        RECT 1552.930 1917.490 1554.110 1918.670 ;
        RECT 1552.930 1739.090 1554.110 1740.270 ;
        RECT 1552.930 1737.490 1554.110 1738.670 ;
        RECT 1552.930 1559.090 1554.110 1560.270 ;
        RECT 1552.930 1557.490 1554.110 1558.670 ;
        RECT 1552.930 1379.090 1554.110 1380.270 ;
        RECT 1552.930 1377.490 1554.110 1378.670 ;
        RECT 1552.930 1199.090 1554.110 1200.270 ;
        RECT 1552.930 1197.490 1554.110 1198.670 ;
        RECT 1552.930 1019.090 1554.110 1020.270 ;
        RECT 1552.930 1017.490 1554.110 1018.670 ;
        RECT 1552.930 839.090 1554.110 840.270 ;
        RECT 1552.930 837.490 1554.110 838.670 ;
        RECT 1552.930 659.090 1554.110 660.270 ;
        RECT 1552.930 657.490 1554.110 658.670 ;
        RECT 1552.930 479.090 1554.110 480.270 ;
        RECT 1552.930 477.490 1554.110 478.670 ;
        RECT 1552.930 299.090 1554.110 300.270 ;
        RECT 1552.930 297.490 1554.110 298.670 ;
        RECT 1552.930 119.090 1554.110 120.270 ;
        RECT 1552.930 117.490 1554.110 118.670 ;
        RECT 1552.930 -16.710 1554.110 -15.530 ;
        RECT 1552.930 -18.310 1554.110 -17.130 ;
        RECT 1732.930 3536.810 1734.110 3537.990 ;
        RECT 1732.930 3535.210 1734.110 3536.390 ;
        RECT 1732.930 3359.090 1734.110 3360.270 ;
        RECT 1732.930 3357.490 1734.110 3358.670 ;
        RECT 1732.930 3179.090 1734.110 3180.270 ;
        RECT 1732.930 3177.490 1734.110 3178.670 ;
        RECT 1732.930 2999.090 1734.110 3000.270 ;
        RECT 1732.930 2997.490 1734.110 2998.670 ;
        RECT 1732.930 2819.090 1734.110 2820.270 ;
        RECT 1732.930 2817.490 1734.110 2818.670 ;
        RECT 1732.930 2639.090 1734.110 2640.270 ;
        RECT 1732.930 2637.490 1734.110 2638.670 ;
        RECT 1732.930 2459.090 1734.110 2460.270 ;
        RECT 1732.930 2457.490 1734.110 2458.670 ;
        RECT 1732.930 2279.090 1734.110 2280.270 ;
        RECT 1732.930 2277.490 1734.110 2278.670 ;
        RECT 1732.930 2099.090 1734.110 2100.270 ;
        RECT 1732.930 2097.490 1734.110 2098.670 ;
        RECT 1732.930 1919.090 1734.110 1920.270 ;
        RECT 1732.930 1917.490 1734.110 1918.670 ;
        RECT 1732.930 1739.090 1734.110 1740.270 ;
        RECT 1732.930 1737.490 1734.110 1738.670 ;
        RECT 1732.930 1559.090 1734.110 1560.270 ;
        RECT 1732.930 1557.490 1734.110 1558.670 ;
        RECT 1732.930 1379.090 1734.110 1380.270 ;
        RECT 1732.930 1377.490 1734.110 1378.670 ;
        RECT 1732.930 1199.090 1734.110 1200.270 ;
        RECT 1732.930 1197.490 1734.110 1198.670 ;
        RECT 1732.930 1019.090 1734.110 1020.270 ;
        RECT 1732.930 1017.490 1734.110 1018.670 ;
        RECT 1732.930 839.090 1734.110 840.270 ;
        RECT 1732.930 837.490 1734.110 838.670 ;
        RECT 1732.930 659.090 1734.110 660.270 ;
        RECT 1732.930 657.490 1734.110 658.670 ;
        RECT 1732.930 479.090 1734.110 480.270 ;
        RECT 1732.930 477.490 1734.110 478.670 ;
        RECT 1732.930 299.090 1734.110 300.270 ;
        RECT 1732.930 297.490 1734.110 298.670 ;
        RECT 1732.930 119.090 1734.110 120.270 ;
        RECT 1732.930 117.490 1734.110 118.670 ;
        RECT 1732.930 -16.710 1734.110 -15.530 ;
        RECT 1732.930 -18.310 1734.110 -17.130 ;
        RECT 1912.930 3536.810 1914.110 3537.990 ;
        RECT 1912.930 3535.210 1914.110 3536.390 ;
        RECT 1912.930 3359.090 1914.110 3360.270 ;
        RECT 1912.930 3357.490 1914.110 3358.670 ;
        RECT 1912.930 3179.090 1914.110 3180.270 ;
        RECT 1912.930 3177.490 1914.110 3178.670 ;
        RECT 1912.930 2999.090 1914.110 3000.270 ;
        RECT 1912.930 2997.490 1914.110 2998.670 ;
        RECT 1912.930 2819.090 1914.110 2820.270 ;
        RECT 1912.930 2817.490 1914.110 2818.670 ;
        RECT 1912.930 2639.090 1914.110 2640.270 ;
        RECT 1912.930 2637.490 1914.110 2638.670 ;
        RECT 1912.930 2459.090 1914.110 2460.270 ;
        RECT 1912.930 2457.490 1914.110 2458.670 ;
        RECT 1912.930 2279.090 1914.110 2280.270 ;
        RECT 1912.930 2277.490 1914.110 2278.670 ;
        RECT 1912.930 2099.090 1914.110 2100.270 ;
        RECT 1912.930 2097.490 1914.110 2098.670 ;
        RECT 1912.930 1919.090 1914.110 1920.270 ;
        RECT 1912.930 1917.490 1914.110 1918.670 ;
        RECT 1912.930 1739.090 1914.110 1740.270 ;
        RECT 1912.930 1737.490 1914.110 1738.670 ;
        RECT 1912.930 1559.090 1914.110 1560.270 ;
        RECT 1912.930 1557.490 1914.110 1558.670 ;
        RECT 1912.930 1379.090 1914.110 1380.270 ;
        RECT 1912.930 1377.490 1914.110 1378.670 ;
        RECT 1912.930 1199.090 1914.110 1200.270 ;
        RECT 1912.930 1197.490 1914.110 1198.670 ;
        RECT 1912.930 1019.090 1914.110 1020.270 ;
        RECT 1912.930 1017.490 1914.110 1018.670 ;
        RECT 1912.930 839.090 1914.110 840.270 ;
        RECT 1912.930 837.490 1914.110 838.670 ;
        RECT 1912.930 659.090 1914.110 660.270 ;
        RECT 1912.930 657.490 1914.110 658.670 ;
        RECT 1912.930 479.090 1914.110 480.270 ;
        RECT 1912.930 477.490 1914.110 478.670 ;
        RECT 1912.930 299.090 1914.110 300.270 ;
        RECT 1912.930 297.490 1914.110 298.670 ;
        RECT 1912.930 119.090 1914.110 120.270 ;
        RECT 1912.930 117.490 1914.110 118.670 ;
        RECT 1912.930 -16.710 1914.110 -15.530 ;
        RECT 1912.930 -18.310 1914.110 -17.130 ;
        RECT 2092.930 3536.810 2094.110 3537.990 ;
        RECT 2092.930 3535.210 2094.110 3536.390 ;
        RECT 2092.930 3359.090 2094.110 3360.270 ;
        RECT 2092.930 3357.490 2094.110 3358.670 ;
        RECT 2092.930 3179.090 2094.110 3180.270 ;
        RECT 2092.930 3177.490 2094.110 3178.670 ;
        RECT 2092.930 2999.090 2094.110 3000.270 ;
        RECT 2092.930 2997.490 2094.110 2998.670 ;
        RECT 2092.930 2819.090 2094.110 2820.270 ;
        RECT 2092.930 2817.490 2094.110 2818.670 ;
        RECT 2092.930 2639.090 2094.110 2640.270 ;
        RECT 2092.930 2637.490 2094.110 2638.670 ;
        RECT 2092.930 2459.090 2094.110 2460.270 ;
        RECT 2092.930 2457.490 2094.110 2458.670 ;
        RECT 2092.930 2279.090 2094.110 2280.270 ;
        RECT 2092.930 2277.490 2094.110 2278.670 ;
        RECT 2092.930 2099.090 2094.110 2100.270 ;
        RECT 2092.930 2097.490 2094.110 2098.670 ;
        RECT 2092.930 1919.090 2094.110 1920.270 ;
        RECT 2092.930 1917.490 2094.110 1918.670 ;
        RECT 2092.930 1739.090 2094.110 1740.270 ;
        RECT 2092.930 1737.490 2094.110 1738.670 ;
        RECT 2092.930 1559.090 2094.110 1560.270 ;
        RECT 2092.930 1557.490 2094.110 1558.670 ;
        RECT 2092.930 1379.090 2094.110 1380.270 ;
        RECT 2092.930 1377.490 2094.110 1378.670 ;
        RECT 2092.930 1199.090 2094.110 1200.270 ;
        RECT 2092.930 1197.490 2094.110 1198.670 ;
        RECT 2092.930 1019.090 2094.110 1020.270 ;
        RECT 2092.930 1017.490 2094.110 1018.670 ;
        RECT 2092.930 839.090 2094.110 840.270 ;
        RECT 2092.930 837.490 2094.110 838.670 ;
        RECT 2092.930 659.090 2094.110 660.270 ;
        RECT 2092.930 657.490 2094.110 658.670 ;
        RECT 2092.930 479.090 2094.110 480.270 ;
        RECT 2092.930 477.490 2094.110 478.670 ;
        RECT 2092.930 299.090 2094.110 300.270 ;
        RECT 2092.930 297.490 2094.110 298.670 ;
        RECT 2092.930 119.090 2094.110 120.270 ;
        RECT 2092.930 117.490 2094.110 118.670 ;
        RECT 2092.930 -16.710 2094.110 -15.530 ;
        RECT 2092.930 -18.310 2094.110 -17.130 ;
        RECT 2272.930 3536.810 2274.110 3537.990 ;
        RECT 2272.930 3535.210 2274.110 3536.390 ;
        RECT 2272.930 3359.090 2274.110 3360.270 ;
        RECT 2272.930 3357.490 2274.110 3358.670 ;
        RECT 2272.930 3179.090 2274.110 3180.270 ;
        RECT 2272.930 3177.490 2274.110 3178.670 ;
        RECT 2272.930 2999.090 2274.110 3000.270 ;
        RECT 2272.930 2997.490 2274.110 2998.670 ;
        RECT 2272.930 2819.090 2274.110 2820.270 ;
        RECT 2272.930 2817.490 2274.110 2818.670 ;
        RECT 2272.930 2639.090 2274.110 2640.270 ;
        RECT 2272.930 2637.490 2274.110 2638.670 ;
        RECT 2272.930 2459.090 2274.110 2460.270 ;
        RECT 2272.930 2457.490 2274.110 2458.670 ;
        RECT 2272.930 2279.090 2274.110 2280.270 ;
        RECT 2272.930 2277.490 2274.110 2278.670 ;
        RECT 2272.930 2099.090 2274.110 2100.270 ;
        RECT 2272.930 2097.490 2274.110 2098.670 ;
        RECT 2272.930 1919.090 2274.110 1920.270 ;
        RECT 2272.930 1917.490 2274.110 1918.670 ;
        RECT 2272.930 1739.090 2274.110 1740.270 ;
        RECT 2272.930 1737.490 2274.110 1738.670 ;
        RECT 2272.930 1559.090 2274.110 1560.270 ;
        RECT 2272.930 1557.490 2274.110 1558.670 ;
        RECT 2272.930 1379.090 2274.110 1380.270 ;
        RECT 2272.930 1377.490 2274.110 1378.670 ;
        RECT 2272.930 1199.090 2274.110 1200.270 ;
        RECT 2272.930 1197.490 2274.110 1198.670 ;
        RECT 2272.930 1019.090 2274.110 1020.270 ;
        RECT 2272.930 1017.490 2274.110 1018.670 ;
        RECT 2272.930 839.090 2274.110 840.270 ;
        RECT 2272.930 837.490 2274.110 838.670 ;
        RECT 2272.930 659.090 2274.110 660.270 ;
        RECT 2272.930 657.490 2274.110 658.670 ;
        RECT 2272.930 479.090 2274.110 480.270 ;
        RECT 2272.930 477.490 2274.110 478.670 ;
        RECT 2272.930 299.090 2274.110 300.270 ;
        RECT 2272.930 297.490 2274.110 298.670 ;
        RECT 2272.930 119.090 2274.110 120.270 ;
        RECT 2272.930 117.490 2274.110 118.670 ;
        RECT 2272.930 -16.710 2274.110 -15.530 ;
        RECT 2272.930 -18.310 2274.110 -17.130 ;
        RECT 2452.930 3536.810 2454.110 3537.990 ;
        RECT 2452.930 3535.210 2454.110 3536.390 ;
        RECT 2452.930 3359.090 2454.110 3360.270 ;
        RECT 2452.930 3357.490 2454.110 3358.670 ;
        RECT 2452.930 3179.090 2454.110 3180.270 ;
        RECT 2452.930 3177.490 2454.110 3178.670 ;
        RECT 2452.930 2999.090 2454.110 3000.270 ;
        RECT 2452.930 2997.490 2454.110 2998.670 ;
        RECT 2452.930 2819.090 2454.110 2820.270 ;
        RECT 2452.930 2817.490 2454.110 2818.670 ;
        RECT 2452.930 2639.090 2454.110 2640.270 ;
        RECT 2452.930 2637.490 2454.110 2638.670 ;
        RECT 2452.930 2459.090 2454.110 2460.270 ;
        RECT 2452.930 2457.490 2454.110 2458.670 ;
        RECT 2452.930 2279.090 2454.110 2280.270 ;
        RECT 2452.930 2277.490 2454.110 2278.670 ;
        RECT 2452.930 2099.090 2454.110 2100.270 ;
        RECT 2452.930 2097.490 2454.110 2098.670 ;
        RECT 2452.930 1919.090 2454.110 1920.270 ;
        RECT 2452.930 1917.490 2454.110 1918.670 ;
        RECT 2452.930 1739.090 2454.110 1740.270 ;
        RECT 2452.930 1737.490 2454.110 1738.670 ;
        RECT 2452.930 1559.090 2454.110 1560.270 ;
        RECT 2452.930 1557.490 2454.110 1558.670 ;
        RECT 2452.930 1379.090 2454.110 1380.270 ;
        RECT 2452.930 1377.490 2454.110 1378.670 ;
        RECT 2452.930 1199.090 2454.110 1200.270 ;
        RECT 2452.930 1197.490 2454.110 1198.670 ;
        RECT 2452.930 1019.090 2454.110 1020.270 ;
        RECT 2452.930 1017.490 2454.110 1018.670 ;
        RECT 2452.930 839.090 2454.110 840.270 ;
        RECT 2452.930 837.490 2454.110 838.670 ;
        RECT 2452.930 659.090 2454.110 660.270 ;
        RECT 2452.930 657.490 2454.110 658.670 ;
        RECT 2452.930 479.090 2454.110 480.270 ;
        RECT 2452.930 477.490 2454.110 478.670 ;
        RECT 2452.930 299.090 2454.110 300.270 ;
        RECT 2452.930 297.490 2454.110 298.670 ;
        RECT 2452.930 119.090 2454.110 120.270 ;
        RECT 2452.930 117.490 2454.110 118.670 ;
        RECT 2452.930 -16.710 2454.110 -15.530 ;
        RECT 2452.930 -18.310 2454.110 -17.130 ;
        RECT 2632.930 3536.810 2634.110 3537.990 ;
        RECT 2632.930 3535.210 2634.110 3536.390 ;
        RECT 2632.930 3359.090 2634.110 3360.270 ;
        RECT 2632.930 3357.490 2634.110 3358.670 ;
        RECT 2632.930 3179.090 2634.110 3180.270 ;
        RECT 2632.930 3177.490 2634.110 3178.670 ;
        RECT 2632.930 2999.090 2634.110 3000.270 ;
        RECT 2632.930 2997.490 2634.110 2998.670 ;
        RECT 2632.930 2819.090 2634.110 2820.270 ;
        RECT 2632.930 2817.490 2634.110 2818.670 ;
        RECT 2632.930 2639.090 2634.110 2640.270 ;
        RECT 2632.930 2637.490 2634.110 2638.670 ;
        RECT 2632.930 2459.090 2634.110 2460.270 ;
        RECT 2632.930 2457.490 2634.110 2458.670 ;
        RECT 2632.930 2279.090 2634.110 2280.270 ;
        RECT 2632.930 2277.490 2634.110 2278.670 ;
        RECT 2632.930 2099.090 2634.110 2100.270 ;
        RECT 2632.930 2097.490 2634.110 2098.670 ;
        RECT 2632.930 1919.090 2634.110 1920.270 ;
        RECT 2632.930 1917.490 2634.110 1918.670 ;
        RECT 2632.930 1739.090 2634.110 1740.270 ;
        RECT 2632.930 1737.490 2634.110 1738.670 ;
        RECT 2632.930 1559.090 2634.110 1560.270 ;
        RECT 2632.930 1557.490 2634.110 1558.670 ;
        RECT 2632.930 1379.090 2634.110 1380.270 ;
        RECT 2632.930 1377.490 2634.110 1378.670 ;
        RECT 2632.930 1199.090 2634.110 1200.270 ;
        RECT 2632.930 1197.490 2634.110 1198.670 ;
        RECT 2632.930 1019.090 2634.110 1020.270 ;
        RECT 2632.930 1017.490 2634.110 1018.670 ;
        RECT 2632.930 839.090 2634.110 840.270 ;
        RECT 2632.930 837.490 2634.110 838.670 ;
        RECT 2632.930 659.090 2634.110 660.270 ;
        RECT 2632.930 657.490 2634.110 658.670 ;
        RECT 2632.930 479.090 2634.110 480.270 ;
        RECT 2632.930 477.490 2634.110 478.670 ;
        RECT 2632.930 299.090 2634.110 300.270 ;
        RECT 2632.930 297.490 2634.110 298.670 ;
        RECT 2632.930 119.090 2634.110 120.270 ;
        RECT 2632.930 117.490 2634.110 118.670 ;
        RECT 2632.930 -16.710 2634.110 -15.530 ;
        RECT 2632.930 -18.310 2634.110 -17.130 ;
        RECT 2812.930 3536.810 2814.110 3537.990 ;
        RECT 2812.930 3535.210 2814.110 3536.390 ;
        RECT 2812.930 3359.090 2814.110 3360.270 ;
        RECT 2812.930 3357.490 2814.110 3358.670 ;
        RECT 2812.930 3179.090 2814.110 3180.270 ;
        RECT 2812.930 3177.490 2814.110 3178.670 ;
        RECT 2812.930 2999.090 2814.110 3000.270 ;
        RECT 2812.930 2997.490 2814.110 2998.670 ;
        RECT 2812.930 2819.090 2814.110 2820.270 ;
        RECT 2812.930 2817.490 2814.110 2818.670 ;
        RECT 2812.930 2639.090 2814.110 2640.270 ;
        RECT 2812.930 2637.490 2814.110 2638.670 ;
        RECT 2812.930 2459.090 2814.110 2460.270 ;
        RECT 2812.930 2457.490 2814.110 2458.670 ;
        RECT 2812.930 2279.090 2814.110 2280.270 ;
        RECT 2812.930 2277.490 2814.110 2278.670 ;
        RECT 2812.930 2099.090 2814.110 2100.270 ;
        RECT 2812.930 2097.490 2814.110 2098.670 ;
        RECT 2812.930 1919.090 2814.110 1920.270 ;
        RECT 2812.930 1917.490 2814.110 1918.670 ;
        RECT 2812.930 1739.090 2814.110 1740.270 ;
        RECT 2812.930 1737.490 2814.110 1738.670 ;
        RECT 2812.930 1559.090 2814.110 1560.270 ;
        RECT 2812.930 1557.490 2814.110 1558.670 ;
        RECT 2812.930 1379.090 2814.110 1380.270 ;
        RECT 2812.930 1377.490 2814.110 1378.670 ;
        RECT 2812.930 1199.090 2814.110 1200.270 ;
        RECT 2812.930 1197.490 2814.110 1198.670 ;
        RECT 2812.930 1019.090 2814.110 1020.270 ;
        RECT 2812.930 1017.490 2814.110 1018.670 ;
        RECT 2812.930 839.090 2814.110 840.270 ;
        RECT 2812.930 837.490 2814.110 838.670 ;
        RECT 2812.930 659.090 2814.110 660.270 ;
        RECT 2812.930 657.490 2814.110 658.670 ;
        RECT 2812.930 479.090 2814.110 480.270 ;
        RECT 2812.930 477.490 2814.110 478.670 ;
        RECT 2812.930 299.090 2814.110 300.270 ;
        RECT 2812.930 297.490 2814.110 298.670 ;
        RECT 2812.930 119.090 2814.110 120.270 ;
        RECT 2812.930 117.490 2814.110 118.670 ;
        RECT 2812.930 -16.710 2814.110 -15.530 ;
        RECT 2812.930 -18.310 2814.110 -17.130 ;
        RECT 2941.310 3536.810 2942.490 3537.990 ;
        RECT 2941.310 3535.210 2942.490 3536.390 ;
        RECT 2941.310 3359.090 2942.490 3360.270 ;
        RECT 2941.310 3357.490 2942.490 3358.670 ;
        RECT 2941.310 3179.090 2942.490 3180.270 ;
        RECT 2941.310 3177.490 2942.490 3178.670 ;
        RECT 2941.310 2999.090 2942.490 3000.270 ;
        RECT 2941.310 2997.490 2942.490 2998.670 ;
        RECT 2941.310 2819.090 2942.490 2820.270 ;
        RECT 2941.310 2817.490 2942.490 2818.670 ;
        RECT 2941.310 2639.090 2942.490 2640.270 ;
        RECT 2941.310 2637.490 2942.490 2638.670 ;
        RECT 2941.310 2459.090 2942.490 2460.270 ;
        RECT 2941.310 2457.490 2942.490 2458.670 ;
        RECT 2941.310 2279.090 2942.490 2280.270 ;
        RECT 2941.310 2277.490 2942.490 2278.670 ;
        RECT 2941.310 2099.090 2942.490 2100.270 ;
        RECT 2941.310 2097.490 2942.490 2098.670 ;
        RECT 2941.310 1919.090 2942.490 1920.270 ;
        RECT 2941.310 1917.490 2942.490 1918.670 ;
        RECT 2941.310 1739.090 2942.490 1740.270 ;
        RECT 2941.310 1737.490 2942.490 1738.670 ;
        RECT 2941.310 1559.090 2942.490 1560.270 ;
        RECT 2941.310 1557.490 2942.490 1558.670 ;
        RECT 2941.310 1379.090 2942.490 1380.270 ;
        RECT 2941.310 1377.490 2942.490 1378.670 ;
        RECT 2941.310 1199.090 2942.490 1200.270 ;
        RECT 2941.310 1197.490 2942.490 1198.670 ;
        RECT 2941.310 1019.090 2942.490 1020.270 ;
        RECT 2941.310 1017.490 2942.490 1018.670 ;
        RECT 2941.310 839.090 2942.490 840.270 ;
        RECT 2941.310 837.490 2942.490 838.670 ;
        RECT 2941.310 659.090 2942.490 660.270 ;
        RECT 2941.310 657.490 2942.490 658.670 ;
        RECT 2941.310 479.090 2942.490 480.270 ;
        RECT 2941.310 477.490 2942.490 478.670 ;
        RECT 2941.310 299.090 2942.490 300.270 ;
        RECT 2941.310 297.490 2942.490 298.670 ;
        RECT 2941.310 119.090 2942.490 120.270 ;
        RECT 2941.310 117.490 2942.490 118.670 ;
        RECT 2941.310 -16.710 2942.490 -15.530 ;
        RECT 2941.310 -18.310 2942.490 -17.130 ;
      LAYER met5 ;
        RECT -23.780 3538.100 -20.780 3538.110 ;
        RECT 112.020 3538.100 115.020 3538.110 ;
        RECT 292.020 3538.100 295.020 3538.110 ;
        RECT 472.020 3538.100 475.020 3538.110 ;
        RECT 652.020 3538.100 655.020 3538.110 ;
        RECT 832.020 3538.100 835.020 3538.110 ;
        RECT 1012.020 3538.100 1015.020 3538.110 ;
        RECT 1192.020 3538.100 1195.020 3538.110 ;
        RECT 1372.020 3538.100 1375.020 3538.110 ;
        RECT 1552.020 3538.100 1555.020 3538.110 ;
        RECT 1732.020 3538.100 1735.020 3538.110 ;
        RECT 1912.020 3538.100 1915.020 3538.110 ;
        RECT 2092.020 3538.100 2095.020 3538.110 ;
        RECT 2272.020 3538.100 2275.020 3538.110 ;
        RECT 2452.020 3538.100 2455.020 3538.110 ;
        RECT 2632.020 3538.100 2635.020 3538.110 ;
        RECT 2812.020 3538.100 2815.020 3538.110 ;
        RECT 2940.400 3538.100 2943.400 3538.110 ;
        RECT -23.780 3535.100 2943.400 3538.100 ;
        RECT -23.780 3535.090 -20.780 3535.100 ;
        RECT 112.020 3535.090 115.020 3535.100 ;
        RECT 292.020 3535.090 295.020 3535.100 ;
        RECT 472.020 3535.090 475.020 3535.100 ;
        RECT 652.020 3535.090 655.020 3535.100 ;
        RECT 832.020 3535.090 835.020 3535.100 ;
        RECT 1012.020 3535.090 1015.020 3535.100 ;
        RECT 1192.020 3535.090 1195.020 3535.100 ;
        RECT 1372.020 3535.090 1375.020 3535.100 ;
        RECT 1552.020 3535.090 1555.020 3535.100 ;
        RECT 1732.020 3535.090 1735.020 3535.100 ;
        RECT 1912.020 3535.090 1915.020 3535.100 ;
        RECT 2092.020 3535.090 2095.020 3535.100 ;
        RECT 2272.020 3535.090 2275.020 3535.100 ;
        RECT 2452.020 3535.090 2455.020 3535.100 ;
        RECT 2632.020 3535.090 2635.020 3535.100 ;
        RECT 2812.020 3535.090 2815.020 3535.100 ;
        RECT 2940.400 3535.090 2943.400 3535.100 ;
        RECT -23.780 3360.380 -20.780 3360.390 ;
        RECT 112.020 3360.380 115.020 3360.390 ;
        RECT 292.020 3360.380 295.020 3360.390 ;
        RECT 472.020 3360.380 475.020 3360.390 ;
        RECT 652.020 3360.380 655.020 3360.390 ;
        RECT 832.020 3360.380 835.020 3360.390 ;
        RECT 1012.020 3360.380 1015.020 3360.390 ;
        RECT 1192.020 3360.380 1195.020 3360.390 ;
        RECT 1372.020 3360.380 1375.020 3360.390 ;
        RECT 1552.020 3360.380 1555.020 3360.390 ;
        RECT 1732.020 3360.380 1735.020 3360.390 ;
        RECT 1912.020 3360.380 1915.020 3360.390 ;
        RECT 2092.020 3360.380 2095.020 3360.390 ;
        RECT 2272.020 3360.380 2275.020 3360.390 ;
        RECT 2452.020 3360.380 2455.020 3360.390 ;
        RECT 2632.020 3360.380 2635.020 3360.390 ;
        RECT 2812.020 3360.380 2815.020 3360.390 ;
        RECT 2940.400 3360.380 2943.400 3360.390 ;
        RECT -23.780 3357.380 2943.400 3360.380 ;
        RECT -23.780 3357.370 -20.780 3357.380 ;
        RECT 112.020 3357.370 115.020 3357.380 ;
        RECT 292.020 3357.370 295.020 3357.380 ;
        RECT 472.020 3357.370 475.020 3357.380 ;
        RECT 652.020 3357.370 655.020 3357.380 ;
        RECT 832.020 3357.370 835.020 3357.380 ;
        RECT 1012.020 3357.370 1015.020 3357.380 ;
        RECT 1192.020 3357.370 1195.020 3357.380 ;
        RECT 1372.020 3357.370 1375.020 3357.380 ;
        RECT 1552.020 3357.370 1555.020 3357.380 ;
        RECT 1732.020 3357.370 1735.020 3357.380 ;
        RECT 1912.020 3357.370 1915.020 3357.380 ;
        RECT 2092.020 3357.370 2095.020 3357.380 ;
        RECT 2272.020 3357.370 2275.020 3357.380 ;
        RECT 2452.020 3357.370 2455.020 3357.380 ;
        RECT 2632.020 3357.370 2635.020 3357.380 ;
        RECT 2812.020 3357.370 2815.020 3357.380 ;
        RECT 2940.400 3357.370 2943.400 3357.380 ;
        RECT -23.780 3180.380 -20.780 3180.390 ;
        RECT 112.020 3180.380 115.020 3180.390 ;
        RECT 292.020 3180.380 295.020 3180.390 ;
        RECT 472.020 3180.380 475.020 3180.390 ;
        RECT 652.020 3180.380 655.020 3180.390 ;
        RECT 832.020 3180.380 835.020 3180.390 ;
        RECT 1012.020 3180.380 1015.020 3180.390 ;
        RECT 1192.020 3180.380 1195.020 3180.390 ;
        RECT 1372.020 3180.380 1375.020 3180.390 ;
        RECT 1552.020 3180.380 1555.020 3180.390 ;
        RECT 1732.020 3180.380 1735.020 3180.390 ;
        RECT 1912.020 3180.380 1915.020 3180.390 ;
        RECT 2092.020 3180.380 2095.020 3180.390 ;
        RECT 2272.020 3180.380 2275.020 3180.390 ;
        RECT 2452.020 3180.380 2455.020 3180.390 ;
        RECT 2632.020 3180.380 2635.020 3180.390 ;
        RECT 2812.020 3180.380 2815.020 3180.390 ;
        RECT 2940.400 3180.380 2943.400 3180.390 ;
        RECT -23.780 3177.380 2943.400 3180.380 ;
        RECT -23.780 3177.370 -20.780 3177.380 ;
        RECT 112.020 3177.370 115.020 3177.380 ;
        RECT 292.020 3177.370 295.020 3177.380 ;
        RECT 472.020 3177.370 475.020 3177.380 ;
        RECT 652.020 3177.370 655.020 3177.380 ;
        RECT 832.020 3177.370 835.020 3177.380 ;
        RECT 1012.020 3177.370 1015.020 3177.380 ;
        RECT 1192.020 3177.370 1195.020 3177.380 ;
        RECT 1372.020 3177.370 1375.020 3177.380 ;
        RECT 1552.020 3177.370 1555.020 3177.380 ;
        RECT 1732.020 3177.370 1735.020 3177.380 ;
        RECT 1912.020 3177.370 1915.020 3177.380 ;
        RECT 2092.020 3177.370 2095.020 3177.380 ;
        RECT 2272.020 3177.370 2275.020 3177.380 ;
        RECT 2452.020 3177.370 2455.020 3177.380 ;
        RECT 2632.020 3177.370 2635.020 3177.380 ;
        RECT 2812.020 3177.370 2815.020 3177.380 ;
        RECT 2940.400 3177.370 2943.400 3177.380 ;
        RECT -23.780 3000.380 -20.780 3000.390 ;
        RECT 112.020 3000.380 115.020 3000.390 ;
        RECT 292.020 3000.380 295.020 3000.390 ;
        RECT 472.020 3000.380 475.020 3000.390 ;
        RECT 652.020 3000.380 655.020 3000.390 ;
        RECT 832.020 3000.380 835.020 3000.390 ;
        RECT 1012.020 3000.380 1015.020 3000.390 ;
        RECT 1192.020 3000.380 1195.020 3000.390 ;
        RECT 1372.020 3000.380 1375.020 3000.390 ;
        RECT 1552.020 3000.380 1555.020 3000.390 ;
        RECT 1732.020 3000.380 1735.020 3000.390 ;
        RECT 1912.020 3000.380 1915.020 3000.390 ;
        RECT 2092.020 3000.380 2095.020 3000.390 ;
        RECT 2272.020 3000.380 2275.020 3000.390 ;
        RECT 2452.020 3000.380 2455.020 3000.390 ;
        RECT 2632.020 3000.380 2635.020 3000.390 ;
        RECT 2812.020 3000.380 2815.020 3000.390 ;
        RECT 2940.400 3000.380 2943.400 3000.390 ;
        RECT -23.780 2997.380 2943.400 3000.380 ;
        RECT -23.780 2997.370 -20.780 2997.380 ;
        RECT 112.020 2997.370 115.020 2997.380 ;
        RECT 292.020 2997.370 295.020 2997.380 ;
        RECT 472.020 2997.370 475.020 2997.380 ;
        RECT 652.020 2997.370 655.020 2997.380 ;
        RECT 832.020 2997.370 835.020 2997.380 ;
        RECT 1012.020 2997.370 1015.020 2997.380 ;
        RECT 1192.020 2997.370 1195.020 2997.380 ;
        RECT 1372.020 2997.370 1375.020 2997.380 ;
        RECT 1552.020 2997.370 1555.020 2997.380 ;
        RECT 1732.020 2997.370 1735.020 2997.380 ;
        RECT 1912.020 2997.370 1915.020 2997.380 ;
        RECT 2092.020 2997.370 2095.020 2997.380 ;
        RECT 2272.020 2997.370 2275.020 2997.380 ;
        RECT 2452.020 2997.370 2455.020 2997.380 ;
        RECT 2632.020 2997.370 2635.020 2997.380 ;
        RECT 2812.020 2997.370 2815.020 2997.380 ;
        RECT 2940.400 2997.370 2943.400 2997.380 ;
        RECT -23.780 2820.380 -20.780 2820.390 ;
        RECT 112.020 2820.380 115.020 2820.390 ;
        RECT 292.020 2820.380 295.020 2820.390 ;
        RECT 472.020 2820.380 475.020 2820.390 ;
        RECT 652.020 2820.380 655.020 2820.390 ;
        RECT 832.020 2820.380 835.020 2820.390 ;
        RECT 1012.020 2820.380 1015.020 2820.390 ;
        RECT 1192.020 2820.380 1195.020 2820.390 ;
        RECT 1372.020 2820.380 1375.020 2820.390 ;
        RECT 1552.020 2820.380 1555.020 2820.390 ;
        RECT 1732.020 2820.380 1735.020 2820.390 ;
        RECT 1912.020 2820.380 1915.020 2820.390 ;
        RECT 2092.020 2820.380 2095.020 2820.390 ;
        RECT 2272.020 2820.380 2275.020 2820.390 ;
        RECT 2452.020 2820.380 2455.020 2820.390 ;
        RECT 2632.020 2820.380 2635.020 2820.390 ;
        RECT 2812.020 2820.380 2815.020 2820.390 ;
        RECT 2940.400 2820.380 2943.400 2820.390 ;
        RECT -23.780 2817.380 2943.400 2820.380 ;
        RECT -23.780 2817.370 -20.780 2817.380 ;
        RECT 112.020 2817.370 115.020 2817.380 ;
        RECT 292.020 2817.370 295.020 2817.380 ;
        RECT 472.020 2817.370 475.020 2817.380 ;
        RECT 652.020 2817.370 655.020 2817.380 ;
        RECT 832.020 2817.370 835.020 2817.380 ;
        RECT 1012.020 2817.370 1015.020 2817.380 ;
        RECT 1192.020 2817.370 1195.020 2817.380 ;
        RECT 1372.020 2817.370 1375.020 2817.380 ;
        RECT 1552.020 2817.370 1555.020 2817.380 ;
        RECT 1732.020 2817.370 1735.020 2817.380 ;
        RECT 1912.020 2817.370 1915.020 2817.380 ;
        RECT 2092.020 2817.370 2095.020 2817.380 ;
        RECT 2272.020 2817.370 2275.020 2817.380 ;
        RECT 2452.020 2817.370 2455.020 2817.380 ;
        RECT 2632.020 2817.370 2635.020 2817.380 ;
        RECT 2812.020 2817.370 2815.020 2817.380 ;
        RECT 2940.400 2817.370 2943.400 2817.380 ;
        RECT -23.780 2640.380 -20.780 2640.390 ;
        RECT 112.020 2640.380 115.020 2640.390 ;
        RECT 292.020 2640.380 295.020 2640.390 ;
        RECT 472.020 2640.380 475.020 2640.390 ;
        RECT 652.020 2640.380 655.020 2640.390 ;
        RECT 832.020 2640.380 835.020 2640.390 ;
        RECT 1012.020 2640.380 1015.020 2640.390 ;
        RECT 1192.020 2640.380 1195.020 2640.390 ;
        RECT 1372.020 2640.380 1375.020 2640.390 ;
        RECT 1552.020 2640.380 1555.020 2640.390 ;
        RECT 1732.020 2640.380 1735.020 2640.390 ;
        RECT 1912.020 2640.380 1915.020 2640.390 ;
        RECT 2092.020 2640.380 2095.020 2640.390 ;
        RECT 2272.020 2640.380 2275.020 2640.390 ;
        RECT 2452.020 2640.380 2455.020 2640.390 ;
        RECT 2632.020 2640.380 2635.020 2640.390 ;
        RECT 2812.020 2640.380 2815.020 2640.390 ;
        RECT 2940.400 2640.380 2943.400 2640.390 ;
        RECT -23.780 2637.380 2943.400 2640.380 ;
        RECT -23.780 2637.370 -20.780 2637.380 ;
        RECT 112.020 2637.370 115.020 2637.380 ;
        RECT 292.020 2637.370 295.020 2637.380 ;
        RECT 472.020 2637.370 475.020 2637.380 ;
        RECT 652.020 2637.370 655.020 2637.380 ;
        RECT 832.020 2637.370 835.020 2637.380 ;
        RECT 1012.020 2637.370 1015.020 2637.380 ;
        RECT 1192.020 2637.370 1195.020 2637.380 ;
        RECT 1372.020 2637.370 1375.020 2637.380 ;
        RECT 1552.020 2637.370 1555.020 2637.380 ;
        RECT 1732.020 2637.370 1735.020 2637.380 ;
        RECT 1912.020 2637.370 1915.020 2637.380 ;
        RECT 2092.020 2637.370 2095.020 2637.380 ;
        RECT 2272.020 2637.370 2275.020 2637.380 ;
        RECT 2452.020 2637.370 2455.020 2637.380 ;
        RECT 2632.020 2637.370 2635.020 2637.380 ;
        RECT 2812.020 2637.370 2815.020 2637.380 ;
        RECT 2940.400 2637.370 2943.400 2637.380 ;
        RECT -23.780 2460.380 -20.780 2460.390 ;
        RECT 112.020 2460.380 115.020 2460.390 ;
        RECT 292.020 2460.380 295.020 2460.390 ;
        RECT 472.020 2460.380 475.020 2460.390 ;
        RECT 652.020 2460.380 655.020 2460.390 ;
        RECT 832.020 2460.380 835.020 2460.390 ;
        RECT 1012.020 2460.380 1015.020 2460.390 ;
        RECT 1192.020 2460.380 1195.020 2460.390 ;
        RECT 1372.020 2460.380 1375.020 2460.390 ;
        RECT 1552.020 2460.380 1555.020 2460.390 ;
        RECT 1732.020 2460.380 1735.020 2460.390 ;
        RECT 1912.020 2460.380 1915.020 2460.390 ;
        RECT 2092.020 2460.380 2095.020 2460.390 ;
        RECT 2272.020 2460.380 2275.020 2460.390 ;
        RECT 2452.020 2460.380 2455.020 2460.390 ;
        RECT 2632.020 2460.380 2635.020 2460.390 ;
        RECT 2812.020 2460.380 2815.020 2460.390 ;
        RECT 2940.400 2460.380 2943.400 2460.390 ;
        RECT -23.780 2457.380 2943.400 2460.380 ;
        RECT -23.780 2457.370 -20.780 2457.380 ;
        RECT 112.020 2457.370 115.020 2457.380 ;
        RECT 292.020 2457.370 295.020 2457.380 ;
        RECT 472.020 2457.370 475.020 2457.380 ;
        RECT 652.020 2457.370 655.020 2457.380 ;
        RECT 832.020 2457.370 835.020 2457.380 ;
        RECT 1012.020 2457.370 1015.020 2457.380 ;
        RECT 1192.020 2457.370 1195.020 2457.380 ;
        RECT 1372.020 2457.370 1375.020 2457.380 ;
        RECT 1552.020 2457.370 1555.020 2457.380 ;
        RECT 1732.020 2457.370 1735.020 2457.380 ;
        RECT 1912.020 2457.370 1915.020 2457.380 ;
        RECT 2092.020 2457.370 2095.020 2457.380 ;
        RECT 2272.020 2457.370 2275.020 2457.380 ;
        RECT 2452.020 2457.370 2455.020 2457.380 ;
        RECT 2632.020 2457.370 2635.020 2457.380 ;
        RECT 2812.020 2457.370 2815.020 2457.380 ;
        RECT 2940.400 2457.370 2943.400 2457.380 ;
        RECT -23.780 2280.380 -20.780 2280.390 ;
        RECT 112.020 2280.380 115.020 2280.390 ;
        RECT 292.020 2280.380 295.020 2280.390 ;
        RECT 472.020 2280.380 475.020 2280.390 ;
        RECT 652.020 2280.380 655.020 2280.390 ;
        RECT 832.020 2280.380 835.020 2280.390 ;
        RECT 1012.020 2280.380 1015.020 2280.390 ;
        RECT 1192.020 2280.380 1195.020 2280.390 ;
        RECT 1372.020 2280.380 1375.020 2280.390 ;
        RECT 1552.020 2280.380 1555.020 2280.390 ;
        RECT 1732.020 2280.380 1735.020 2280.390 ;
        RECT 1912.020 2280.380 1915.020 2280.390 ;
        RECT 2092.020 2280.380 2095.020 2280.390 ;
        RECT 2272.020 2280.380 2275.020 2280.390 ;
        RECT 2452.020 2280.380 2455.020 2280.390 ;
        RECT 2632.020 2280.380 2635.020 2280.390 ;
        RECT 2812.020 2280.380 2815.020 2280.390 ;
        RECT 2940.400 2280.380 2943.400 2280.390 ;
        RECT -23.780 2277.380 2943.400 2280.380 ;
        RECT -23.780 2277.370 -20.780 2277.380 ;
        RECT 112.020 2277.370 115.020 2277.380 ;
        RECT 292.020 2277.370 295.020 2277.380 ;
        RECT 472.020 2277.370 475.020 2277.380 ;
        RECT 652.020 2277.370 655.020 2277.380 ;
        RECT 832.020 2277.370 835.020 2277.380 ;
        RECT 1012.020 2277.370 1015.020 2277.380 ;
        RECT 1192.020 2277.370 1195.020 2277.380 ;
        RECT 1372.020 2277.370 1375.020 2277.380 ;
        RECT 1552.020 2277.370 1555.020 2277.380 ;
        RECT 1732.020 2277.370 1735.020 2277.380 ;
        RECT 1912.020 2277.370 1915.020 2277.380 ;
        RECT 2092.020 2277.370 2095.020 2277.380 ;
        RECT 2272.020 2277.370 2275.020 2277.380 ;
        RECT 2452.020 2277.370 2455.020 2277.380 ;
        RECT 2632.020 2277.370 2635.020 2277.380 ;
        RECT 2812.020 2277.370 2815.020 2277.380 ;
        RECT 2940.400 2277.370 2943.400 2277.380 ;
        RECT -23.780 2100.380 -20.780 2100.390 ;
        RECT 112.020 2100.380 115.020 2100.390 ;
        RECT 292.020 2100.380 295.020 2100.390 ;
        RECT 472.020 2100.380 475.020 2100.390 ;
        RECT 652.020 2100.380 655.020 2100.390 ;
        RECT 832.020 2100.380 835.020 2100.390 ;
        RECT 1012.020 2100.380 1015.020 2100.390 ;
        RECT 1192.020 2100.380 1195.020 2100.390 ;
        RECT 1372.020 2100.380 1375.020 2100.390 ;
        RECT 1552.020 2100.380 1555.020 2100.390 ;
        RECT 1732.020 2100.380 1735.020 2100.390 ;
        RECT 1912.020 2100.380 1915.020 2100.390 ;
        RECT 2092.020 2100.380 2095.020 2100.390 ;
        RECT 2272.020 2100.380 2275.020 2100.390 ;
        RECT 2452.020 2100.380 2455.020 2100.390 ;
        RECT 2632.020 2100.380 2635.020 2100.390 ;
        RECT 2812.020 2100.380 2815.020 2100.390 ;
        RECT 2940.400 2100.380 2943.400 2100.390 ;
        RECT -23.780 2097.380 2943.400 2100.380 ;
        RECT -23.780 2097.370 -20.780 2097.380 ;
        RECT 112.020 2097.370 115.020 2097.380 ;
        RECT 292.020 2097.370 295.020 2097.380 ;
        RECT 472.020 2097.370 475.020 2097.380 ;
        RECT 652.020 2097.370 655.020 2097.380 ;
        RECT 832.020 2097.370 835.020 2097.380 ;
        RECT 1012.020 2097.370 1015.020 2097.380 ;
        RECT 1192.020 2097.370 1195.020 2097.380 ;
        RECT 1372.020 2097.370 1375.020 2097.380 ;
        RECT 1552.020 2097.370 1555.020 2097.380 ;
        RECT 1732.020 2097.370 1735.020 2097.380 ;
        RECT 1912.020 2097.370 1915.020 2097.380 ;
        RECT 2092.020 2097.370 2095.020 2097.380 ;
        RECT 2272.020 2097.370 2275.020 2097.380 ;
        RECT 2452.020 2097.370 2455.020 2097.380 ;
        RECT 2632.020 2097.370 2635.020 2097.380 ;
        RECT 2812.020 2097.370 2815.020 2097.380 ;
        RECT 2940.400 2097.370 2943.400 2097.380 ;
        RECT -23.780 1920.380 -20.780 1920.390 ;
        RECT 112.020 1920.380 115.020 1920.390 ;
        RECT 292.020 1920.380 295.020 1920.390 ;
        RECT 472.020 1920.380 475.020 1920.390 ;
        RECT 652.020 1920.380 655.020 1920.390 ;
        RECT 832.020 1920.380 835.020 1920.390 ;
        RECT 1012.020 1920.380 1015.020 1920.390 ;
        RECT 1192.020 1920.380 1195.020 1920.390 ;
        RECT 1372.020 1920.380 1375.020 1920.390 ;
        RECT 1552.020 1920.380 1555.020 1920.390 ;
        RECT 1732.020 1920.380 1735.020 1920.390 ;
        RECT 1912.020 1920.380 1915.020 1920.390 ;
        RECT 2092.020 1920.380 2095.020 1920.390 ;
        RECT 2272.020 1920.380 2275.020 1920.390 ;
        RECT 2452.020 1920.380 2455.020 1920.390 ;
        RECT 2632.020 1920.380 2635.020 1920.390 ;
        RECT 2812.020 1920.380 2815.020 1920.390 ;
        RECT 2940.400 1920.380 2943.400 1920.390 ;
        RECT -23.780 1917.380 2943.400 1920.380 ;
        RECT -23.780 1917.370 -20.780 1917.380 ;
        RECT 112.020 1917.370 115.020 1917.380 ;
        RECT 292.020 1917.370 295.020 1917.380 ;
        RECT 472.020 1917.370 475.020 1917.380 ;
        RECT 652.020 1917.370 655.020 1917.380 ;
        RECT 832.020 1917.370 835.020 1917.380 ;
        RECT 1012.020 1917.370 1015.020 1917.380 ;
        RECT 1192.020 1917.370 1195.020 1917.380 ;
        RECT 1372.020 1917.370 1375.020 1917.380 ;
        RECT 1552.020 1917.370 1555.020 1917.380 ;
        RECT 1732.020 1917.370 1735.020 1917.380 ;
        RECT 1912.020 1917.370 1915.020 1917.380 ;
        RECT 2092.020 1917.370 2095.020 1917.380 ;
        RECT 2272.020 1917.370 2275.020 1917.380 ;
        RECT 2452.020 1917.370 2455.020 1917.380 ;
        RECT 2632.020 1917.370 2635.020 1917.380 ;
        RECT 2812.020 1917.370 2815.020 1917.380 ;
        RECT 2940.400 1917.370 2943.400 1917.380 ;
        RECT -23.780 1740.380 -20.780 1740.390 ;
        RECT 112.020 1740.380 115.020 1740.390 ;
        RECT 292.020 1740.380 295.020 1740.390 ;
        RECT 472.020 1740.380 475.020 1740.390 ;
        RECT 652.020 1740.380 655.020 1740.390 ;
        RECT 832.020 1740.380 835.020 1740.390 ;
        RECT 1012.020 1740.380 1015.020 1740.390 ;
        RECT 1192.020 1740.380 1195.020 1740.390 ;
        RECT 1372.020 1740.380 1375.020 1740.390 ;
        RECT 1552.020 1740.380 1555.020 1740.390 ;
        RECT 1732.020 1740.380 1735.020 1740.390 ;
        RECT 1912.020 1740.380 1915.020 1740.390 ;
        RECT 2092.020 1740.380 2095.020 1740.390 ;
        RECT 2272.020 1740.380 2275.020 1740.390 ;
        RECT 2452.020 1740.380 2455.020 1740.390 ;
        RECT 2632.020 1740.380 2635.020 1740.390 ;
        RECT 2812.020 1740.380 2815.020 1740.390 ;
        RECT 2940.400 1740.380 2943.400 1740.390 ;
        RECT -23.780 1737.380 2943.400 1740.380 ;
        RECT -23.780 1737.370 -20.780 1737.380 ;
        RECT 112.020 1737.370 115.020 1737.380 ;
        RECT 292.020 1737.370 295.020 1737.380 ;
        RECT 472.020 1737.370 475.020 1737.380 ;
        RECT 652.020 1737.370 655.020 1737.380 ;
        RECT 832.020 1737.370 835.020 1737.380 ;
        RECT 1012.020 1737.370 1015.020 1737.380 ;
        RECT 1192.020 1737.370 1195.020 1737.380 ;
        RECT 1372.020 1737.370 1375.020 1737.380 ;
        RECT 1552.020 1737.370 1555.020 1737.380 ;
        RECT 1732.020 1737.370 1735.020 1737.380 ;
        RECT 1912.020 1737.370 1915.020 1737.380 ;
        RECT 2092.020 1737.370 2095.020 1737.380 ;
        RECT 2272.020 1737.370 2275.020 1737.380 ;
        RECT 2452.020 1737.370 2455.020 1737.380 ;
        RECT 2632.020 1737.370 2635.020 1737.380 ;
        RECT 2812.020 1737.370 2815.020 1737.380 ;
        RECT 2940.400 1737.370 2943.400 1737.380 ;
        RECT -23.780 1560.380 -20.780 1560.390 ;
        RECT 112.020 1560.380 115.020 1560.390 ;
        RECT 292.020 1560.380 295.020 1560.390 ;
        RECT 472.020 1560.380 475.020 1560.390 ;
        RECT 652.020 1560.380 655.020 1560.390 ;
        RECT 832.020 1560.380 835.020 1560.390 ;
        RECT 1012.020 1560.380 1015.020 1560.390 ;
        RECT 1192.020 1560.380 1195.020 1560.390 ;
        RECT 1372.020 1560.380 1375.020 1560.390 ;
        RECT 1552.020 1560.380 1555.020 1560.390 ;
        RECT 1732.020 1560.380 1735.020 1560.390 ;
        RECT 1912.020 1560.380 1915.020 1560.390 ;
        RECT 2092.020 1560.380 2095.020 1560.390 ;
        RECT 2272.020 1560.380 2275.020 1560.390 ;
        RECT 2452.020 1560.380 2455.020 1560.390 ;
        RECT 2632.020 1560.380 2635.020 1560.390 ;
        RECT 2812.020 1560.380 2815.020 1560.390 ;
        RECT 2940.400 1560.380 2943.400 1560.390 ;
        RECT -23.780 1557.380 2943.400 1560.380 ;
        RECT -23.780 1557.370 -20.780 1557.380 ;
        RECT 112.020 1557.370 115.020 1557.380 ;
        RECT 292.020 1557.370 295.020 1557.380 ;
        RECT 472.020 1557.370 475.020 1557.380 ;
        RECT 652.020 1557.370 655.020 1557.380 ;
        RECT 832.020 1557.370 835.020 1557.380 ;
        RECT 1012.020 1557.370 1015.020 1557.380 ;
        RECT 1192.020 1557.370 1195.020 1557.380 ;
        RECT 1372.020 1557.370 1375.020 1557.380 ;
        RECT 1552.020 1557.370 1555.020 1557.380 ;
        RECT 1732.020 1557.370 1735.020 1557.380 ;
        RECT 1912.020 1557.370 1915.020 1557.380 ;
        RECT 2092.020 1557.370 2095.020 1557.380 ;
        RECT 2272.020 1557.370 2275.020 1557.380 ;
        RECT 2452.020 1557.370 2455.020 1557.380 ;
        RECT 2632.020 1557.370 2635.020 1557.380 ;
        RECT 2812.020 1557.370 2815.020 1557.380 ;
        RECT 2940.400 1557.370 2943.400 1557.380 ;
        RECT -23.780 1380.380 -20.780 1380.390 ;
        RECT 112.020 1380.380 115.020 1380.390 ;
        RECT 292.020 1380.380 295.020 1380.390 ;
        RECT 472.020 1380.380 475.020 1380.390 ;
        RECT 652.020 1380.380 655.020 1380.390 ;
        RECT 832.020 1380.380 835.020 1380.390 ;
        RECT 1012.020 1380.380 1015.020 1380.390 ;
        RECT 1192.020 1380.380 1195.020 1380.390 ;
        RECT 1372.020 1380.380 1375.020 1380.390 ;
        RECT 1552.020 1380.380 1555.020 1380.390 ;
        RECT 1732.020 1380.380 1735.020 1380.390 ;
        RECT 1912.020 1380.380 1915.020 1380.390 ;
        RECT 2092.020 1380.380 2095.020 1380.390 ;
        RECT 2272.020 1380.380 2275.020 1380.390 ;
        RECT 2452.020 1380.380 2455.020 1380.390 ;
        RECT 2632.020 1380.380 2635.020 1380.390 ;
        RECT 2812.020 1380.380 2815.020 1380.390 ;
        RECT 2940.400 1380.380 2943.400 1380.390 ;
        RECT -23.780 1377.380 2943.400 1380.380 ;
        RECT -23.780 1377.370 -20.780 1377.380 ;
        RECT 112.020 1377.370 115.020 1377.380 ;
        RECT 292.020 1377.370 295.020 1377.380 ;
        RECT 472.020 1377.370 475.020 1377.380 ;
        RECT 652.020 1377.370 655.020 1377.380 ;
        RECT 832.020 1377.370 835.020 1377.380 ;
        RECT 1012.020 1377.370 1015.020 1377.380 ;
        RECT 1192.020 1377.370 1195.020 1377.380 ;
        RECT 1372.020 1377.370 1375.020 1377.380 ;
        RECT 1552.020 1377.370 1555.020 1377.380 ;
        RECT 1732.020 1377.370 1735.020 1377.380 ;
        RECT 1912.020 1377.370 1915.020 1377.380 ;
        RECT 2092.020 1377.370 2095.020 1377.380 ;
        RECT 2272.020 1377.370 2275.020 1377.380 ;
        RECT 2452.020 1377.370 2455.020 1377.380 ;
        RECT 2632.020 1377.370 2635.020 1377.380 ;
        RECT 2812.020 1377.370 2815.020 1377.380 ;
        RECT 2940.400 1377.370 2943.400 1377.380 ;
        RECT -23.780 1200.380 -20.780 1200.390 ;
        RECT 112.020 1200.380 115.020 1200.390 ;
        RECT 292.020 1200.380 295.020 1200.390 ;
        RECT 472.020 1200.380 475.020 1200.390 ;
        RECT 652.020 1200.380 655.020 1200.390 ;
        RECT 832.020 1200.380 835.020 1200.390 ;
        RECT 1012.020 1200.380 1015.020 1200.390 ;
        RECT 1192.020 1200.380 1195.020 1200.390 ;
        RECT 1372.020 1200.380 1375.020 1200.390 ;
        RECT 1552.020 1200.380 1555.020 1200.390 ;
        RECT 1732.020 1200.380 1735.020 1200.390 ;
        RECT 1912.020 1200.380 1915.020 1200.390 ;
        RECT 2092.020 1200.380 2095.020 1200.390 ;
        RECT 2272.020 1200.380 2275.020 1200.390 ;
        RECT 2452.020 1200.380 2455.020 1200.390 ;
        RECT 2632.020 1200.380 2635.020 1200.390 ;
        RECT 2812.020 1200.380 2815.020 1200.390 ;
        RECT 2940.400 1200.380 2943.400 1200.390 ;
        RECT -23.780 1197.380 2943.400 1200.380 ;
        RECT -23.780 1197.370 -20.780 1197.380 ;
        RECT 112.020 1197.370 115.020 1197.380 ;
        RECT 292.020 1197.370 295.020 1197.380 ;
        RECT 472.020 1197.370 475.020 1197.380 ;
        RECT 652.020 1197.370 655.020 1197.380 ;
        RECT 832.020 1197.370 835.020 1197.380 ;
        RECT 1012.020 1197.370 1015.020 1197.380 ;
        RECT 1192.020 1197.370 1195.020 1197.380 ;
        RECT 1372.020 1197.370 1375.020 1197.380 ;
        RECT 1552.020 1197.370 1555.020 1197.380 ;
        RECT 1732.020 1197.370 1735.020 1197.380 ;
        RECT 1912.020 1197.370 1915.020 1197.380 ;
        RECT 2092.020 1197.370 2095.020 1197.380 ;
        RECT 2272.020 1197.370 2275.020 1197.380 ;
        RECT 2452.020 1197.370 2455.020 1197.380 ;
        RECT 2632.020 1197.370 2635.020 1197.380 ;
        RECT 2812.020 1197.370 2815.020 1197.380 ;
        RECT 2940.400 1197.370 2943.400 1197.380 ;
        RECT -23.780 1020.380 -20.780 1020.390 ;
        RECT 112.020 1020.380 115.020 1020.390 ;
        RECT 292.020 1020.380 295.020 1020.390 ;
        RECT 472.020 1020.380 475.020 1020.390 ;
        RECT 652.020 1020.380 655.020 1020.390 ;
        RECT 832.020 1020.380 835.020 1020.390 ;
        RECT 1012.020 1020.380 1015.020 1020.390 ;
        RECT 1192.020 1020.380 1195.020 1020.390 ;
        RECT 1372.020 1020.380 1375.020 1020.390 ;
        RECT 1552.020 1020.380 1555.020 1020.390 ;
        RECT 1732.020 1020.380 1735.020 1020.390 ;
        RECT 1912.020 1020.380 1915.020 1020.390 ;
        RECT 2092.020 1020.380 2095.020 1020.390 ;
        RECT 2272.020 1020.380 2275.020 1020.390 ;
        RECT 2452.020 1020.380 2455.020 1020.390 ;
        RECT 2632.020 1020.380 2635.020 1020.390 ;
        RECT 2812.020 1020.380 2815.020 1020.390 ;
        RECT 2940.400 1020.380 2943.400 1020.390 ;
        RECT -23.780 1017.380 2943.400 1020.380 ;
        RECT -23.780 1017.370 -20.780 1017.380 ;
        RECT 112.020 1017.370 115.020 1017.380 ;
        RECT 292.020 1017.370 295.020 1017.380 ;
        RECT 472.020 1017.370 475.020 1017.380 ;
        RECT 652.020 1017.370 655.020 1017.380 ;
        RECT 832.020 1017.370 835.020 1017.380 ;
        RECT 1012.020 1017.370 1015.020 1017.380 ;
        RECT 1192.020 1017.370 1195.020 1017.380 ;
        RECT 1372.020 1017.370 1375.020 1017.380 ;
        RECT 1552.020 1017.370 1555.020 1017.380 ;
        RECT 1732.020 1017.370 1735.020 1017.380 ;
        RECT 1912.020 1017.370 1915.020 1017.380 ;
        RECT 2092.020 1017.370 2095.020 1017.380 ;
        RECT 2272.020 1017.370 2275.020 1017.380 ;
        RECT 2452.020 1017.370 2455.020 1017.380 ;
        RECT 2632.020 1017.370 2635.020 1017.380 ;
        RECT 2812.020 1017.370 2815.020 1017.380 ;
        RECT 2940.400 1017.370 2943.400 1017.380 ;
        RECT -23.780 840.380 -20.780 840.390 ;
        RECT 112.020 840.380 115.020 840.390 ;
        RECT 292.020 840.380 295.020 840.390 ;
        RECT 472.020 840.380 475.020 840.390 ;
        RECT 652.020 840.380 655.020 840.390 ;
        RECT 832.020 840.380 835.020 840.390 ;
        RECT 1012.020 840.380 1015.020 840.390 ;
        RECT 1192.020 840.380 1195.020 840.390 ;
        RECT 1372.020 840.380 1375.020 840.390 ;
        RECT 1552.020 840.380 1555.020 840.390 ;
        RECT 1732.020 840.380 1735.020 840.390 ;
        RECT 1912.020 840.380 1915.020 840.390 ;
        RECT 2092.020 840.380 2095.020 840.390 ;
        RECT 2272.020 840.380 2275.020 840.390 ;
        RECT 2452.020 840.380 2455.020 840.390 ;
        RECT 2632.020 840.380 2635.020 840.390 ;
        RECT 2812.020 840.380 2815.020 840.390 ;
        RECT 2940.400 840.380 2943.400 840.390 ;
        RECT -23.780 837.380 2943.400 840.380 ;
        RECT -23.780 837.370 -20.780 837.380 ;
        RECT 112.020 837.370 115.020 837.380 ;
        RECT 292.020 837.370 295.020 837.380 ;
        RECT 472.020 837.370 475.020 837.380 ;
        RECT 652.020 837.370 655.020 837.380 ;
        RECT 832.020 837.370 835.020 837.380 ;
        RECT 1012.020 837.370 1015.020 837.380 ;
        RECT 1192.020 837.370 1195.020 837.380 ;
        RECT 1372.020 837.370 1375.020 837.380 ;
        RECT 1552.020 837.370 1555.020 837.380 ;
        RECT 1732.020 837.370 1735.020 837.380 ;
        RECT 1912.020 837.370 1915.020 837.380 ;
        RECT 2092.020 837.370 2095.020 837.380 ;
        RECT 2272.020 837.370 2275.020 837.380 ;
        RECT 2452.020 837.370 2455.020 837.380 ;
        RECT 2632.020 837.370 2635.020 837.380 ;
        RECT 2812.020 837.370 2815.020 837.380 ;
        RECT 2940.400 837.370 2943.400 837.380 ;
        RECT -23.780 660.380 -20.780 660.390 ;
        RECT 112.020 660.380 115.020 660.390 ;
        RECT 292.020 660.380 295.020 660.390 ;
        RECT 472.020 660.380 475.020 660.390 ;
        RECT 652.020 660.380 655.020 660.390 ;
        RECT 832.020 660.380 835.020 660.390 ;
        RECT 1012.020 660.380 1015.020 660.390 ;
        RECT 1192.020 660.380 1195.020 660.390 ;
        RECT 1372.020 660.380 1375.020 660.390 ;
        RECT 1552.020 660.380 1555.020 660.390 ;
        RECT 1732.020 660.380 1735.020 660.390 ;
        RECT 1912.020 660.380 1915.020 660.390 ;
        RECT 2092.020 660.380 2095.020 660.390 ;
        RECT 2272.020 660.380 2275.020 660.390 ;
        RECT 2452.020 660.380 2455.020 660.390 ;
        RECT 2632.020 660.380 2635.020 660.390 ;
        RECT 2812.020 660.380 2815.020 660.390 ;
        RECT 2940.400 660.380 2943.400 660.390 ;
        RECT -23.780 657.380 2943.400 660.380 ;
        RECT -23.780 657.370 -20.780 657.380 ;
        RECT 112.020 657.370 115.020 657.380 ;
        RECT 292.020 657.370 295.020 657.380 ;
        RECT 472.020 657.370 475.020 657.380 ;
        RECT 652.020 657.370 655.020 657.380 ;
        RECT 832.020 657.370 835.020 657.380 ;
        RECT 1012.020 657.370 1015.020 657.380 ;
        RECT 1192.020 657.370 1195.020 657.380 ;
        RECT 1372.020 657.370 1375.020 657.380 ;
        RECT 1552.020 657.370 1555.020 657.380 ;
        RECT 1732.020 657.370 1735.020 657.380 ;
        RECT 1912.020 657.370 1915.020 657.380 ;
        RECT 2092.020 657.370 2095.020 657.380 ;
        RECT 2272.020 657.370 2275.020 657.380 ;
        RECT 2452.020 657.370 2455.020 657.380 ;
        RECT 2632.020 657.370 2635.020 657.380 ;
        RECT 2812.020 657.370 2815.020 657.380 ;
        RECT 2940.400 657.370 2943.400 657.380 ;
        RECT -23.780 480.380 -20.780 480.390 ;
        RECT 112.020 480.380 115.020 480.390 ;
        RECT 292.020 480.380 295.020 480.390 ;
        RECT 472.020 480.380 475.020 480.390 ;
        RECT 652.020 480.380 655.020 480.390 ;
        RECT 832.020 480.380 835.020 480.390 ;
        RECT 1012.020 480.380 1015.020 480.390 ;
        RECT 1192.020 480.380 1195.020 480.390 ;
        RECT 1372.020 480.380 1375.020 480.390 ;
        RECT 1552.020 480.380 1555.020 480.390 ;
        RECT 1732.020 480.380 1735.020 480.390 ;
        RECT 1912.020 480.380 1915.020 480.390 ;
        RECT 2092.020 480.380 2095.020 480.390 ;
        RECT 2272.020 480.380 2275.020 480.390 ;
        RECT 2452.020 480.380 2455.020 480.390 ;
        RECT 2632.020 480.380 2635.020 480.390 ;
        RECT 2812.020 480.380 2815.020 480.390 ;
        RECT 2940.400 480.380 2943.400 480.390 ;
        RECT -23.780 477.380 2943.400 480.380 ;
        RECT -23.780 477.370 -20.780 477.380 ;
        RECT 112.020 477.370 115.020 477.380 ;
        RECT 292.020 477.370 295.020 477.380 ;
        RECT 472.020 477.370 475.020 477.380 ;
        RECT 652.020 477.370 655.020 477.380 ;
        RECT 832.020 477.370 835.020 477.380 ;
        RECT 1012.020 477.370 1015.020 477.380 ;
        RECT 1192.020 477.370 1195.020 477.380 ;
        RECT 1372.020 477.370 1375.020 477.380 ;
        RECT 1552.020 477.370 1555.020 477.380 ;
        RECT 1732.020 477.370 1735.020 477.380 ;
        RECT 1912.020 477.370 1915.020 477.380 ;
        RECT 2092.020 477.370 2095.020 477.380 ;
        RECT 2272.020 477.370 2275.020 477.380 ;
        RECT 2452.020 477.370 2455.020 477.380 ;
        RECT 2632.020 477.370 2635.020 477.380 ;
        RECT 2812.020 477.370 2815.020 477.380 ;
        RECT 2940.400 477.370 2943.400 477.380 ;
        RECT -23.780 300.380 -20.780 300.390 ;
        RECT 112.020 300.380 115.020 300.390 ;
        RECT 292.020 300.380 295.020 300.390 ;
        RECT 472.020 300.380 475.020 300.390 ;
        RECT 652.020 300.380 655.020 300.390 ;
        RECT 832.020 300.380 835.020 300.390 ;
        RECT 1012.020 300.380 1015.020 300.390 ;
        RECT 1192.020 300.380 1195.020 300.390 ;
        RECT 1372.020 300.380 1375.020 300.390 ;
        RECT 1552.020 300.380 1555.020 300.390 ;
        RECT 1732.020 300.380 1735.020 300.390 ;
        RECT 1912.020 300.380 1915.020 300.390 ;
        RECT 2092.020 300.380 2095.020 300.390 ;
        RECT 2272.020 300.380 2275.020 300.390 ;
        RECT 2452.020 300.380 2455.020 300.390 ;
        RECT 2632.020 300.380 2635.020 300.390 ;
        RECT 2812.020 300.380 2815.020 300.390 ;
        RECT 2940.400 300.380 2943.400 300.390 ;
        RECT -23.780 297.380 2943.400 300.380 ;
        RECT -23.780 297.370 -20.780 297.380 ;
        RECT 112.020 297.370 115.020 297.380 ;
        RECT 292.020 297.370 295.020 297.380 ;
        RECT 472.020 297.370 475.020 297.380 ;
        RECT 652.020 297.370 655.020 297.380 ;
        RECT 832.020 297.370 835.020 297.380 ;
        RECT 1012.020 297.370 1015.020 297.380 ;
        RECT 1192.020 297.370 1195.020 297.380 ;
        RECT 1372.020 297.370 1375.020 297.380 ;
        RECT 1552.020 297.370 1555.020 297.380 ;
        RECT 1732.020 297.370 1735.020 297.380 ;
        RECT 1912.020 297.370 1915.020 297.380 ;
        RECT 2092.020 297.370 2095.020 297.380 ;
        RECT 2272.020 297.370 2275.020 297.380 ;
        RECT 2452.020 297.370 2455.020 297.380 ;
        RECT 2632.020 297.370 2635.020 297.380 ;
        RECT 2812.020 297.370 2815.020 297.380 ;
        RECT 2940.400 297.370 2943.400 297.380 ;
        RECT -23.780 120.380 -20.780 120.390 ;
        RECT 112.020 120.380 115.020 120.390 ;
        RECT 292.020 120.380 295.020 120.390 ;
        RECT 472.020 120.380 475.020 120.390 ;
        RECT 652.020 120.380 655.020 120.390 ;
        RECT 832.020 120.380 835.020 120.390 ;
        RECT 1012.020 120.380 1015.020 120.390 ;
        RECT 1192.020 120.380 1195.020 120.390 ;
        RECT 1372.020 120.380 1375.020 120.390 ;
        RECT 1552.020 120.380 1555.020 120.390 ;
        RECT 1732.020 120.380 1735.020 120.390 ;
        RECT 1912.020 120.380 1915.020 120.390 ;
        RECT 2092.020 120.380 2095.020 120.390 ;
        RECT 2272.020 120.380 2275.020 120.390 ;
        RECT 2452.020 120.380 2455.020 120.390 ;
        RECT 2632.020 120.380 2635.020 120.390 ;
        RECT 2812.020 120.380 2815.020 120.390 ;
        RECT 2940.400 120.380 2943.400 120.390 ;
        RECT -23.780 117.380 2943.400 120.380 ;
        RECT -23.780 117.370 -20.780 117.380 ;
        RECT 112.020 117.370 115.020 117.380 ;
        RECT 292.020 117.370 295.020 117.380 ;
        RECT 472.020 117.370 475.020 117.380 ;
        RECT 652.020 117.370 655.020 117.380 ;
        RECT 832.020 117.370 835.020 117.380 ;
        RECT 1012.020 117.370 1015.020 117.380 ;
        RECT 1192.020 117.370 1195.020 117.380 ;
        RECT 1372.020 117.370 1375.020 117.380 ;
        RECT 1552.020 117.370 1555.020 117.380 ;
        RECT 1732.020 117.370 1735.020 117.380 ;
        RECT 1912.020 117.370 1915.020 117.380 ;
        RECT 2092.020 117.370 2095.020 117.380 ;
        RECT 2272.020 117.370 2275.020 117.380 ;
        RECT 2452.020 117.370 2455.020 117.380 ;
        RECT 2632.020 117.370 2635.020 117.380 ;
        RECT 2812.020 117.370 2815.020 117.380 ;
        RECT 2940.400 117.370 2943.400 117.380 ;
        RECT -23.780 -15.420 -20.780 -15.410 ;
        RECT 112.020 -15.420 115.020 -15.410 ;
        RECT 292.020 -15.420 295.020 -15.410 ;
        RECT 472.020 -15.420 475.020 -15.410 ;
        RECT 652.020 -15.420 655.020 -15.410 ;
        RECT 832.020 -15.420 835.020 -15.410 ;
        RECT 1012.020 -15.420 1015.020 -15.410 ;
        RECT 1192.020 -15.420 1195.020 -15.410 ;
        RECT 1372.020 -15.420 1375.020 -15.410 ;
        RECT 1552.020 -15.420 1555.020 -15.410 ;
        RECT 1732.020 -15.420 1735.020 -15.410 ;
        RECT 1912.020 -15.420 1915.020 -15.410 ;
        RECT 2092.020 -15.420 2095.020 -15.410 ;
        RECT 2272.020 -15.420 2275.020 -15.410 ;
        RECT 2452.020 -15.420 2455.020 -15.410 ;
        RECT 2632.020 -15.420 2635.020 -15.410 ;
        RECT 2812.020 -15.420 2815.020 -15.410 ;
        RECT 2940.400 -15.420 2943.400 -15.410 ;
        RECT -23.780 -18.420 2943.400 -15.420 ;
        RECT -23.780 -18.430 -20.780 -18.420 ;
        RECT 112.020 -18.430 115.020 -18.420 ;
        RECT 292.020 -18.430 295.020 -18.420 ;
        RECT 472.020 -18.430 475.020 -18.420 ;
        RECT 652.020 -18.430 655.020 -18.420 ;
        RECT 832.020 -18.430 835.020 -18.420 ;
        RECT 1012.020 -18.430 1015.020 -18.420 ;
        RECT 1192.020 -18.430 1195.020 -18.420 ;
        RECT 1372.020 -18.430 1375.020 -18.420 ;
        RECT 1552.020 -18.430 1555.020 -18.420 ;
        RECT 1732.020 -18.430 1735.020 -18.420 ;
        RECT 1912.020 -18.430 1915.020 -18.420 ;
        RECT 2092.020 -18.430 2095.020 -18.420 ;
        RECT 2272.020 -18.430 2275.020 -18.420 ;
        RECT 2452.020 -18.430 2455.020 -18.420 ;
        RECT 2632.020 -18.430 2635.020 -18.420 ;
        RECT 2812.020 -18.430 2815.020 -18.420 ;
        RECT 2940.400 -18.430 2943.400 -18.420 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -28.380 -23.020 -25.380 3542.700 ;
        RECT 40.020 -27.620 43.020 3547.300 ;
        RECT 220.020 -27.620 223.020 3547.300 ;
        RECT 400.020 -27.620 403.020 3547.300 ;
        RECT 580.020 -27.620 583.020 3547.300 ;
        RECT 760.020 -27.620 763.020 3547.300 ;
        RECT 940.020 -27.620 943.020 3547.300 ;
        RECT 1120.020 -27.620 1123.020 3547.300 ;
        RECT 1300.020 -27.620 1303.020 3547.300 ;
        RECT 1480.020 -27.620 1483.020 3547.300 ;
        RECT 1660.020 -27.620 1663.020 3547.300 ;
        RECT 1840.020 -27.620 1843.020 3547.300 ;
        RECT 2020.020 -27.620 2023.020 3547.300 ;
        RECT 2200.020 -27.620 2203.020 3547.300 ;
        RECT 2380.020 -27.620 2383.020 3547.300 ;
        RECT 2560.020 -27.620 2563.020 3547.300 ;
        RECT 2740.020 -27.620 2743.020 3547.300 ;
        RECT 2945.000 -23.020 2948.000 3542.700 ;
      LAYER via4 ;
        RECT -27.470 3541.410 -26.290 3542.590 ;
        RECT -27.470 3539.810 -26.290 3540.990 ;
        RECT -27.470 3467.090 -26.290 3468.270 ;
        RECT -27.470 3465.490 -26.290 3466.670 ;
        RECT -27.470 3287.090 -26.290 3288.270 ;
        RECT -27.470 3285.490 -26.290 3286.670 ;
        RECT -27.470 3107.090 -26.290 3108.270 ;
        RECT -27.470 3105.490 -26.290 3106.670 ;
        RECT -27.470 2927.090 -26.290 2928.270 ;
        RECT -27.470 2925.490 -26.290 2926.670 ;
        RECT -27.470 2747.090 -26.290 2748.270 ;
        RECT -27.470 2745.490 -26.290 2746.670 ;
        RECT -27.470 2567.090 -26.290 2568.270 ;
        RECT -27.470 2565.490 -26.290 2566.670 ;
        RECT -27.470 2387.090 -26.290 2388.270 ;
        RECT -27.470 2385.490 -26.290 2386.670 ;
        RECT -27.470 2207.090 -26.290 2208.270 ;
        RECT -27.470 2205.490 -26.290 2206.670 ;
        RECT -27.470 2027.090 -26.290 2028.270 ;
        RECT -27.470 2025.490 -26.290 2026.670 ;
        RECT -27.470 1847.090 -26.290 1848.270 ;
        RECT -27.470 1845.490 -26.290 1846.670 ;
        RECT -27.470 1667.090 -26.290 1668.270 ;
        RECT -27.470 1665.490 -26.290 1666.670 ;
        RECT -27.470 1487.090 -26.290 1488.270 ;
        RECT -27.470 1485.490 -26.290 1486.670 ;
        RECT -27.470 1307.090 -26.290 1308.270 ;
        RECT -27.470 1305.490 -26.290 1306.670 ;
        RECT -27.470 1127.090 -26.290 1128.270 ;
        RECT -27.470 1125.490 -26.290 1126.670 ;
        RECT -27.470 947.090 -26.290 948.270 ;
        RECT -27.470 945.490 -26.290 946.670 ;
        RECT -27.470 767.090 -26.290 768.270 ;
        RECT -27.470 765.490 -26.290 766.670 ;
        RECT -27.470 587.090 -26.290 588.270 ;
        RECT -27.470 585.490 -26.290 586.670 ;
        RECT -27.470 407.090 -26.290 408.270 ;
        RECT -27.470 405.490 -26.290 406.670 ;
        RECT -27.470 227.090 -26.290 228.270 ;
        RECT -27.470 225.490 -26.290 226.670 ;
        RECT -27.470 47.090 -26.290 48.270 ;
        RECT -27.470 45.490 -26.290 46.670 ;
        RECT -27.470 -21.310 -26.290 -20.130 ;
        RECT -27.470 -22.910 -26.290 -21.730 ;
        RECT 40.930 3541.410 42.110 3542.590 ;
        RECT 40.930 3539.810 42.110 3540.990 ;
        RECT 40.930 3467.090 42.110 3468.270 ;
        RECT 40.930 3465.490 42.110 3466.670 ;
        RECT 40.930 3287.090 42.110 3288.270 ;
        RECT 40.930 3285.490 42.110 3286.670 ;
        RECT 40.930 3107.090 42.110 3108.270 ;
        RECT 40.930 3105.490 42.110 3106.670 ;
        RECT 40.930 2927.090 42.110 2928.270 ;
        RECT 40.930 2925.490 42.110 2926.670 ;
        RECT 40.930 2747.090 42.110 2748.270 ;
        RECT 40.930 2745.490 42.110 2746.670 ;
        RECT 40.930 2567.090 42.110 2568.270 ;
        RECT 40.930 2565.490 42.110 2566.670 ;
        RECT 40.930 2387.090 42.110 2388.270 ;
        RECT 40.930 2385.490 42.110 2386.670 ;
        RECT 40.930 2207.090 42.110 2208.270 ;
        RECT 40.930 2205.490 42.110 2206.670 ;
        RECT 40.930 2027.090 42.110 2028.270 ;
        RECT 40.930 2025.490 42.110 2026.670 ;
        RECT 40.930 1847.090 42.110 1848.270 ;
        RECT 40.930 1845.490 42.110 1846.670 ;
        RECT 40.930 1667.090 42.110 1668.270 ;
        RECT 40.930 1665.490 42.110 1666.670 ;
        RECT 40.930 1487.090 42.110 1488.270 ;
        RECT 40.930 1485.490 42.110 1486.670 ;
        RECT 40.930 1307.090 42.110 1308.270 ;
        RECT 40.930 1305.490 42.110 1306.670 ;
        RECT 40.930 1127.090 42.110 1128.270 ;
        RECT 40.930 1125.490 42.110 1126.670 ;
        RECT 40.930 947.090 42.110 948.270 ;
        RECT 40.930 945.490 42.110 946.670 ;
        RECT 40.930 767.090 42.110 768.270 ;
        RECT 40.930 765.490 42.110 766.670 ;
        RECT 40.930 587.090 42.110 588.270 ;
        RECT 40.930 585.490 42.110 586.670 ;
        RECT 40.930 407.090 42.110 408.270 ;
        RECT 40.930 405.490 42.110 406.670 ;
        RECT 40.930 227.090 42.110 228.270 ;
        RECT 40.930 225.490 42.110 226.670 ;
        RECT 40.930 47.090 42.110 48.270 ;
        RECT 40.930 45.490 42.110 46.670 ;
        RECT 40.930 -21.310 42.110 -20.130 ;
        RECT 40.930 -22.910 42.110 -21.730 ;
        RECT 220.930 3541.410 222.110 3542.590 ;
        RECT 220.930 3539.810 222.110 3540.990 ;
        RECT 220.930 3467.090 222.110 3468.270 ;
        RECT 220.930 3465.490 222.110 3466.670 ;
        RECT 220.930 3287.090 222.110 3288.270 ;
        RECT 220.930 3285.490 222.110 3286.670 ;
        RECT 220.930 3107.090 222.110 3108.270 ;
        RECT 220.930 3105.490 222.110 3106.670 ;
        RECT 220.930 2927.090 222.110 2928.270 ;
        RECT 220.930 2925.490 222.110 2926.670 ;
        RECT 220.930 2747.090 222.110 2748.270 ;
        RECT 220.930 2745.490 222.110 2746.670 ;
        RECT 220.930 2567.090 222.110 2568.270 ;
        RECT 220.930 2565.490 222.110 2566.670 ;
        RECT 220.930 2387.090 222.110 2388.270 ;
        RECT 220.930 2385.490 222.110 2386.670 ;
        RECT 220.930 2207.090 222.110 2208.270 ;
        RECT 220.930 2205.490 222.110 2206.670 ;
        RECT 220.930 2027.090 222.110 2028.270 ;
        RECT 220.930 2025.490 222.110 2026.670 ;
        RECT 220.930 1847.090 222.110 1848.270 ;
        RECT 220.930 1845.490 222.110 1846.670 ;
        RECT 220.930 1667.090 222.110 1668.270 ;
        RECT 220.930 1665.490 222.110 1666.670 ;
        RECT 220.930 1487.090 222.110 1488.270 ;
        RECT 220.930 1485.490 222.110 1486.670 ;
        RECT 220.930 1307.090 222.110 1308.270 ;
        RECT 220.930 1305.490 222.110 1306.670 ;
        RECT 220.930 1127.090 222.110 1128.270 ;
        RECT 220.930 1125.490 222.110 1126.670 ;
        RECT 220.930 947.090 222.110 948.270 ;
        RECT 220.930 945.490 222.110 946.670 ;
        RECT 220.930 767.090 222.110 768.270 ;
        RECT 220.930 765.490 222.110 766.670 ;
        RECT 220.930 587.090 222.110 588.270 ;
        RECT 220.930 585.490 222.110 586.670 ;
        RECT 220.930 407.090 222.110 408.270 ;
        RECT 220.930 405.490 222.110 406.670 ;
        RECT 220.930 227.090 222.110 228.270 ;
        RECT 220.930 225.490 222.110 226.670 ;
        RECT 220.930 47.090 222.110 48.270 ;
        RECT 220.930 45.490 222.110 46.670 ;
        RECT 220.930 -21.310 222.110 -20.130 ;
        RECT 220.930 -22.910 222.110 -21.730 ;
        RECT 400.930 3541.410 402.110 3542.590 ;
        RECT 400.930 3539.810 402.110 3540.990 ;
        RECT 400.930 3467.090 402.110 3468.270 ;
        RECT 400.930 3465.490 402.110 3466.670 ;
        RECT 400.930 3287.090 402.110 3288.270 ;
        RECT 400.930 3285.490 402.110 3286.670 ;
        RECT 400.930 3107.090 402.110 3108.270 ;
        RECT 400.930 3105.490 402.110 3106.670 ;
        RECT 400.930 2927.090 402.110 2928.270 ;
        RECT 400.930 2925.490 402.110 2926.670 ;
        RECT 400.930 2747.090 402.110 2748.270 ;
        RECT 400.930 2745.490 402.110 2746.670 ;
        RECT 400.930 2567.090 402.110 2568.270 ;
        RECT 400.930 2565.490 402.110 2566.670 ;
        RECT 400.930 2387.090 402.110 2388.270 ;
        RECT 400.930 2385.490 402.110 2386.670 ;
        RECT 400.930 2207.090 402.110 2208.270 ;
        RECT 400.930 2205.490 402.110 2206.670 ;
        RECT 400.930 2027.090 402.110 2028.270 ;
        RECT 400.930 2025.490 402.110 2026.670 ;
        RECT 400.930 1847.090 402.110 1848.270 ;
        RECT 400.930 1845.490 402.110 1846.670 ;
        RECT 400.930 1667.090 402.110 1668.270 ;
        RECT 400.930 1665.490 402.110 1666.670 ;
        RECT 400.930 1487.090 402.110 1488.270 ;
        RECT 400.930 1485.490 402.110 1486.670 ;
        RECT 400.930 1307.090 402.110 1308.270 ;
        RECT 400.930 1305.490 402.110 1306.670 ;
        RECT 400.930 1127.090 402.110 1128.270 ;
        RECT 400.930 1125.490 402.110 1126.670 ;
        RECT 400.930 947.090 402.110 948.270 ;
        RECT 400.930 945.490 402.110 946.670 ;
        RECT 400.930 767.090 402.110 768.270 ;
        RECT 400.930 765.490 402.110 766.670 ;
        RECT 400.930 587.090 402.110 588.270 ;
        RECT 400.930 585.490 402.110 586.670 ;
        RECT 400.930 407.090 402.110 408.270 ;
        RECT 400.930 405.490 402.110 406.670 ;
        RECT 400.930 227.090 402.110 228.270 ;
        RECT 400.930 225.490 402.110 226.670 ;
        RECT 400.930 47.090 402.110 48.270 ;
        RECT 400.930 45.490 402.110 46.670 ;
        RECT 400.930 -21.310 402.110 -20.130 ;
        RECT 400.930 -22.910 402.110 -21.730 ;
        RECT 580.930 3541.410 582.110 3542.590 ;
        RECT 580.930 3539.810 582.110 3540.990 ;
        RECT 580.930 3467.090 582.110 3468.270 ;
        RECT 580.930 3465.490 582.110 3466.670 ;
        RECT 580.930 3287.090 582.110 3288.270 ;
        RECT 580.930 3285.490 582.110 3286.670 ;
        RECT 580.930 3107.090 582.110 3108.270 ;
        RECT 580.930 3105.490 582.110 3106.670 ;
        RECT 580.930 2927.090 582.110 2928.270 ;
        RECT 580.930 2925.490 582.110 2926.670 ;
        RECT 580.930 2747.090 582.110 2748.270 ;
        RECT 580.930 2745.490 582.110 2746.670 ;
        RECT 580.930 2567.090 582.110 2568.270 ;
        RECT 580.930 2565.490 582.110 2566.670 ;
        RECT 580.930 2387.090 582.110 2388.270 ;
        RECT 580.930 2385.490 582.110 2386.670 ;
        RECT 580.930 2207.090 582.110 2208.270 ;
        RECT 580.930 2205.490 582.110 2206.670 ;
        RECT 580.930 2027.090 582.110 2028.270 ;
        RECT 580.930 2025.490 582.110 2026.670 ;
        RECT 580.930 1847.090 582.110 1848.270 ;
        RECT 580.930 1845.490 582.110 1846.670 ;
        RECT 580.930 1667.090 582.110 1668.270 ;
        RECT 580.930 1665.490 582.110 1666.670 ;
        RECT 580.930 1487.090 582.110 1488.270 ;
        RECT 580.930 1485.490 582.110 1486.670 ;
        RECT 580.930 1307.090 582.110 1308.270 ;
        RECT 580.930 1305.490 582.110 1306.670 ;
        RECT 580.930 1127.090 582.110 1128.270 ;
        RECT 580.930 1125.490 582.110 1126.670 ;
        RECT 580.930 947.090 582.110 948.270 ;
        RECT 580.930 945.490 582.110 946.670 ;
        RECT 580.930 767.090 582.110 768.270 ;
        RECT 580.930 765.490 582.110 766.670 ;
        RECT 580.930 587.090 582.110 588.270 ;
        RECT 580.930 585.490 582.110 586.670 ;
        RECT 580.930 407.090 582.110 408.270 ;
        RECT 580.930 405.490 582.110 406.670 ;
        RECT 580.930 227.090 582.110 228.270 ;
        RECT 580.930 225.490 582.110 226.670 ;
        RECT 580.930 47.090 582.110 48.270 ;
        RECT 580.930 45.490 582.110 46.670 ;
        RECT 580.930 -21.310 582.110 -20.130 ;
        RECT 580.930 -22.910 582.110 -21.730 ;
        RECT 760.930 3541.410 762.110 3542.590 ;
        RECT 760.930 3539.810 762.110 3540.990 ;
        RECT 760.930 3467.090 762.110 3468.270 ;
        RECT 760.930 3465.490 762.110 3466.670 ;
        RECT 760.930 3287.090 762.110 3288.270 ;
        RECT 760.930 3285.490 762.110 3286.670 ;
        RECT 760.930 3107.090 762.110 3108.270 ;
        RECT 760.930 3105.490 762.110 3106.670 ;
        RECT 760.930 2927.090 762.110 2928.270 ;
        RECT 760.930 2925.490 762.110 2926.670 ;
        RECT 760.930 2747.090 762.110 2748.270 ;
        RECT 760.930 2745.490 762.110 2746.670 ;
        RECT 760.930 2567.090 762.110 2568.270 ;
        RECT 760.930 2565.490 762.110 2566.670 ;
        RECT 760.930 2387.090 762.110 2388.270 ;
        RECT 760.930 2385.490 762.110 2386.670 ;
        RECT 760.930 2207.090 762.110 2208.270 ;
        RECT 760.930 2205.490 762.110 2206.670 ;
        RECT 760.930 2027.090 762.110 2028.270 ;
        RECT 760.930 2025.490 762.110 2026.670 ;
        RECT 760.930 1847.090 762.110 1848.270 ;
        RECT 760.930 1845.490 762.110 1846.670 ;
        RECT 760.930 1667.090 762.110 1668.270 ;
        RECT 760.930 1665.490 762.110 1666.670 ;
        RECT 760.930 1487.090 762.110 1488.270 ;
        RECT 760.930 1485.490 762.110 1486.670 ;
        RECT 760.930 1307.090 762.110 1308.270 ;
        RECT 760.930 1305.490 762.110 1306.670 ;
        RECT 760.930 1127.090 762.110 1128.270 ;
        RECT 760.930 1125.490 762.110 1126.670 ;
        RECT 760.930 947.090 762.110 948.270 ;
        RECT 760.930 945.490 762.110 946.670 ;
        RECT 760.930 767.090 762.110 768.270 ;
        RECT 760.930 765.490 762.110 766.670 ;
        RECT 760.930 587.090 762.110 588.270 ;
        RECT 760.930 585.490 762.110 586.670 ;
        RECT 760.930 407.090 762.110 408.270 ;
        RECT 760.930 405.490 762.110 406.670 ;
        RECT 760.930 227.090 762.110 228.270 ;
        RECT 760.930 225.490 762.110 226.670 ;
        RECT 760.930 47.090 762.110 48.270 ;
        RECT 760.930 45.490 762.110 46.670 ;
        RECT 760.930 -21.310 762.110 -20.130 ;
        RECT 760.930 -22.910 762.110 -21.730 ;
        RECT 940.930 3541.410 942.110 3542.590 ;
        RECT 940.930 3539.810 942.110 3540.990 ;
        RECT 940.930 3467.090 942.110 3468.270 ;
        RECT 940.930 3465.490 942.110 3466.670 ;
        RECT 940.930 3287.090 942.110 3288.270 ;
        RECT 940.930 3285.490 942.110 3286.670 ;
        RECT 940.930 3107.090 942.110 3108.270 ;
        RECT 940.930 3105.490 942.110 3106.670 ;
        RECT 940.930 2927.090 942.110 2928.270 ;
        RECT 940.930 2925.490 942.110 2926.670 ;
        RECT 940.930 2747.090 942.110 2748.270 ;
        RECT 940.930 2745.490 942.110 2746.670 ;
        RECT 940.930 2567.090 942.110 2568.270 ;
        RECT 940.930 2565.490 942.110 2566.670 ;
        RECT 940.930 2387.090 942.110 2388.270 ;
        RECT 940.930 2385.490 942.110 2386.670 ;
        RECT 940.930 2207.090 942.110 2208.270 ;
        RECT 940.930 2205.490 942.110 2206.670 ;
        RECT 940.930 2027.090 942.110 2028.270 ;
        RECT 940.930 2025.490 942.110 2026.670 ;
        RECT 940.930 1847.090 942.110 1848.270 ;
        RECT 940.930 1845.490 942.110 1846.670 ;
        RECT 940.930 1667.090 942.110 1668.270 ;
        RECT 940.930 1665.490 942.110 1666.670 ;
        RECT 940.930 1487.090 942.110 1488.270 ;
        RECT 940.930 1485.490 942.110 1486.670 ;
        RECT 940.930 1307.090 942.110 1308.270 ;
        RECT 940.930 1305.490 942.110 1306.670 ;
        RECT 940.930 1127.090 942.110 1128.270 ;
        RECT 940.930 1125.490 942.110 1126.670 ;
        RECT 940.930 947.090 942.110 948.270 ;
        RECT 940.930 945.490 942.110 946.670 ;
        RECT 940.930 767.090 942.110 768.270 ;
        RECT 940.930 765.490 942.110 766.670 ;
        RECT 940.930 587.090 942.110 588.270 ;
        RECT 940.930 585.490 942.110 586.670 ;
        RECT 940.930 407.090 942.110 408.270 ;
        RECT 940.930 405.490 942.110 406.670 ;
        RECT 940.930 227.090 942.110 228.270 ;
        RECT 940.930 225.490 942.110 226.670 ;
        RECT 940.930 47.090 942.110 48.270 ;
        RECT 940.930 45.490 942.110 46.670 ;
        RECT 940.930 -21.310 942.110 -20.130 ;
        RECT 940.930 -22.910 942.110 -21.730 ;
        RECT 1120.930 3541.410 1122.110 3542.590 ;
        RECT 1120.930 3539.810 1122.110 3540.990 ;
        RECT 1120.930 3467.090 1122.110 3468.270 ;
        RECT 1120.930 3465.490 1122.110 3466.670 ;
        RECT 1120.930 3287.090 1122.110 3288.270 ;
        RECT 1120.930 3285.490 1122.110 3286.670 ;
        RECT 1120.930 3107.090 1122.110 3108.270 ;
        RECT 1120.930 3105.490 1122.110 3106.670 ;
        RECT 1120.930 2927.090 1122.110 2928.270 ;
        RECT 1120.930 2925.490 1122.110 2926.670 ;
        RECT 1120.930 2747.090 1122.110 2748.270 ;
        RECT 1120.930 2745.490 1122.110 2746.670 ;
        RECT 1120.930 2567.090 1122.110 2568.270 ;
        RECT 1120.930 2565.490 1122.110 2566.670 ;
        RECT 1120.930 2387.090 1122.110 2388.270 ;
        RECT 1120.930 2385.490 1122.110 2386.670 ;
        RECT 1120.930 2207.090 1122.110 2208.270 ;
        RECT 1120.930 2205.490 1122.110 2206.670 ;
        RECT 1120.930 2027.090 1122.110 2028.270 ;
        RECT 1120.930 2025.490 1122.110 2026.670 ;
        RECT 1120.930 1847.090 1122.110 1848.270 ;
        RECT 1120.930 1845.490 1122.110 1846.670 ;
        RECT 1120.930 1667.090 1122.110 1668.270 ;
        RECT 1120.930 1665.490 1122.110 1666.670 ;
        RECT 1120.930 1487.090 1122.110 1488.270 ;
        RECT 1120.930 1485.490 1122.110 1486.670 ;
        RECT 1120.930 1307.090 1122.110 1308.270 ;
        RECT 1120.930 1305.490 1122.110 1306.670 ;
        RECT 1120.930 1127.090 1122.110 1128.270 ;
        RECT 1120.930 1125.490 1122.110 1126.670 ;
        RECT 1120.930 947.090 1122.110 948.270 ;
        RECT 1120.930 945.490 1122.110 946.670 ;
        RECT 1120.930 767.090 1122.110 768.270 ;
        RECT 1120.930 765.490 1122.110 766.670 ;
        RECT 1120.930 587.090 1122.110 588.270 ;
        RECT 1120.930 585.490 1122.110 586.670 ;
        RECT 1120.930 407.090 1122.110 408.270 ;
        RECT 1120.930 405.490 1122.110 406.670 ;
        RECT 1120.930 227.090 1122.110 228.270 ;
        RECT 1120.930 225.490 1122.110 226.670 ;
        RECT 1120.930 47.090 1122.110 48.270 ;
        RECT 1120.930 45.490 1122.110 46.670 ;
        RECT 1120.930 -21.310 1122.110 -20.130 ;
        RECT 1120.930 -22.910 1122.110 -21.730 ;
        RECT 1300.930 3541.410 1302.110 3542.590 ;
        RECT 1300.930 3539.810 1302.110 3540.990 ;
        RECT 1300.930 3467.090 1302.110 3468.270 ;
        RECT 1300.930 3465.490 1302.110 3466.670 ;
        RECT 1300.930 3287.090 1302.110 3288.270 ;
        RECT 1300.930 3285.490 1302.110 3286.670 ;
        RECT 1300.930 3107.090 1302.110 3108.270 ;
        RECT 1300.930 3105.490 1302.110 3106.670 ;
        RECT 1300.930 2927.090 1302.110 2928.270 ;
        RECT 1300.930 2925.490 1302.110 2926.670 ;
        RECT 1300.930 2747.090 1302.110 2748.270 ;
        RECT 1300.930 2745.490 1302.110 2746.670 ;
        RECT 1300.930 2567.090 1302.110 2568.270 ;
        RECT 1300.930 2565.490 1302.110 2566.670 ;
        RECT 1300.930 2387.090 1302.110 2388.270 ;
        RECT 1300.930 2385.490 1302.110 2386.670 ;
        RECT 1300.930 2207.090 1302.110 2208.270 ;
        RECT 1300.930 2205.490 1302.110 2206.670 ;
        RECT 1300.930 2027.090 1302.110 2028.270 ;
        RECT 1300.930 2025.490 1302.110 2026.670 ;
        RECT 1300.930 1847.090 1302.110 1848.270 ;
        RECT 1300.930 1845.490 1302.110 1846.670 ;
        RECT 1300.930 1667.090 1302.110 1668.270 ;
        RECT 1300.930 1665.490 1302.110 1666.670 ;
        RECT 1300.930 1487.090 1302.110 1488.270 ;
        RECT 1300.930 1485.490 1302.110 1486.670 ;
        RECT 1300.930 1307.090 1302.110 1308.270 ;
        RECT 1300.930 1305.490 1302.110 1306.670 ;
        RECT 1300.930 1127.090 1302.110 1128.270 ;
        RECT 1300.930 1125.490 1302.110 1126.670 ;
        RECT 1300.930 947.090 1302.110 948.270 ;
        RECT 1300.930 945.490 1302.110 946.670 ;
        RECT 1300.930 767.090 1302.110 768.270 ;
        RECT 1300.930 765.490 1302.110 766.670 ;
        RECT 1300.930 587.090 1302.110 588.270 ;
        RECT 1300.930 585.490 1302.110 586.670 ;
        RECT 1300.930 407.090 1302.110 408.270 ;
        RECT 1300.930 405.490 1302.110 406.670 ;
        RECT 1300.930 227.090 1302.110 228.270 ;
        RECT 1300.930 225.490 1302.110 226.670 ;
        RECT 1300.930 47.090 1302.110 48.270 ;
        RECT 1300.930 45.490 1302.110 46.670 ;
        RECT 1300.930 -21.310 1302.110 -20.130 ;
        RECT 1300.930 -22.910 1302.110 -21.730 ;
        RECT 1480.930 3541.410 1482.110 3542.590 ;
        RECT 1480.930 3539.810 1482.110 3540.990 ;
        RECT 1480.930 3467.090 1482.110 3468.270 ;
        RECT 1480.930 3465.490 1482.110 3466.670 ;
        RECT 1480.930 3287.090 1482.110 3288.270 ;
        RECT 1480.930 3285.490 1482.110 3286.670 ;
        RECT 1480.930 3107.090 1482.110 3108.270 ;
        RECT 1480.930 3105.490 1482.110 3106.670 ;
        RECT 1480.930 2927.090 1482.110 2928.270 ;
        RECT 1480.930 2925.490 1482.110 2926.670 ;
        RECT 1480.930 2747.090 1482.110 2748.270 ;
        RECT 1480.930 2745.490 1482.110 2746.670 ;
        RECT 1480.930 2567.090 1482.110 2568.270 ;
        RECT 1480.930 2565.490 1482.110 2566.670 ;
        RECT 1480.930 2387.090 1482.110 2388.270 ;
        RECT 1480.930 2385.490 1482.110 2386.670 ;
        RECT 1480.930 2207.090 1482.110 2208.270 ;
        RECT 1480.930 2205.490 1482.110 2206.670 ;
        RECT 1480.930 2027.090 1482.110 2028.270 ;
        RECT 1480.930 2025.490 1482.110 2026.670 ;
        RECT 1480.930 1847.090 1482.110 1848.270 ;
        RECT 1480.930 1845.490 1482.110 1846.670 ;
        RECT 1480.930 1667.090 1482.110 1668.270 ;
        RECT 1480.930 1665.490 1482.110 1666.670 ;
        RECT 1480.930 1487.090 1482.110 1488.270 ;
        RECT 1480.930 1485.490 1482.110 1486.670 ;
        RECT 1480.930 1307.090 1482.110 1308.270 ;
        RECT 1480.930 1305.490 1482.110 1306.670 ;
        RECT 1480.930 1127.090 1482.110 1128.270 ;
        RECT 1480.930 1125.490 1482.110 1126.670 ;
        RECT 1480.930 947.090 1482.110 948.270 ;
        RECT 1480.930 945.490 1482.110 946.670 ;
        RECT 1480.930 767.090 1482.110 768.270 ;
        RECT 1480.930 765.490 1482.110 766.670 ;
        RECT 1480.930 587.090 1482.110 588.270 ;
        RECT 1480.930 585.490 1482.110 586.670 ;
        RECT 1480.930 407.090 1482.110 408.270 ;
        RECT 1480.930 405.490 1482.110 406.670 ;
        RECT 1480.930 227.090 1482.110 228.270 ;
        RECT 1480.930 225.490 1482.110 226.670 ;
        RECT 1480.930 47.090 1482.110 48.270 ;
        RECT 1480.930 45.490 1482.110 46.670 ;
        RECT 1480.930 -21.310 1482.110 -20.130 ;
        RECT 1480.930 -22.910 1482.110 -21.730 ;
        RECT 1660.930 3541.410 1662.110 3542.590 ;
        RECT 1660.930 3539.810 1662.110 3540.990 ;
        RECT 1660.930 3467.090 1662.110 3468.270 ;
        RECT 1660.930 3465.490 1662.110 3466.670 ;
        RECT 1660.930 3287.090 1662.110 3288.270 ;
        RECT 1660.930 3285.490 1662.110 3286.670 ;
        RECT 1660.930 3107.090 1662.110 3108.270 ;
        RECT 1660.930 3105.490 1662.110 3106.670 ;
        RECT 1660.930 2927.090 1662.110 2928.270 ;
        RECT 1660.930 2925.490 1662.110 2926.670 ;
        RECT 1660.930 2747.090 1662.110 2748.270 ;
        RECT 1660.930 2745.490 1662.110 2746.670 ;
        RECT 1660.930 2567.090 1662.110 2568.270 ;
        RECT 1660.930 2565.490 1662.110 2566.670 ;
        RECT 1660.930 2387.090 1662.110 2388.270 ;
        RECT 1660.930 2385.490 1662.110 2386.670 ;
        RECT 1660.930 2207.090 1662.110 2208.270 ;
        RECT 1660.930 2205.490 1662.110 2206.670 ;
        RECT 1660.930 2027.090 1662.110 2028.270 ;
        RECT 1660.930 2025.490 1662.110 2026.670 ;
        RECT 1660.930 1847.090 1662.110 1848.270 ;
        RECT 1660.930 1845.490 1662.110 1846.670 ;
        RECT 1660.930 1667.090 1662.110 1668.270 ;
        RECT 1660.930 1665.490 1662.110 1666.670 ;
        RECT 1660.930 1487.090 1662.110 1488.270 ;
        RECT 1660.930 1485.490 1662.110 1486.670 ;
        RECT 1660.930 1307.090 1662.110 1308.270 ;
        RECT 1660.930 1305.490 1662.110 1306.670 ;
        RECT 1660.930 1127.090 1662.110 1128.270 ;
        RECT 1660.930 1125.490 1662.110 1126.670 ;
        RECT 1660.930 947.090 1662.110 948.270 ;
        RECT 1660.930 945.490 1662.110 946.670 ;
        RECT 1660.930 767.090 1662.110 768.270 ;
        RECT 1660.930 765.490 1662.110 766.670 ;
        RECT 1660.930 587.090 1662.110 588.270 ;
        RECT 1660.930 585.490 1662.110 586.670 ;
        RECT 1660.930 407.090 1662.110 408.270 ;
        RECT 1660.930 405.490 1662.110 406.670 ;
        RECT 1660.930 227.090 1662.110 228.270 ;
        RECT 1660.930 225.490 1662.110 226.670 ;
        RECT 1660.930 47.090 1662.110 48.270 ;
        RECT 1660.930 45.490 1662.110 46.670 ;
        RECT 1660.930 -21.310 1662.110 -20.130 ;
        RECT 1660.930 -22.910 1662.110 -21.730 ;
        RECT 1840.930 3541.410 1842.110 3542.590 ;
        RECT 1840.930 3539.810 1842.110 3540.990 ;
        RECT 1840.930 3467.090 1842.110 3468.270 ;
        RECT 1840.930 3465.490 1842.110 3466.670 ;
        RECT 1840.930 3287.090 1842.110 3288.270 ;
        RECT 1840.930 3285.490 1842.110 3286.670 ;
        RECT 1840.930 3107.090 1842.110 3108.270 ;
        RECT 1840.930 3105.490 1842.110 3106.670 ;
        RECT 1840.930 2927.090 1842.110 2928.270 ;
        RECT 1840.930 2925.490 1842.110 2926.670 ;
        RECT 1840.930 2747.090 1842.110 2748.270 ;
        RECT 1840.930 2745.490 1842.110 2746.670 ;
        RECT 1840.930 2567.090 1842.110 2568.270 ;
        RECT 1840.930 2565.490 1842.110 2566.670 ;
        RECT 1840.930 2387.090 1842.110 2388.270 ;
        RECT 1840.930 2385.490 1842.110 2386.670 ;
        RECT 1840.930 2207.090 1842.110 2208.270 ;
        RECT 1840.930 2205.490 1842.110 2206.670 ;
        RECT 1840.930 2027.090 1842.110 2028.270 ;
        RECT 1840.930 2025.490 1842.110 2026.670 ;
        RECT 1840.930 1847.090 1842.110 1848.270 ;
        RECT 1840.930 1845.490 1842.110 1846.670 ;
        RECT 1840.930 1667.090 1842.110 1668.270 ;
        RECT 1840.930 1665.490 1842.110 1666.670 ;
        RECT 1840.930 1487.090 1842.110 1488.270 ;
        RECT 1840.930 1485.490 1842.110 1486.670 ;
        RECT 1840.930 1307.090 1842.110 1308.270 ;
        RECT 1840.930 1305.490 1842.110 1306.670 ;
        RECT 1840.930 1127.090 1842.110 1128.270 ;
        RECT 1840.930 1125.490 1842.110 1126.670 ;
        RECT 1840.930 947.090 1842.110 948.270 ;
        RECT 1840.930 945.490 1842.110 946.670 ;
        RECT 1840.930 767.090 1842.110 768.270 ;
        RECT 1840.930 765.490 1842.110 766.670 ;
        RECT 1840.930 587.090 1842.110 588.270 ;
        RECT 1840.930 585.490 1842.110 586.670 ;
        RECT 1840.930 407.090 1842.110 408.270 ;
        RECT 1840.930 405.490 1842.110 406.670 ;
        RECT 1840.930 227.090 1842.110 228.270 ;
        RECT 1840.930 225.490 1842.110 226.670 ;
        RECT 1840.930 47.090 1842.110 48.270 ;
        RECT 1840.930 45.490 1842.110 46.670 ;
        RECT 1840.930 -21.310 1842.110 -20.130 ;
        RECT 1840.930 -22.910 1842.110 -21.730 ;
        RECT 2020.930 3541.410 2022.110 3542.590 ;
        RECT 2020.930 3539.810 2022.110 3540.990 ;
        RECT 2020.930 3467.090 2022.110 3468.270 ;
        RECT 2020.930 3465.490 2022.110 3466.670 ;
        RECT 2020.930 3287.090 2022.110 3288.270 ;
        RECT 2020.930 3285.490 2022.110 3286.670 ;
        RECT 2020.930 3107.090 2022.110 3108.270 ;
        RECT 2020.930 3105.490 2022.110 3106.670 ;
        RECT 2020.930 2927.090 2022.110 2928.270 ;
        RECT 2020.930 2925.490 2022.110 2926.670 ;
        RECT 2020.930 2747.090 2022.110 2748.270 ;
        RECT 2020.930 2745.490 2022.110 2746.670 ;
        RECT 2020.930 2567.090 2022.110 2568.270 ;
        RECT 2020.930 2565.490 2022.110 2566.670 ;
        RECT 2020.930 2387.090 2022.110 2388.270 ;
        RECT 2020.930 2385.490 2022.110 2386.670 ;
        RECT 2020.930 2207.090 2022.110 2208.270 ;
        RECT 2020.930 2205.490 2022.110 2206.670 ;
        RECT 2020.930 2027.090 2022.110 2028.270 ;
        RECT 2020.930 2025.490 2022.110 2026.670 ;
        RECT 2020.930 1847.090 2022.110 1848.270 ;
        RECT 2020.930 1845.490 2022.110 1846.670 ;
        RECT 2020.930 1667.090 2022.110 1668.270 ;
        RECT 2020.930 1665.490 2022.110 1666.670 ;
        RECT 2020.930 1487.090 2022.110 1488.270 ;
        RECT 2020.930 1485.490 2022.110 1486.670 ;
        RECT 2020.930 1307.090 2022.110 1308.270 ;
        RECT 2020.930 1305.490 2022.110 1306.670 ;
        RECT 2020.930 1127.090 2022.110 1128.270 ;
        RECT 2020.930 1125.490 2022.110 1126.670 ;
        RECT 2020.930 947.090 2022.110 948.270 ;
        RECT 2020.930 945.490 2022.110 946.670 ;
        RECT 2020.930 767.090 2022.110 768.270 ;
        RECT 2020.930 765.490 2022.110 766.670 ;
        RECT 2020.930 587.090 2022.110 588.270 ;
        RECT 2020.930 585.490 2022.110 586.670 ;
        RECT 2020.930 407.090 2022.110 408.270 ;
        RECT 2020.930 405.490 2022.110 406.670 ;
        RECT 2020.930 227.090 2022.110 228.270 ;
        RECT 2020.930 225.490 2022.110 226.670 ;
        RECT 2020.930 47.090 2022.110 48.270 ;
        RECT 2020.930 45.490 2022.110 46.670 ;
        RECT 2020.930 -21.310 2022.110 -20.130 ;
        RECT 2020.930 -22.910 2022.110 -21.730 ;
        RECT 2200.930 3541.410 2202.110 3542.590 ;
        RECT 2200.930 3539.810 2202.110 3540.990 ;
        RECT 2200.930 3467.090 2202.110 3468.270 ;
        RECT 2200.930 3465.490 2202.110 3466.670 ;
        RECT 2200.930 3287.090 2202.110 3288.270 ;
        RECT 2200.930 3285.490 2202.110 3286.670 ;
        RECT 2200.930 3107.090 2202.110 3108.270 ;
        RECT 2200.930 3105.490 2202.110 3106.670 ;
        RECT 2200.930 2927.090 2202.110 2928.270 ;
        RECT 2200.930 2925.490 2202.110 2926.670 ;
        RECT 2200.930 2747.090 2202.110 2748.270 ;
        RECT 2200.930 2745.490 2202.110 2746.670 ;
        RECT 2200.930 2567.090 2202.110 2568.270 ;
        RECT 2200.930 2565.490 2202.110 2566.670 ;
        RECT 2200.930 2387.090 2202.110 2388.270 ;
        RECT 2200.930 2385.490 2202.110 2386.670 ;
        RECT 2200.930 2207.090 2202.110 2208.270 ;
        RECT 2200.930 2205.490 2202.110 2206.670 ;
        RECT 2200.930 2027.090 2202.110 2028.270 ;
        RECT 2200.930 2025.490 2202.110 2026.670 ;
        RECT 2200.930 1847.090 2202.110 1848.270 ;
        RECT 2200.930 1845.490 2202.110 1846.670 ;
        RECT 2200.930 1667.090 2202.110 1668.270 ;
        RECT 2200.930 1665.490 2202.110 1666.670 ;
        RECT 2200.930 1487.090 2202.110 1488.270 ;
        RECT 2200.930 1485.490 2202.110 1486.670 ;
        RECT 2200.930 1307.090 2202.110 1308.270 ;
        RECT 2200.930 1305.490 2202.110 1306.670 ;
        RECT 2200.930 1127.090 2202.110 1128.270 ;
        RECT 2200.930 1125.490 2202.110 1126.670 ;
        RECT 2200.930 947.090 2202.110 948.270 ;
        RECT 2200.930 945.490 2202.110 946.670 ;
        RECT 2200.930 767.090 2202.110 768.270 ;
        RECT 2200.930 765.490 2202.110 766.670 ;
        RECT 2200.930 587.090 2202.110 588.270 ;
        RECT 2200.930 585.490 2202.110 586.670 ;
        RECT 2200.930 407.090 2202.110 408.270 ;
        RECT 2200.930 405.490 2202.110 406.670 ;
        RECT 2200.930 227.090 2202.110 228.270 ;
        RECT 2200.930 225.490 2202.110 226.670 ;
        RECT 2200.930 47.090 2202.110 48.270 ;
        RECT 2200.930 45.490 2202.110 46.670 ;
        RECT 2200.930 -21.310 2202.110 -20.130 ;
        RECT 2200.930 -22.910 2202.110 -21.730 ;
        RECT 2380.930 3541.410 2382.110 3542.590 ;
        RECT 2380.930 3539.810 2382.110 3540.990 ;
        RECT 2380.930 3467.090 2382.110 3468.270 ;
        RECT 2380.930 3465.490 2382.110 3466.670 ;
        RECT 2380.930 3287.090 2382.110 3288.270 ;
        RECT 2380.930 3285.490 2382.110 3286.670 ;
        RECT 2380.930 3107.090 2382.110 3108.270 ;
        RECT 2380.930 3105.490 2382.110 3106.670 ;
        RECT 2380.930 2927.090 2382.110 2928.270 ;
        RECT 2380.930 2925.490 2382.110 2926.670 ;
        RECT 2380.930 2747.090 2382.110 2748.270 ;
        RECT 2380.930 2745.490 2382.110 2746.670 ;
        RECT 2380.930 2567.090 2382.110 2568.270 ;
        RECT 2380.930 2565.490 2382.110 2566.670 ;
        RECT 2380.930 2387.090 2382.110 2388.270 ;
        RECT 2380.930 2385.490 2382.110 2386.670 ;
        RECT 2380.930 2207.090 2382.110 2208.270 ;
        RECT 2380.930 2205.490 2382.110 2206.670 ;
        RECT 2380.930 2027.090 2382.110 2028.270 ;
        RECT 2380.930 2025.490 2382.110 2026.670 ;
        RECT 2380.930 1847.090 2382.110 1848.270 ;
        RECT 2380.930 1845.490 2382.110 1846.670 ;
        RECT 2380.930 1667.090 2382.110 1668.270 ;
        RECT 2380.930 1665.490 2382.110 1666.670 ;
        RECT 2380.930 1487.090 2382.110 1488.270 ;
        RECT 2380.930 1485.490 2382.110 1486.670 ;
        RECT 2380.930 1307.090 2382.110 1308.270 ;
        RECT 2380.930 1305.490 2382.110 1306.670 ;
        RECT 2380.930 1127.090 2382.110 1128.270 ;
        RECT 2380.930 1125.490 2382.110 1126.670 ;
        RECT 2380.930 947.090 2382.110 948.270 ;
        RECT 2380.930 945.490 2382.110 946.670 ;
        RECT 2380.930 767.090 2382.110 768.270 ;
        RECT 2380.930 765.490 2382.110 766.670 ;
        RECT 2380.930 587.090 2382.110 588.270 ;
        RECT 2380.930 585.490 2382.110 586.670 ;
        RECT 2380.930 407.090 2382.110 408.270 ;
        RECT 2380.930 405.490 2382.110 406.670 ;
        RECT 2380.930 227.090 2382.110 228.270 ;
        RECT 2380.930 225.490 2382.110 226.670 ;
        RECT 2380.930 47.090 2382.110 48.270 ;
        RECT 2380.930 45.490 2382.110 46.670 ;
        RECT 2380.930 -21.310 2382.110 -20.130 ;
        RECT 2380.930 -22.910 2382.110 -21.730 ;
        RECT 2560.930 3541.410 2562.110 3542.590 ;
        RECT 2560.930 3539.810 2562.110 3540.990 ;
        RECT 2560.930 3467.090 2562.110 3468.270 ;
        RECT 2560.930 3465.490 2562.110 3466.670 ;
        RECT 2560.930 3287.090 2562.110 3288.270 ;
        RECT 2560.930 3285.490 2562.110 3286.670 ;
        RECT 2560.930 3107.090 2562.110 3108.270 ;
        RECT 2560.930 3105.490 2562.110 3106.670 ;
        RECT 2560.930 2927.090 2562.110 2928.270 ;
        RECT 2560.930 2925.490 2562.110 2926.670 ;
        RECT 2560.930 2747.090 2562.110 2748.270 ;
        RECT 2560.930 2745.490 2562.110 2746.670 ;
        RECT 2560.930 2567.090 2562.110 2568.270 ;
        RECT 2560.930 2565.490 2562.110 2566.670 ;
        RECT 2560.930 2387.090 2562.110 2388.270 ;
        RECT 2560.930 2385.490 2562.110 2386.670 ;
        RECT 2560.930 2207.090 2562.110 2208.270 ;
        RECT 2560.930 2205.490 2562.110 2206.670 ;
        RECT 2560.930 2027.090 2562.110 2028.270 ;
        RECT 2560.930 2025.490 2562.110 2026.670 ;
        RECT 2560.930 1847.090 2562.110 1848.270 ;
        RECT 2560.930 1845.490 2562.110 1846.670 ;
        RECT 2560.930 1667.090 2562.110 1668.270 ;
        RECT 2560.930 1665.490 2562.110 1666.670 ;
        RECT 2560.930 1487.090 2562.110 1488.270 ;
        RECT 2560.930 1485.490 2562.110 1486.670 ;
        RECT 2560.930 1307.090 2562.110 1308.270 ;
        RECT 2560.930 1305.490 2562.110 1306.670 ;
        RECT 2560.930 1127.090 2562.110 1128.270 ;
        RECT 2560.930 1125.490 2562.110 1126.670 ;
        RECT 2560.930 947.090 2562.110 948.270 ;
        RECT 2560.930 945.490 2562.110 946.670 ;
        RECT 2560.930 767.090 2562.110 768.270 ;
        RECT 2560.930 765.490 2562.110 766.670 ;
        RECT 2560.930 587.090 2562.110 588.270 ;
        RECT 2560.930 585.490 2562.110 586.670 ;
        RECT 2560.930 407.090 2562.110 408.270 ;
        RECT 2560.930 405.490 2562.110 406.670 ;
        RECT 2560.930 227.090 2562.110 228.270 ;
        RECT 2560.930 225.490 2562.110 226.670 ;
        RECT 2560.930 47.090 2562.110 48.270 ;
        RECT 2560.930 45.490 2562.110 46.670 ;
        RECT 2560.930 -21.310 2562.110 -20.130 ;
        RECT 2560.930 -22.910 2562.110 -21.730 ;
        RECT 2740.930 3541.410 2742.110 3542.590 ;
        RECT 2740.930 3539.810 2742.110 3540.990 ;
        RECT 2740.930 3467.090 2742.110 3468.270 ;
        RECT 2740.930 3465.490 2742.110 3466.670 ;
        RECT 2740.930 3287.090 2742.110 3288.270 ;
        RECT 2740.930 3285.490 2742.110 3286.670 ;
        RECT 2740.930 3107.090 2742.110 3108.270 ;
        RECT 2740.930 3105.490 2742.110 3106.670 ;
        RECT 2740.930 2927.090 2742.110 2928.270 ;
        RECT 2740.930 2925.490 2742.110 2926.670 ;
        RECT 2740.930 2747.090 2742.110 2748.270 ;
        RECT 2740.930 2745.490 2742.110 2746.670 ;
        RECT 2740.930 2567.090 2742.110 2568.270 ;
        RECT 2740.930 2565.490 2742.110 2566.670 ;
        RECT 2740.930 2387.090 2742.110 2388.270 ;
        RECT 2740.930 2385.490 2742.110 2386.670 ;
        RECT 2740.930 2207.090 2742.110 2208.270 ;
        RECT 2740.930 2205.490 2742.110 2206.670 ;
        RECT 2740.930 2027.090 2742.110 2028.270 ;
        RECT 2740.930 2025.490 2742.110 2026.670 ;
        RECT 2740.930 1847.090 2742.110 1848.270 ;
        RECT 2740.930 1845.490 2742.110 1846.670 ;
        RECT 2740.930 1667.090 2742.110 1668.270 ;
        RECT 2740.930 1665.490 2742.110 1666.670 ;
        RECT 2740.930 1487.090 2742.110 1488.270 ;
        RECT 2740.930 1485.490 2742.110 1486.670 ;
        RECT 2740.930 1307.090 2742.110 1308.270 ;
        RECT 2740.930 1305.490 2742.110 1306.670 ;
        RECT 2740.930 1127.090 2742.110 1128.270 ;
        RECT 2740.930 1125.490 2742.110 1126.670 ;
        RECT 2740.930 947.090 2742.110 948.270 ;
        RECT 2740.930 945.490 2742.110 946.670 ;
        RECT 2740.930 767.090 2742.110 768.270 ;
        RECT 2740.930 765.490 2742.110 766.670 ;
        RECT 2740.930 587.090 2742.110 588.270 ;
        RECT 2740.930 585.490 2742.110 586.670 ;
        RECT 2740.930 407.090 2742.110 408.270 ;
        RECT 2740.930 405.490 2742.110 406.670 ;
        RECT 2740.930 227.090 2742.110 228.270 ;
        RECT 2740.930 225.490 2742.110 226.670 ;
        RECT 2740.930 47.090 2742.110 48.270 ;
        RECT 2740.930 45.490 2742.110 46.670 ;
        RECT 2740.930 -21.310 2742.110 -20.130 ;
        RECT 2740.930 -22.910 2742.110 -21.730 ;
        RECT 2945.910 3541.410 2947.090 3542.590 ;
        RECT 2945.910 3539.810 2947.090 3540.990 ;
        RECT 2945.910 3467.090 2947.090 3468.270 ;
        RECT 2945.910 3465.490 2947.090 3466.670 ;
        RECT 2945.910 3287.090 2947.090 3288.270 ;
        RECT 2945.910 3285.490 2947.090 3286.670 ;
        RECT 2945.910 3107.090 2947.090 3108.270 ;
        RECT 2945.910 3105.490 2947.090 3106.670 ;
        RECT 2945.910 2927.090 2947.090 2928.270 ;
        RECT 2945.910 2925.490 2947.090 2926.670 ;
        RECT 2945.910 2747.090 2947.090 2748.270 ;
        RECT 2945.910 2745.490 2947.090 2746.670 ;
        RECT 2945.910 2567.090 2947.090 2568.270 ;
        RECT 2945.910 2565.490 2947.090 2566.670 ;
        RECT 2945.910 2387.090 2947.090 2388.270 ;
        RECT 2945.910 2385.490 2947.090 2386.670 ;
        RECT 2945.910 2207.090 2947.090 2208.270 ;
        RECT 2945.910 2205.490 2947.090 2206.670 ;
        RECT 2945.910 2027.090 2947.090 2028.270 ;
        RECT 2945.910 2025.490 2947.090 2026.670 ;
        RECT 2945.910 1847.090 2947.090 1848.270 ;
        RECT 2945.910 1845.490 2947.090 1846.670 ;
        RECT 2945.910 1667.090 2947.090 1668.270 ;
        RECT 2945.910 1665.490 2947.090 1666.670 ;
        RECT 2945.910 1487.090 2947.090 1488.270 ;
        RECT 2945.910 1485.490 2947.090 1486.670 ;
        RECT 2945.910 1307.090 2947.090 1308.270 ;
        RECT 2945.910 1305.490 2947.090 1306.670 ;
        RECT 2945.910 1127.090 2947.090 1128.270 ;
        RECT 2945.910 1125.490 2947.090 1126.670 ;
        RECT 2945.910 947.090 2947.090 948.270 ;
        RECT 2945.910 945.490 2947.090 946.670 ;
        RECT 2945.910 767.090 2947.090 768.270 ;
        RECT 2945.910 765.490 2947.090 766.670 ;
        RECT 2945.910 587.090 2947.090 588.270 ;
        RECT 2945.910 585.490 2947.090 586.670 ;
        RECT 2945.910 407.090 2947.090 408.270 ;
        RECT 2945.910 405.490 2947.090 406.670 ;
        RECT 2945.910 227.090 2947.090 228.270 ;
        RECT 2945.910 225.490 2947.090 226.670 ;
        RECT 2945.910 47.090 2947.090 48.270 ;
        RECT 2945.910 45.490 2947.090 46.670 ;
        RECT 2945.910 -21.310 2947.090 -20.130 ;
        RECT 2945.910 -22.910 2947.090 -21.730 ;
      LAYER met5 ;
        RECT -28.380 3542.700 -25.380 3542.710 ;
        RECT 40.020 3542.700 43.020 3542.710 ;
        RECT 220.020 3542.700 223.020 3542.710 ;
        RECT 400.020 3542.700 403.020 3542.710 ;
        RECT 580.020 3542.700 583.020 3542.710 ;
        RECT 760.020 3542.700 763.020 3542.710 ;
        RECT 940.020 3542.700 943.020 3542.710 ;
        RECT 1120.020 3542.700 1123.020 3542.710 ;
        RECT 1300.020 3542.700 1303.020 3542.710 ;
        RECT 1480.020 3542.700 1483.020 3542.710 ;
        RECT 1660.020 3542.700 1663.020 3542.710 ;
        RECT 1840.020 3542.700 1843.020 3542.710 ;
        RECT 2020.020 3542.700 2023.020 3542.710 ;
        RECT 2200.020 3542.700 2203.020 3542.710 ;
        RECT 2380.020 3542.700 2383.020 3542.710 ;
        RECT 2560.020 3542.700 2563.020 3542.710 ;
        RECT 2740.020 3542.700 2743.020 3542.710 ;
        RECT 2945.000 3542.700 2948.000 3542.710 ;
        RECT -28.380 3539.700 2948.000 3542.700 ;
        RECT -28.380 3539.690 -25.380 3539.700 ;
        RECT 40.020 3539.690 43.020 3539.700 ;
        RECT 220.020 3539.690 223.020 3539.700 ;
        RECT 400.020 3539.690 403.020 3539.700 ;
        RECT 580.020 3539.690 583.020 3539.700 ;
        RECT 760.020 3539.690 763.020 3539.700 ;
        RECT 940.020 3539.690 943.020 3539.700 ;
        RECT 1120.020 3539.690 1123.020 3539.700 ;
        RECT 1300.020 3539.690 1303.020 3539.700 ;
        RECT 1480.020 3539.690 1483.020 3539.700 ;
        RECT 1660.020 3539.690 1663.020 3539.700 ;
        RECT 1840.020 3539.690 1843.020 3539.700 ;
        RECT 2020.020 3539.690 2023.020 3539.700 ;
        RECT 2200.020 3539.690 2203.020 3539.700 ;
        RECT 2380.020 3539.690 2383.020 3539.700 ;
        RECT 2560.020 3539.690 2563.020 3539.700 ;
        RECT 2740.020 3539.690 2743.020 3539.700 ;
        RECT 2945.000 3539.690 2948.000 3539.700 ;
        RECT -28.380 3468.380 -25.380 3468.390 ;
        RECT 40.020 3468.380 43.020 3468.390 ;
        RECT 220.020 3468.380 223.020 3468.390 ;
        RECT 400.020 3468.380 403.020 3468.390 ;
        RECT 580.020 3468.380 583.020 3468.390 ;
        RECT 760.020 3468.380 763.020 3468.390 ;
        RECT 940.020 3468.380 943.020 3468.390 ;
        RECT 1120.020 3468.380 1123.020 3468.390 ;
        RECT 1300.020 3468.380 1303.020 3468.390 ;
        RECT 1480.020 3468.380 1483.020 3468.390 ;
        RECT 1660.020 3468.380 1663.020 3468.390 ;
        RECT 1840.020 3468.380 1843.020 3468.390 ;
        RECT 2020.020 3468.380 2023.020 3468.390 ;
        RECT 2200.020 3468.380 2203.020 3468.390 ;
        RECT 2380.020 3468.380 2383.020 3468.390 ;
        RECT 2560.020 3468.380 2563.020 3468.390 ;
        RECT 2740.020 3468.380 2743.020 3468.390 ;
        RECT 2945.000 3468.380 2948.000 3468.390 ;
        RECT -32.980 3465.380 2952.600 3468.380 ;
        RECT -28.380 3465.370 -25.380 3465.380 ;
        RECT 40.020 3465.370 43.020 3465.380 ;
        RECT 220.020 3465.370 223.020 3465.380 ;
        RECT 400.020 3465.370 403.020 3465.380 ;
        RECT 580.020 3465.370 583.020 3465.380 ;
        RECT 760.020 3465.370 763.020 3465.380 ;
        RECT 940.020 3465.370 943.020 3465.380 ;
        RECT 1120.020 3465.370 1123.020 3465.380 ;
        RECT 1300.020 3465.370 1303.020 3465.380 ;
        RECT 1480.020 3465.370 1483.020 3465.380 ;
        RECT 1660.020 3465.370 1663.020 3465.380 ;
        RECT 1840.020 3465.370 1843.020 3465.380 ;
        RECT 2020.020 3465.370 2023.020 3465.380 ;
        RECT 2200.020 3465.370 2203.020 3465.380 ;
        RECT 2380.020 3465.370 2383.020 3465.380 ;
        RECT 2560.020 3465.370 2563.020 3465.380 ;
        RECT 2740.020 3465.370 2743.020 3465.380 ;
        RECT 2945.000 3465.370 2948.000 3465.380 ;
        RECT -28.380 3288.380 -25.380 3288.390 ;
        RECT 40.020 3288.380 43.020 3288.390 ;
        RECT 220.020 3288.380 223.020 3288.390 ;
        RECT 400.020 3288.380 403.020 3288.390 ;
        RECT 580.020 3288.380 583.020 3288.390 ;
        RECT 760.020 3288.380 763.020 3288.390 ;
        RECT 940.020 3288.380 943.020 3288.390 ;
        RECT 1120.020 3288.380 1123.020 3288.390 ;
        RECT 1300.020 3288.380 1303.020 3288.390 ;
        RECT 1480.020 3288.380 1483.020 3288.390 ;
        RECT 1660.020 3288.380 1663.020 3288.390 ;
        RECT 1840.020 3288.380 1843.020 3288.390 ;
        RECT 2020.020 3288.380 2023.020 3288.390 ;
        RECT 2200.020 3288.380 2203.020 3288.390 ;
        RECT 2380.020 3288.380 2383.020 3288.390 ;
        RECT 2560.020 3288.380 2563.020 3288.390 ;
        RECT 2740.020 3288.380 2743.020 3288.390 ;
        RECT 2945.000 3288.380 2948.000 3288.390 ;
        RECT -32.980 3285.380 2952.600 3288.380 ;
        RECT -28.380 3285.370 -25.380 3285.380 ;
        RECT 40.020 3285.370 43.020 3285.380 ;
        RECT 220.020 3285.370 223.020 3285.380 ;
        RECT 400.020 3285.370 403.020 3285.380 ;
        RECT 580.020 3285.370 583.020 3285.380 ;
        RECT 760.020 3285.370 763.020 3285.380 ;
        RECT 940.020 3285.370 943.020 3285.380 ;
        RECT 1120.020 3285.370 1123.020 3285.380 ;
        RECT 1300.020 3285.370 1303.020 3285.380 ;
        RECT 1480.020 3285.370 1483.020 3285.380 ;
        RECT 1660.020 3285.370 1663.020 3285.380 ;
        RECT 1840.020 3285.370 1843.020 3285.380 ;
        RECT 2020.020 3285.370 2023.020 3285.380 ;
        RECT 2200.020 3285.370 2203.020 3285.380 ;
        RECT 2380.020 3285.370 2383.020 3285.380 ;
        RECT 2560.020 3285.370 2563.020 3285.380 ;
        RECT 2740.020 3285.370 2743.020 3285.380 ;
        RECT 2945.000 3285.370 2948.000 3285.380 ;
        RECT -28.380 3108.380 -25.380 3108.390 ;
        RECT 40.020 3108.380 43.020 3108.390 ;
        RECT 220.020 3108.380 223.020 3108.390 ;
        RECT 400.020 3108.380 403.020 3108.390 ;
        RECT 580.020 3108.380 583.020 3108.390 ;
        RECT 760.020 3108.380 763.020 3108.390 ;
        RECT 940.020 3108.380 943.020 3108.390 ;
        RECT 1120.020 3108.380 1123.020 3108.390 ;
        RECT 1300.020 3108.380 1303.020 3108.390 ;
        RECT 1480.020 3108.380 1483.020 3108.390 ;
        RECT 1660.020 3108.380 1663.020 3108.390 ;
        RECT 1840.020 3108.380 1843.020 3108.390 ;
        RECT 2020.020 3108.380 2023.020 3108.390 ;
        RECT 2200.020 3108.380 2203.020 3108.390 ;
        RECT 2380.020 3108.380 2383.020 3108.390 ;
        RECT 2560.020 3108.380 2563.020 3108.390 ;
        RECT 2740.020 3108.380 2743.020 3108.390 ;
        RECT 2945.000 3108.380 2948.000 3108.390 ;
        RECT -32.980 3105.380 2952.600 3108.380 ;
        RECT -28.380 3105.370 -25.380 3105.380 ;
        RECT 40.020 3105.370 43.020 3105.380 ;
        RECT 220.020 3105.370 223.020 3105.380 ;
        RECT 400.020 3105.370 403.020 3105.380 ;
        RECT 580.020 3105.370 583.020 3105.380 ;
        RECT 760.020 3105.370 763.020 3105.380 ;
        RECT 940.020 3105.370 943.020 3105.380 ;
        RECT 1120.020 3105.370 1123.020 3105.380 ;
        RECT 1300.020 3105.370 1303.020 3105.380 ;
        RECT 1480.020 3105.370 1483.020 3105.380 ;
        RECT 1660.020 3105.370 1663.020 3105.380 ;
        RECT 1840.020 3105.370 1843.020 3105.380 ;
        RECT 2020.020 3105.370 2023.020 3105.380 ;
        RECT 2200.020 3105.370 2203.020 3105.380 ;
        RECT 2380.020 3105.370 2383.020 3105.380 ;
        RECT 2560.020 3105.370 2563.020 3105.380 ;
        RECT 2740.020 3105.370 2743.020 3105.380 ;
        RECT 2945.000 3105.370 2948.000 3105.380 ;
        RECT -28.380 2928.380 -25.380 2928.390 ;
        RECT 40.020 2928.380 43.020 2928.390 ;
        RECT 220.020 2928.380 223.020 2928.390 ;
        RECT 400.020 2928.380 403.020 2928.390 ;
        RECT 580.020 2928.380 583.020 2928.390 ;
        RECT 760.020 2928.380 763.020 2928.390 ;
        RECT 940.020 2928.380 943.020 2928.390 ;
        RECT 1120.020 2928.380 1123.020 2928.390 ;
        RECT 1300.020 2928.380 1303.020 2928.390 ;
        RECT 1480.020 2928.380 1483.020 2928.390 ;
        RECT 1660.020 2928.380 1663.020 2928.390 ;
        RECT 1840.020 2928.380 1843.020 2928.390 ;
        RECT 2020.020 2928.380 2023.020 2928.390 ;
        RECT 2200.020 2928.380 2203.020 2928.390 ;
        RECT 2380.020 2928.380 2383.020 2928.390 ;
        RECT 2560.020 2928.380 2563.020 2928.390 ;
        RECT 2740.020 2928.380 2743.020 2928.390 ;
        RECT 2945.000 2928.380 2948.000 2928.390 ;
        RECT -32.980 2925.380 2952.600 2928.380 ;
        RECT -28.380 2925.370 -25.380 2925.380 ;
        RECT 40.020 2925.370 43.020 2925.380 ;
        RECT 220.020 2925.370 223.020 2925.380 ;
        RECT 400.020 2925.370 403.020 2925.380 ;
        RECT 580.020 2925.370 583.020 2925.380 ;
        RECT 760.020 2925.370 763.020 2925.380 ;
        RECT 940.020 2925.370 943.020 2925.380 ;
        RECT 1120.020 2925.370 1123.020 2925.380 ;
        RECT 1300.020 2925.370 1303.020 2925.380 ;
        RECT 1480.020 2925.370 1483.020 2925.380 ;
        RECT 1660.020 2925.370 1663.020 2925.380 ;
        RECT 1840.020 2925.370 1843.020 2925.380 ;
        RECT 2020.020 2925.370 2023.020 2925.380 ;
        RECT 2200.020 2925.370 2203.020 2925.380 ;
        RECT 2380.020 2925.370 2383.020 2925.380 ;
        RECT 2560.020 2925.370 2563.020 2925.380 ;
        RECT 2740.020 2925.370 2743.020 2925.380 ;
        RECT 2945.000 2925.370 2948.000 2925.380 ;
        RECT -28.380 2748.380 -25.380 2748.390 ;
        RECT 40.020 2748.380 43.020 2748.390 ;
        RECT 220.020 2748.380 223.020 2748.390 ;
        RECT 400.020 2748.380 403.020 2748.390 ;
        RECT 580.020 2748.380 583.020 2748.390 ;
        RECT 760.020 2748.380 763.020 2748.390 ;
        RECT 940.020 2748.380 943.020 2748.390 ;
        RECT 1120.020 2748.380 1123.020 2748.390 ;
        RECT 1300.020 2748.380 1303.020 2748.390 ;
        RECT 1480.020 2748.380 1483.020 2748.390 ;
        RECT 1660.020 2748.380 1663.020 2748.390 ;
        RECT 1840.020 2748.380 1843.020 2748.390 ;
        RECT 2020.020 2748.380 2023.020 2748.390 ;
        RECT 2200.020 2748.380 2203.020 2748.390 ;
        RECT 2380.020 2748.380 2383.020 2748.390 ;
        RECT 2560.020 2748.380 2563.020 2748.390 ;
        RECT 2740.020 2748.380 2743.020 2748.390 ;
        RECT 2945.000 2748.380 2948.000 2748.390 ;
        RECT -32.980 2745.380 2952.600 2748.380 ;
        RECT -28.380 2745.370 -25.380 2745.380 ;
        RECT 40.020 2745.370 43.020 2745.380 ;
        RECT 220.020 2745.370 223.020 2745.380 ;
        RECT 400.020 2745.370 403.020 2745.380 ;
        RECT 580.020 2745.370 583.020 2745.380 ;
        RECT 760.020 2745.370 763.020 2745.380 ;
        RECT 940.020 2745.370 943.020 2745.380 ;
        RECT 1120.020 2745.370 1123.020 2745.380 ;
        RECT 1300.020 2745.370 1303.020 2745.380 ;
        RECT 1480.020 2745.370 1483.020 2745.380 ;
        RECT 1660.020 2745.370 1663.020 2745.380 ;
        RECT 1840.020 2745.370 1843.020 2745.380 ;
        RECT 2020.020 2745.370 2023.020 2745.380 ;
        RECT 2200.020 2745.370 2203.020 2745.380 ;
        RECT 2380.020 2745.370 2383.020 2745.380 ;
        RECT 2560.020 2745.370 2563.020 2745.380 ;
        RECT 2740.020 2745.370 2743.020 2745.380 ;
        RECT 2945.000 2745.370 2948.000 2745.380 ;
        RECT -28.380 2568.380 -25.380 2568.390 ;
        RECT 40.020 2568.380 43.020 2568.390 ;
        RECT 220.020 2568.380 223.020 2568.390 ;
        RECT 400.020 2568.380 403.020 2568.390 ;
        RECT 580.020 2568.380 583.020 2568.390 ;
        RECT 760.020 2568.380 763.020 2568.390 ;
        RECT 940.020 2568.380 943.020 2568.390 ;
        RECT 1120.020 2568.380 1123.020 2568.390 ;
        RECT 1300.020 2568.380 1303.020 2568.390 ;
        RECT 1480.020 2568.380 1483.020 2568.390 ;
        RECT 1660.020 2568.380 1663.020 2568.390 ;
        RECT 1840.020 2568.380 1843.020 2568.390 ;
        RECT 2020.020 2568.380 2023.020 2568.390 ;
        RECT 2200.020 2568.380 2203.020 2568.390 ;
        RECT 2380.020 2568.380 2383.020 2568.390 ;
        RECT 2560.020 2568.380 2563.020 2568.390 ;
        RECT 2740.020 2568.380 2743.020 2568.390 ;
        RECT 2945.000 2568.380 2948.000 2568.390 ;
        RECT -32.980 2565.380 2952.600 2568.380 ;
        RECT -28.380 2565.370 -25.380 2565.380 ;
        RECT 40.020 2565.370 43.020 2565.380 ;
        RECT 220.020 2565.370 223.020 2565.380 ;
        RECT 400.020 2565.370 403.020 2565.380 ;
        RECT 580.020 2565.370 583.020 2565.380 ;
        RECT 760.020 2565.370 763.020 2565.380 ;
        RECT 940.020 2565.370 943.020 2565.380 ;
        RECT 1120.020 2565.370 1123.020 2565.380 ;
        RECT 1300.020 2565.370 1303.020 2565.380 ;
        RECT 1480.020 2565.370 1483.020 2565.380 ;
        RECT 1660.020 2565.370 1663.020 2565.380 ;
        RECT 1840.020 2565.370 1843.020 2565.380 ;
        RECT 2020.020 2565.370 2023.020 2565.380 ;
        RECT 2200.020 2565.370 2203.020 2565.380 ;
        RECT 2380.020 2565.370 2383.020 2565.380 ;
        RECT 2560.020 2565.370 2563.020 2565.380 ;
        RECT 2740.020 2565.370 2743.020 2565.380 ;
        RECT 2945.000 2565.370 2948.000 2565.380 ;
        RECT -28.380 2388.380 -25.380 2388.390 ;
        RECT 40.020 2388.380 43.020 2388.390 ;
        RECT 220.020 2388.380 223.020 2388.390 ;
        RECT 400.020 2388.380 403.020 2388.390 ;
        RECT 580.020 2388.380 583.020 2388.390 ;
        RECT 760.020 2388.380 763.020 2388.390 ;
        RECT 940.020 2388.380 943.020 2388.390 ;
        RECT 1120.020 2388.380 1123.020 2388.390 ;
        RECT 1300.020 2388.380 1303.020 2388.390 ;
        RECT 1480.020 2388.380 1483.020 2388.390 ;
        RECT 1660.020 2388.380 1663.020 2388.390 ;
        RECT 1840.020 2388.380 1843.020 2388.390 ;
        RECT 2020.020 2388.380 2023.020 2388.390 ;
        RECT 2200.020 2388.380 2203.020 2388.390 ;
        RECT 2380.020 2388.380 2383.020 2388.390 ;
        RECT 2560.020 2388.380 2563.020 2388.390 ;
        RECT 2740.020 2388.380 2743.020 2388.390 ;
        RECT 2945.000 2388.380 2948.000 2388.390 ;
        RECT -32.980 2385.380 2952.600 2388.380 ;
        RECT -28.380 2385.370 -25.380 2385.380 ;
        RECT 40.020 2385.370 43.020 2385.380 ;
        RECT 220.020 2385.370 223.020 2385.380 ;
        RECT 400.020 2385.370 403.020 2385.380 ;
        RECT 580.020 2385.370 583.020 2385.380 ;
        RECT 760.020 2385.370 763.020 2385.380 ;
        RECT 940.020 2385.370 943.020 2385.380 ;
        RECT 1120.020 2385.370 1123.020 2385.380 ;
        RECT 1300.020 2385.370 1303.020 2385.380 ;
        RECT 1480.020 2385.370 1483.020 2385.380 ;
        RECT 1660.020 2385.370 1663.020 2385.380 ;
        RECT 1840.020 2385.370 1843.020 2385.380 ;
        RECT 2020.020 2385.370 2023.020 2385.380 ;
        RECT 2200.020 2385.370 2203.020 2385.380 ;
        RECT 2380.020 2385.370 2383.020 2385.380 ;
        RECT 2560.020 2385.370 2563.020 2385.380 ;
        RECT 2740.020 2385.370 2743.020 2385.380 ;
        RECT 2945.000 2385.370 2948.000 2385.380 ;
        RECT -28.380 2208.380 -25.380 2208.390 ;
        RECT 40.020 2208.380 43.020 2208.390 ;
        RECT 220.020 2208.380 223.020 2208.390 ;
        RECT 400.020 2208.380 403.020 2208.390 ;
        RECT 580.020 2208.380 583.020 2208.390 ;
        RECT 760.020 2208.380 763.020 2208.390 ;
        RECT 940.020 2208.380 943.020 2208.390 ;
        RECT 1120.020 2208.380 1123.020 2208.390 ;
        RECT 1300.020 2208.380 1303.020 2208.390 ;
        RECT 1480.020 2208.380 1483.020 2208.390 ;
        RECT 1660.020 2208.380 1663.020 2208.390 ;
        RECT 1840.020 2208.380 1843.020 2208.390 ;
        RECT 2020.020 2208.380 2023.020 2208.390 ;
        RECT 2200.020 2208.380 2203.020 2208.390 ;
        RECT 2380.020 2208.380 2383.020 2208.390 ;
        RECT 2560.020 2208.380 2563.020 2208.390 ;
        RECT 2740.020 2208.380 2743.020 2208.390 ;
        RECT 2945.000 2208.380 2948.000 2208.390 ;
        RECT -32.980 2205.380 2952.600 2208.380 ;
        RECT -28.380 2205.370 -25.380 2205.380 ;
        RECT 40.020 2205.370 43.020 2205.380 ;
        RECT 220.020 2205.370 223.020 2205.380 ;
        RECT 400.020 2205.370 403.020 2205.380 ;
        RECT 580.020 2205.370 583.020 2205.380 ;
        RECT 760.020 2205.370 763.020 2205.380 ;
        RECT 940.020 2205.370 943.020 2205.380 ;
        RECT 1120.020 2205.370 1123.020 2205.380 ;
        RECT 1300.020 2205.370 1303.020 2205.380 ;
        RECT 1480.020 2205.370 1483.020 2205.380 ;
        RECT 1660.020 2205.370 1663.020 2205.380 ;
        RECT 1840.020 2205.370 1843.020 2205.380 ;
        RECT 2020.020 2205.370 2023.020 2205.380 ;
        RECT 2200.020 2205.370 2203.020 2205.380 ;
        RECT 2380.020 2205.370 2383.020 2205.380 ;
        RECT 2560.020 2205.370 2563.020 2205.380 ;
        RECT 2740.020 2205.370 2743.020 2205.380 ;
        RECT 2945.000 2205.370 2948.000 2205.380 ;
        RECT -28.380 2028.380 -25.380 2028.390 ;
        RECT 40.020 2028.380 43.020 2028.390 ;
        RECT 220.020 2028.380 223.020 2028.390 ;
        RECT 400.020 2028.380 403.020 2028.390 ;
        RECT 580.020 2028.380 583.020 2028.390 ;
        RECT 760.020 2028.380 763.020 2028.390 ;
        RECT 940.020 2028.380 943.020 2028.390 ;
        RECT 1120.020 2028.380 1123.020 2028.390 ;
        RECT 1300.020 2028.380 1303.020 2028.390 ;
        RECT 1480.020 2028.380 1483.020 2028.390 ;
        RECT 1660.020 2028.380 1663.020 2028.390 ;
        RECT 1840.020 2028.380 1843.020 2028.390 ;
        RECT 2020.020 2028.380 2023.020 2028.390 ;
        RECT 2200.020 2028.380 2203.020 2028.390 ;
        RECT 2380.020 2028.380 2383.020 2028.390 ;
        RECT 2560.020 2028.380 2563.020 2028.390 ;
        RECT 2740.020 2028.380 2743.020 2028.390 ;
        RECT 2945.000 2028.380 2948.000 2028.390 ;
        RECT -32.980 2025.380 2952.600 2028.380 ;
        RECT -28.380 2025.370 -25.380 2025.380 ;
        RECT 40.020 2025.370 43.020 2025.380 ;
        RECT 220.020 2025.370 223.020 2025.380 ;
        RECT 400.020 2025.370 403.020 2025.380 ;
        RECT 580.020 2025.370 583.020 2025.380 ;
        RECT 760.020 2025.370 763.020 2025.380 ;
        RECT 940.020 2025.370 943.020 2025.380 ;
        RECT 1120.020 2025.370 1123.020 2025.380 ;
        RECT 1300.020 2025.370 1303.020 2025.380 ;
        RECT 1480.020 2025.370 1483.020 2025.380 ;
        RECT 1660.020 2025.370 1663.020 2025.380 ;
        RECT 1840.020 2025.370 1843.020 2025.380 ;
        RECT 2020.020 2025.370 2023.020 2025.380 ;
        RECT 2200.020 2025.370 2203.020 2025.380 ;
        RECT 2380.020 2025.370 2383.020 2025.380 ;
        RECT 2560.020 2025.370 2563.020 2025.380 ;
        RECT 2740.020 2025.370 2743.020 2025.380 ;
        RECT 2945.000 2025.370 2948.000 2025.380 ;
        RECT -28.380 1848.380 -25.380 1848.390 ;
        RECT 40.020 1848.380 43.020 1848.390 ;
        RECT 220.020 1848.380 223.020 1848.390 ;
        RECT 400.020 1848.380 403.020 1848.390 ;
        RECT 580.020 1848.380 583.020 1848.390 ;
        RECT 760.020 1848.380 763.020 1848.390 ;
        RECT 940.020 1848.380 943.020 1848.390 ;
        RECT 1120.020 1848.380 1123.020 1848.390 ;
        RECT 1300.020 1848.380 1303.020 1848.390 ;
        RECT 1480.020 1848.380 1483.020 1848.390 ;
        RECT 1660.020 1848.380 1663.020 1848.390 ;
        RECT 1840.020 1848.380 1843.020 1848.390 ;
        RECT 2020.020 1848.380 2023.020 1848.390 ;
        RECT 2200.020 1848.380 2203.020 1848.390 ;
        RECT 2380.020 1848.380 2383.020 1848.390 ;
        RECT 2560.020 1848.380 2563.020 1848.390 ;
        RECT 2740.020 1848.380 2743.020 1848.390 ;
        RECT 2945.000 1848.380 2948.000 1848.390 ;
        RECT -32.980 1845.380 2952.600 1848.380 ;
        RECT -28.380 1845.370 -25.380 1845.380 ;
        RECT 40.020 1845.370 43.020 1845.380 ;
        RECT 220.020 1845.370 223.020 1845.380 ;
        RECT 400.020 1845.370 403.020 1845.380 ;
        RECT 580.020 1845.370 583.020 1845.380 ;
        RECT 760.020 1845.370 763.020 1845.380 ;
        RECT 940.020 1845.370 943.020 1845.380 ;
        RECT 1120.020 1845.370 1123.020 1845.380 ;
        RECT 1300.020 1845.370 1303.020 1845.380 ;
        RECT 1480.020 1845.370 1483.020 1845.380 ;
        RECT 1660.020 1845.370 1663.020 1845.380 ;
        RECT 1840.020 1845.370 1843.020 1845.380 ;
        RECT 2020.020 1845.370 2023.020 1845.380 ;
        RECT 2200.020 1845.370 2203.020 1845.380 ;
        RECT 2380.020 1845.370 2383.020 1845.380 ;
        RECT 2560.020 1845.370 2563.020 1845.380 ;
        RECT 2740.020 1845.370 2743.020 1845.380 ;
        RECT 2945.000 1845.370 2948.000 1845.380 ;
        RECT -28.380 1668.380 -25.380 1668.390 ;
        RECT 40.020 1668.380 43.020 1668.390 ;
        RECT 220.020 1668.380 223.020 1668.390 ;
        RECT 400.020 1668.380 403.020 1668.390 ;
        RECT 580.020 1668.380 583.020 1668.390 ;
        RECT 760.020 1668.380 763.020 1668.390 ;
        RECT 940.020 1668.380 943.020 1668.390 ;
        RECT 1120.020 1668.380 1123.020 1668.390 ;
        RECT 1300.020 1668.380 1303.020 1668.390 ;
        RECT 1480.020 1668.380 1483.020 1668.390 ;
        RECT 1660.020 1668.380 1663.020 1668.390 ;
        RECT 1840.020 1668.380 1843.020 1668.390 ;
        RECT 2020.020 1668.380 2023.020 1668.390 ;
        RECT 2200.020 1668.380 2203.020 1668.390 ;
        RECT 2380.020 1668.380 2383.020 1668.390 ;
        RECT 2560.020 1668.380 2563.020 1668.390 ;
        RECT 2740.020 1668.380 2743.020 1668.390 ;
        RECT 2945.000 1668.380 2948.000 1668.390 ;
        RECT -32.980 1665.380 2952.600 1668.380 ;
        RECT -28.380 1665.370 -25.380 1665.380 ;
        RECT 40.020 1665.370 43.020 1665.380 ;
        RECT 220.020 1665.370 223.020 1665.380 ;
        RECT 400.020 1665.370 403.020 1665.380 ;
        RECT 580.020 1665.370 583.020 1665.380 ;
        RECT 760.020 1665.370 763.020 1665.380 ;
        RECT 940.020 1665.370 943.020 1665.380 ;
        RECT 1120.020 1665.370 1123.020 1665.380 ;
        RECT 1300.020 1665.370 1303.020 1665.380 ;
        RECT 1480.020 1665.370 1483.020 1665.380 ;
        RECT 1660.020 1665.370 1663.020 1665.380 ;
        RECT 1840.020 1665.370 1843.020 1665.380 ;
        RECT 2020.020 1665.370 2023.020 1665.380 ;
        RECT 2200.020 1665.370 2203.020 1665.380 ;
        RECT 2380.020 1665.370 2383.020 1665.380 ;
        RECT 2560.020 1665.370 2563.020 1665.380 ;
        RECT 2740.020 1665.370 2743.020 1665.380 ;
        RECT 2945.000 1665.370 2948.000 1665.380 ;
        RECT -28.380 1488.380 -25.380 1488.390 ;
        RECT 40.020 1488.380 43.020 1488.390 ;
        RECT 220.020 1488.380 223.020 1488.390 ;
        RECT 400.020 1488.380 403.020 1488.390 ;
        RECT 580.020 1488.380 583.020 1488.390 ;
        RECT 760.020 1488.380 763.020 1488.390 ;
        RECT 940.020 1488.380 943.020 1488.390 ;
        RECT 1120.020 1488.380 1123.020 1488.390 ;
        RECT 1300.020 1488.380 1303.020 1488.390 ;
        RECT 1480.020 1488.380 1483.020 1488.390 ;
        RECT 1660.020 1488.380 1663.020 1488.390 ;
        RECT 1840.020 1488.380 1843.020 1488.390 ;
        RECT 2020.020 1488.380 2023.020 1488.390 ;
        RECT 2200.020 1488.380 2203.020 1488.390 ;
        RECT 2380.020 1488.380 2383.020 1488.390 ;
        RECT 2560.020 1488.380 2563.020 1488.390 ;
        RECT 2740.020 1488.380 2743.020 1488.390 ;
        RECT 2945.000 1488.380 2948.000 1488.390 ;
        RECT -32.980 1485.380 2952.600 1488.380 ;
        RECT -28.380 1485.370 -25.380 1485.380 ;
        RECT 40.020 1485.370 43.020 1485.380 ;
        RECT 220.020 1485.370 223.020 1485.380 ;
        RECT 400.020 1485.370 403.020 1485.380 ;
        RECT 580.020 1485.370 583.020 1485.380 ;
        RECT 760.020 1485.370 763.020 1485.380 ;
        RECT 940.020 1485.370 943.020 1485.380 ;
        RECT 1120.020 1485.370 1123.020 1485.380 ;
        RECT 1300.020 1485.370 1303.020 1485.380 ;
        RECT 1480.020 1485.370 1483.020 1485.380 ;
        RECT 1660.020 1485.370 1663.020 1485.380 ;
        RECT 1840.020 1485.370 1843.020 1485.380 ;
        RECT 2020.020 1485.370 2023.020 1485.380 ;
        RECT 2200.020 1485.370 2203.020 1485.380 ;
        RECT 2380.020 1485.370 2383.020 1485.380 ;
        RECT 2560.020 1485.370 2563.020 1485.380 ;
        RECT 2740.020 1485.370 2743.020 1485.380 ;
        RECT 2945.000 1485.370 2948.000 1485.380 ;
        RECT -28.380 1308.380 -25.380 1308.390 ;
        RECT 40.020 1308.380 43.020 1308.390 ;
        RECT 220.020 1308.380 223.020 1308.390 ;
        RECT 400.020 1308.380 403.020 1308.390 ;
        RECT 580.020 1308.380 583.020 1308.390 ;
        RECT 760.020 1308.380 763.020 1308.390 ;
        RECT 940.020 1308.380 943.020 1308.390 ;
        RECT 1120.020 1308.380 1123.020 1308.390 ;
        RECT 1300.020 1308.380 1303.020 1308.390 ;
        RECT 1480.020 1308.380 1483.020 1308.390 ;
        RECT 1660.020 1308.380 1663.020 1308.390 ;
        RECT 1840.020 1308.380 1843.020 1308.390 ;
        RECT 2020.020 1308.380 2023.020 1308.390 ;
        RECT 2200.020 1308.380 2203.020 1308.390 ;
        RECT 2380.020 1308.380 2383.020 1308.390 ;
        RECT 2560.020 1308.380 2563.020 1308.390 ;
        RECT 2740.020 1308.380 2743.020 1308.390 ;
        RECT 2945.000 1308.380 2948.000 1308.390 ;
        RECT -32.980 1305.380 2952.600 1308.380 ;
        RECT -28.380 1305.370 -25.380 1305.380 ;
        RECT 40.020 1305.370 43.020 1305.380 ;
        RECT 220.020 1305.370 223.020 1305.380 ;
        RECT 400.020 1305.370 403.020 1305.380 ;
        RECT 580.020 1305.370 583.020 1305.380 ;
        RECT 760.020 1305.370 763.020 1305.380 ;
        RECT 940.020 1305.370 943.020 1305.380 ;
        RECT 1120.020 1305.370 1123.020 1305.380 ;
        RECT 1300.020 1305.370 1303.020 1305.380 ;
        RECT 1480.020 1305.370 1483.020 1305.380 ;
        RECT 1660.020 1305.370 1663.020 1305.380 ;
        RECT 1840.020 1305.370 1843.020 1305.380 ;
        RECT 2020.020 1305.370 2023.020 1305.380 ;
        RECT 2200.020 1305.370 2203.020 1305.380 ;
        RECT 2380.020 1305.370 2383.020 1305.380 ;
        RECT 2560.020 1305.370 2563.020 1305.380 ;
        RECT 2740.020 1305.370 2743.020 1305.380 ;
        RECT 2945.000 1305.370 2948.000 1305.380 ;
        RECT -28.380 1128.380 -25.380 1128.390 ;
        RECT 40.020 1128.380 43.020 1128.390 ;
        RECT 220.020 1128.380 223.020 1128.390 ;
        RECT 400.020 1128.380 403.020 1128.390 ;
        RECT 580.020 1128.380 583.020 1128.390 ;
        RECT 760.020 1128.380 763.020 1128.390 ;
        RECT 940.020 1128.380 943.020 1128.390 ;
        RECT 1120.020 1128.380 1123.020 1128.390 ;
        RECT 1300.020 1128.380 1303.020 1128.390 ;
        RECT 1480.020 1128.380 1483.020 1128.390 ;
        RECT 1660.020 1128.380 1663.020 1128.390 ;
        RECT 1840.020 1128.380 1843.020 1128.390 ;
        RECT 2020.020 1128.380 2023.020 1128.390 ;
        RECT 2200.020 1128.380 2203.020 1128.390 ;
        RECT 2380.020 1128.380 2383.020 1128.390 ;
        RECT 2560.020 1128.380 2563.020 1128.390 ;
        RECT 2740.020 1128.380 2743.020 1128.390 ;
        RECT 2945.000 1128.380 2948.000 1128.390 ;
        RECT -32.980 1125.380 2952.600 1128.380 ;
        RECT -28.380 1125.370 -25.380 1125.380 ;
        RECT 40.020 1125.370 43.020 1125.380 ;
        RECT 220.020 1125.370 223.020 1125.380 ;
        RECT 400.020 1125.370 403.020 1125.380 ;
        RECT 580.020 1125.370 583.020 1125.380 ;
        RECT 760.020 1125.370 763.020 1125.380 ;
        RECT 940.020 1125.370 943.020 1125.380 ;
        RECT 1120.020 1125.370 1123.020 1125.380 ;
        RECT 1300.020 1125.370 1303.020 1125.380 ;
        RECT 1480.020 1125.370 1483.020 1125.380 ;
        RECT 1660.020 1125.370 1663.020 1125.380 ;
        RECT 1840.020 1125.370 1843.020 1125.380 ;
        RECT 2020.020 1125.370 2023.020 1125.380 ;
        RECT 2200.020 1125.370 2203.020 1125.380 ;
        RECT 2380.020 1125.370 2383.020 1125.380 ;
        RECT 2560.020 1125.370 2563.020 1125.380 ;
        RECT 2740.020 1125.370 2743.020 1125.380 ;
        RECT 2945.000 1125.370 2948.000 1125.380 ;
        RECT -28.380 948.380 -25.380 948.390 ;
        RECT 40.020 948.380 43.020 948.390 ;
        RECT 220.020 948.380 223.020 948.390 ;
        RECT 400.020 948.380 403.020 948.390 ;
        RECT 580.020 948.380 583.020 948.390 ;
        RECT 760.020 948.380 763.020 948.390 ;
        RECT 940.020 948.380 943.020 948.390 ;
        RECT 1120.020 948.380 1123.020 948.390 ;
        RECT 1300.020 948.380 1303.020 948.390 ;
        RECT 1480.020 948.380 1483.020 948.390 ;
        RECT 1660.020 948.380 1663.020 948.390 ;
        RECT 1840.020 948.380 1843.020 948.390 ;
        RECT 2020.020 948.380 2023.020 948.390 ;
        RECT 2200.020 948.380 2203.020 948.390 ;
        RECT 2380.020 948.380 2383.020 948.390 ;
        RECT 2560.020 948.380 2563.020 948.390 ;
        RECT 2740.020 948.380 2743.020 948.390 ;
        RECT 2945.000 948.380 2948.000 948.390 ;
        RECT -32.980 945.380 2952.600 948.380 ;
        RECT -28.380 945.370 -25.380 945.380 ;
        RECT 40.020 945.370 43.020 945.380 ;
        RECT 220.020 945.370 223.020 945.380 ;
        RECT 400.020 945.370 403.020 945.380 ;
        RECT 580.020 945.370 583.020 945.380 ;
        RECT 760.020 945.370 763.020 945.380 ;
        RECT 940.020 945.370 943.020 945.380 ;
        RECT 1120.020 945.370 1123.020 945.380 ;
        RECT 1300.020 945.370 1303.020 945.380 ;
        RECT 1480.020 945.370 1483.020 945.380 ;
        RECT 1660.020 945.370 1663.020 945.380 ;
        RECT 1840.020 945.370 1843.020 945.380 ;
        RECT 2020.020 945.370 2023.020 945.380 ;
        RECT 2200.020 945.370 2203.020 945.380 ;
        RECT 2380.020 945.370 2383.020 945.380 ;
        RECT 2560.020 945.370 2563.020 945.380 ;
        RECT 2740.020 945.370 2743.020 945.380 ;
        RECT 2945.000 945.370 2948.000 945.380 ;
        RECT -28.380 768.380 -25.380 768.390 ;
        RECT 40.020 768.380 43.020 768.390 ;
        RECT 220.020 768.380 223.020 768.390 ;
        RECT 400.020 768.380 403.020 768.390 ;
        RECT 580.020 768.380 583.020 768.390 ;
        RECT 760.020 768.380 763.020 768.390 ;
        RECT 940.020 768.380 943.020 768.390 ;
        RECT 1120.020 768.380 1123.020 768.390 ;
        RECT 1300.020 768.380 1303.020 768.390 ;
        RECT 1480.020 768.380 1483.020 768.390 ;
        RECT 1660.020 768.380 1663.020 768.390 ;
        RECT 1840.020 768.380 1843.020 768.390 ;
        RECT 2020.020 768.380 2023.020 768.390 ;
        RECT 2200.020 768.380 2203.020 768.390 ;
        RECT 2380.020 768.380 2383.020 768.390 ;
        RECT 2560.020 768.380 2563.020 768.390 ;
        RECT 2740.020 768.380 2743.020 768.390 ;
        RECT 2945.000 768.380 2948.000 768.390 ;
        RECT -32.980 765.380 2952.600 768.380 ;
        RECT -28.380 765.370 -25.380 765.380 ;
        RECT 40.020 765.370 43.020 765.380 ;
        RECT 220.020 765.370 223.020 765.380 ;
        RECT 400.020 765.370 403.020 765.380 ;
        RECT 580.020 765.370 583.020 765.380 ;
        RECT 760.020 765.370 763.020 765.380 ;
        RECT 940.020 765.370 943.020 765.380 ;
        RECT 1120.020 765.370 1123.020 765.380 ;
        RECT 1300.020 765.370 1303.020 765.380 ;
        RECT 1480.020 765.370 1483.020 765.380 ;
        RECT 1660.020 765.370 1663.020 765.380 ;
        RECT 1840.020 765.370 1843.020 765.380 ;
        RECT 2020.020 765.370 2023.020 765.380 ;
        RECT 2200.020 765.370 2203.020 765.380 ;
        RECT 2380.020 765.370 2383.020 765.380 ;
        RECT 2560.020 765.370 2563.020 765.380 ;
        RECT 2740.020 765.370 2743.020 765.380 ;
        RECT 2945.000 765.370 2948.000 765.380 ;
        RECT -28.380 588.380 -25.380 588.390 ;
        RECT 40.020 588.380 43.020 588.390 ;
        RECT 220.020 588.380 223.020 588.390 ;
        RECT 400.020 588.380 403.020 588.390 ;
        RECT 580.020 588.380 583.020 588.390 ;
        RECT 760.020 588.380 763.020 588.390 ;
        RECT 940.020 588.380 943.020 588.390 ;
        RECT 1120.020 588.380 1123.020 588.390 ;
        RECT 1300.020 588.380 1303.020 588.390 ;
        RECT 1480.020 588.380 1483.020 588.390 ;
        RECT 1660.020 588.380 1663.020 588.390 ;
        RECT 1840.020 588.380 1843.020 588.390 ;
        RECT 2020.020 588.380 2023.020 588.390 ;
        RECT 2200.020 588.380 2203.020 588.390 ;
        RECT 2380.020 588.380 2383.020 588.390 ;
        RECT 2560.020 588.380 2563.020 588.390 ;
        RECT 2740.020 588.380 2743.020 588.390 ;
        RECT 2945.000 588.380 2948.000 588.390 ;
        RECT -32.980 585.380 2952.600 588.380 ;
        RECT -28.380 585.370 -25.380 585.380 ;
        RECT 40.020 585.370 43.020 585.380 ;
        RECT 220.020 585.370 223.020 585.380 ;
        RECT 400.020 585.370 403.020 585.380 ;
        RECT 580.020 585.370 583.020 585.380 ;
        RECT 760.020 585.370 763.020 585.380 ;
        RECT 940.020 585.370 943.020 585.380 ;
        RECT 1120.020 585.370 1123.020 585.380 ;
        RECT 1300.020 585.370 1303.020 585.380 ;
        RECT 1480.020 585.370 1483.020 585.380 ;
        RECT 1660.020 585.370 1663.020 585.380 ;
        RECT 1840.020 585.370 1843.020 585.380 ;
        RECT 2020.020 585.370 2023.020 585.380 ;
        RECT 2200.020 585.370 2203.020 585.380 ;
        RECT 2380.020 585.370 2383.020 585.380 ;
        RECT 2560.020 585.370 2563.020 585.380 ;
        RECT 2740.020 585.370 2743.020 585.380 ;
        RECT 2945.000 585.370 2948.000 585.380 ;
        RECT -28.380 408.380 -25.380 408.390 ;
        RECT 40.020 408.380 43.020 408.390 ;
        RECT 220.020 408.380 223.020 408.390 ;
        RECT 400.020 408.380 403.020 408.390 ;
        RECT 580.020 408.380 583.020 408.390 ;
        RECT 760.020 408.380 763.020 408.390 ;
        RECT 940.020 408.380 943.020 408.390 ;
        RECT 1120.020 408.380 1123.020 408.390 ;
        RECT 1300.020 408.380 1303.020 408.390 ;
        RECT 1480.020 408.380 1483.020 408.390 ;
        RECT 1660.020 408.380 1663.020 408.390 ;
        RECT 1840.020 408.380 1843.020 408.390 ;
        RECT 2020.020 408.380 2023.020 408.390 ;
        RECT 2200.020 408.380 2203.020 408.390 ;
        RECT 2380.020 408.380 2383.020 408.390 ;
        RECT 2560.020 408.380 2563.020 408.390 ;
        RECT 2740.020 408.380 2743.020 408.390 ;
        RECT 2945.000 408.380 2948.000 408.390 ;
        RECT -32.980 405.380 2952.600 408.380 ;
        RECT -28.380 405.370 -25.380 405.380 ;
        RECT 40.020 405.370 43.020 405.380 ;
        RECT 220.020 405.370 223.020 405.380 ;
        RECT 400.020 405.370 403.020 405.380 ;
        RECT 580.020 405.370 583.020 405.380 ;
        RECT 760.020 405.370 763.020 405.380 ;
        RECT 940.020 405.370 943.020 405.380 ;
        RECT 1120.020 405.370 1123.020 405.380 ;
        RECT 1300.020 405.370 1303.020 405.380 ;
        RECT 1480.020 405.370 1483.020 405.380 ;
        RECT 1660.020 405.370 1663.020 405.380 ;
        RECT 1840.020 405.370 1843.020 405.380 ;
        RECT 2020.020 405.370 2023.020 405.380 ;
        RECT 2200.020 405.370 2203.020 405.380 ;
        RECT 2380.020 405.370 2383.020 405.380 ;
        RECT 2560.020 405.370 2563.020 405.380 ;
        RECT 2740.020 405.370 2743.020 405.380 ;
        RECT 2945.000 405.370 2948.000 405.380 ;
        RECT -28.380 228.380 -25.380 228.390 ;
        RECT 40.020 228.380 43.020 228.390 ;
        RECT 220.020 228.380 223.020 228.390 ;
        RECT 400.020 228.380 403.020 228.390 ;
        RECT 580.020 228.380 583.020 228.390 ;
        RECT 760.020 228.380 763.020 228.390 ;
        RECT 940.020 228.380 943.020 228.390 ;
        RECT 1120.020 228.380 1123.020 228.390 ;
        RECT 1300.020 228.380 1303.020 228.390 ;
        RECT 1480.020 228.380 1483.020 228.390 ;
        RECT 1660.020 228.380 1663.020 228.390 ;
        RECT 1840.020 228.380 1843.020 228.390 ;
        RECT 2020.020 228.380 2023.020 228.390 ;
        RECT 2200.020 228.380 2203.020 228.390 ;
        RECT 2380.020 228.380 2383.020 228.390 ;
        RECT 2560.020 228.380 2563.020 228.390 ;
        RECT 2740.020 228.380 2743.020 228.390 ;
        RECT 2945.000 228.380 2948.000 228.390 ;
        RECT -32.980 225.380 2952.600 228.380 ;
        RECT -28.380 225.370 -25.380 225.380 ;
        RECT 40.020 225.370 43.020 225.380 ;
        RECT 220.020 225.370 223.020 225.380 ;
        RECT 400.020 225.370 403.020 225.380 ;
        RECT 580.020 225.370 583.020 225.380 ;
        RECT 760.020 225.370 763.020 225.380 ;
        RECT 940.020 225.370 943.020 225.380 ;
        RECT 1120.020 225.370 1123.020 225.380 ;
        RECT 1300.020 225.370 1303.020 225.380 ;
        RECT 1480.020 225.370 1483.020 225.380 ;
        RECT 1660.020 225.370 1663.020 225.380 ;
        RECT 1840.020 225.370 1843.020 225.380 ;
        RECT 2020.020 225.370 2023.020 225.380 ;
        RECT 2200.020 225.370 2203.020 225.380 ;
        RECT 2380.020 225.370 2383.020 225.380 ;
        RECT 2560.020 225.370 2563.020 225.380 ;
        RECT 2740.020 225.370 2743.020 225.380 ;
        RECT 2945.000 225.370 2948.000 225.380 ;
        RECT -28.380 48.380 -25.380 48.390 ;
        RECT 40.020 48.380 43.020 48.390 ;
        RECT 220.020 48.380 223.020 48.390 ;
        RECT 400.020 48.380 403.020 48.390 ;
        RECT 580.020 48.380 583.020 48.390 ;
        RECT 760.020 48.380 763.020 48.390 ;
        RECT 940.020 48.380 943.020 48.390 ;
        RECT 1120.020 48.380 1123.020 48.390 ;
        RECT 1300.020 48.380 1303.020 48.390 ;
        RECT 1480.020 48.380 1483.020 48.390 ;
        RECT 1660.020 48.380 1663.020 48.390 ;
        RECT 1840.020 48.380 1843.020 48.390 ;
        RECT 2020.020 48.380 2023.020 48.390 ;
        RECT 2200.020 48.380 2203.020 48.390 ;
        RECT 2380.020 48.380 2383.020 48.390 ;
        RECT 2560.020 48.380 2563.020 48.390 ;
        RECT 2740.020 48.380 2743.020 48.390 ;
        RECT 2945.000 48.380 2948.000 48.390 ;
        RECT -32.980 45.380 2952.600 48.380 ;
        RECT -28.380 45.370 -25.380 45.380 ;
        RECT 40.020 45.370 43.020 45.380 ;
        RECT 220.020 45.370 223.020 45.380 ;
        RECT 400.020 45.370 403.020 45.380 ;
        RECT 580.020 45.370 583.020 45.380 ;
        RECT 760.020 45.370 763.020 45.380 ;
        RECT 940.020 45.370 943.020 45.380 ;
        RECT 1120.020 45.370 1123.020 45.380 ;
        RECT 1300.020 45.370 1303.020 45.380 ;
        RECT 1480.020 45.370 1483.020 45.380 ;
        RECT 1660.020 45.370 1663.020 45.380 ;
        RECT 1840.020 45.370 1843.020 45.380 ;
        RECT 2020.020 45.370 2023.020 45.380 ;
        RECT 2200.020 45.370 2203.020 45.380 ;
        RECT 2380.020 45.370 2383.020 45.380 ;
        RECT 2560.020 45.370 2563.020 45.380 ;
        RECT 2740.020 45.370 2743.020 45.380 ;
        RECT 2945.000 45.370 2948.000 45.380 ;
        RECT -28.380 -20.020 -25.380 -20.010 ;
        RECT 40.020 -20.020 43.020 -20.010 ;
        RECT 220.020 -20.020 223.020 -20.010 ;
        RECT 400.020 -20.020 403.020 -20.010 ;
        RECT 580.020 -20.020 583.020 -20.010 ;
        RECT 760.020 -20.020 763.020 -20.010 ;
        RECT 940.020 -20.020 943.020 -20.010 ;
        RECT 1120.020 -20.020 1123.020 -20.010 ;
        RECT 1300.020 -20.020 1303.020 -20.010 ;
        RECT 1480.020 -20.020 1483.020 -20.010 ;
        RECT 1660.020 -20.020 1663.020 -20.010 ;
        RECT 1840.020 -20.020 1843.020 -20.010 ;
        RECT 2020.020 -20.020 2023.020 -20.010 ;
        RECT 2200.020 -20.020 2203.020 -20.010 ;
        RECT 2380.020 -20.020 2383.020 -20.010 ;
        RECT 2560.020 -20.020 2563.020 -20.010 ;
        RECT 2740.020 -20.020 2743.020 -20.010 ;
        RECT 2945.000 -20.020 2948.000 -20.010 ;
        RECT -28.380 -23.020 2948.000 -20.020 ;
        RECT -28.380 -23.030 -25.380 -23.020 ;
        RECT 40.020 -23.030 43.020 -23.020 ;
        RECT 220.020 -23.030 223.020 -23.020 ;
        RECT 400.020 -23.030 403.020 -23.020 ;
        RECT 580.020 -23.030 583.020 -23.020 ;
        RECT 760.020 -23.030 763.020 -23.020 ;
        RECT 940.020 -23.030 943.020 -23.020 ;
        RECT 1120.020 -23.030 1123.020 -23.020 ;
        RECT 1300.020 -23.030 1303.020 -23.020 ;
        RECT 1480.020 -23.030 1483.020 -23.020 ;
        RECT 1660.020 -23.030 1663.020 -23.020 ;
        RECT 1840.020 -23.030 1843.020 -23.020 ;
        RECT 2020.020 -23.030 2023.020 -23.020 ;
        RECT 2200.020 -23.030 2203.020 -23.020 ;
        RECT 2380.020 -23.030 2383.020 -23.020 ;
        RECT 2560.020 -23.030 2563.020 -23.020 ;
        RECT 2740.020 -23.030 2743.020 -23.020 ;
        RECT 2945.000 -23.030 2948.000 -23.020 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -32.980 -27.620 -29.980 3547.300 ;
        RECT 130.020 -27.620 133.020 3547.300 ;
        RECT 310.020 -27.620 313.020 3547.300 ;
        RECT 490.020 -27.620 493.020 3547.300 ;
        RECT 670.020 -27.620 673.020 3547.300 ;
        RECT 850.020 -27.620 853.020 3547.300 ;
        RECT 1030.020 -27.620 1033.020 3547.300 ;
        RECT 1210.020 -27.620 1213.020 3547.300 ;
        RECT 1390.020 -27.620 1393.020 3547.300 ;
        RECT 1570.020 -27.620 1573.020 3547.300 ;
        RECT 1750.020 -27.620 1753.020 3547.300 ;
        RECT 1930.020 -27.620 1933.020 3547.300 ;
        RECT 2110.020 -27.620 2113.020 3547.300 ;
        RECT 2290.020 -27.620 2293.020 3547.300 ;
        RECT 2470.020 -27.620 2473.020 3547.300 ;
        RECT 2650.020 -27.620 2653.020 3547.300 ;
        RECT 2830.020 -27.620 2833.020 3547.300 ;
        RECT 2949.600 -27.620 2952.600 3547.300 ;
      LAYER via4 ;
        RECT -32.070 3546.010 -30.890 3547.190 ;
        RECT -32.070 3544.410 -30.890 3545.590 ;
        RECT -32.070 3377.090 -30.890 3378.270 ;
        RECT -32.070 3375.490 -30.890 3376.670 ;
        RECT -32.070 3197.090 -30.890 3198.270 ;
        RECT -32.070 3195.490 -30.890 3196.670 ;
        RECT -32.070 3017.090 -30.890 3018.270 ;
        RECT -32.070 3015.490 -30.890 3016.670 ;
        RECT -32.070 2837.090 -30.890 2838.270 ;
        RECT -32.070 2835.490 -30.890 2836.670 ;
        RECT -32.070 2657.090 -30.890 2658.270 ;
        RECT -32.070 2655.490 -30.890 2656.670 ;
        RECT -32.070 2477.090 -30.890 2478.270 ;
        RECT -32.070 2475.490 -30.890 2476.670 ;
        RECT -32.070 2297.090 -30.890 2298.270 ;
        RECT -32.070 2295.490 -30.890 2296.670 ;
        RECT -32.070 2117.090 -30.890 2118.270 ;
        RECT -32.070 2115.490 -30.890 2116.670 ;
        RECT -32.070 1937.090 -30.890 1938.270 ;
        RECT -32.070 1935.490 -30.890 1936.670 ;
        RECT -32.070 1757.090 -30.890 1758.270 ;
        RECT -32.070 1755.490 -30.890 1756.670 ;
        RECT -32.070 1577.090 -30.890 1578.270 ;
        RECT -32.070 1575.490 -30.890 1576.670 ;
        RECT -32.070 1397.090 -30.890 1398.270 ;
        RECT -32.070 1395.490 -30.890 1396.670 ;
        RECT -32.070 1217.090 -30.890 1218.270 ;
        RECT -32.070 1215.490 -30.890 1216.670 ;
        RECT -32.070 1037.090 -30.890 1038.270 ;
        RECT -32.070 1035.490 -30.890 1036.670 ;
        RECT -32.070 857.090 -30.890 858.270 ;
        RECT -32.070 855.490 -30.890 856.670 ;
        RECT -32.070 677.090 -30.890 678.270 ;
        RECT -32.070 675.490 -30.890 676.670 ;
        RECT -32.070 497.090 -30.890 498.270 ;
        RECT -32.070 495.490 -30.890 496.670 ;
        RECT -32.070 317.090 -30.890 318.270 ;
        RECT -32.070 315.490 -30.890 316.670 ;
        RECT -32.070 137.090 -30.890 138.270 ;
        RECT -32.070 135.490 -30.890 136.670 ;
        RECT -32.070 -25.910 -30.890 -24.730 ;
        RECT -32.070 -27.510 -30.890 -26.330 ;
        RECT 130.930 3546.010 132.110 3547.190 ;
        RECT 130.930 3544.410 132.110 3545.590 ;
        RECT 130.930 3377.090 132.110 3378.270 ;
        RECT 130.930 3375.490 132.110 3376.670 ;
        RECT 130.930 3197.090 132.110 3198.270 ;
        RECT 130.930 3195.490 132.110 3196.670 ;
        RECT 130.930 3017.090 132.110 3018.270 ;
        RECT 130.930 3015.490 132.110 3016.670 ;
        RECT 130.930 2837.090 132.110 2838.270 ;
        RECT 130.930 2835.490 132.110 2836.670 ;
        RECT 130.930 2657.090 132.110 2658.270 ;
        RECT 130.930 2655.490 132.110 2656.670 ;
        RECT 130.930 2477.090 132.110 2478.270 ;
        RECT 130.930 2475.490 132.110 2476.670 ;
        RECT 130.930 2297.090 132.110 2298.270 ;
        RECT 130.930 2295.490 132.110 2296.670 ;
        RECT 130.930 2117.090 132.110 2118.270 ;
        RECT 130.930 2115.490 132.110 2116.670 ;
        RECT 130.930 1937.090 132.110 1938.270 ;
        RECT 130.930 1935.490 132.110 1936.670 ;
        RECT 130.930 1757.090 132.110 1758.270 ;
        RECT 130.930 1755.490 132.110 1756.670 ;
        RECT 130.930 1577.090 132.110 1578.270 ;
        RECT 130.930 1575.490 132.110 1576.670 ;
        RECT 130.930 1397.090 132.110 1398.270 ;
        RECT 130.930 1395.490 132.110 1396.670 ;
        RECT 130.930 1217.090 132.110 1218.270 ;
        RECT 130.930 1215.490 132.110 1216.670 ;
        RECT 130.930 1037.090 132.110 1038.270 ;
        RECT 130.930 1035.490 132.110 1036.670 ;
        RECT 130.930 857.090 132.110 858.270 ;
        RECT 130.930 855.490 132.110 856.670 ;
        RECT 130.930 677.090 132.110 678.270 ;
        RECT 130.930 675.490 132.110 676.670 ;
        RECT 130.930 497.090 132.110 498.270 ;
        RECT 130.930 495.490 132.110 496.670 ;
        RECT 130.930 317.090 132.110 318.270 ;
        RECT 130.930 315.490 132.110 316.670 ;
        RECT 130.930 137.090 132.110 138.270 ;
        RECT 130.930 135.490 132.110 136.670 ;
        RECT 130.930 -25.910 132.110 -24.730 ;
        RECT 130.930 -27.510 132.110 -26.330 ;
        RECT 310.930 3546.010 312.110 3547.190 ;
        RECT 310.930 3544.410 312.110 3545.590 ;
        RECT 310.930 3377.090 312.110 3378.270 ;
        RECT 310.930 3375.490 312.110 3376.670 ;
        RECT 310.930 3197.090 312.110 3198.270 ;
        RECT 310.930 3195.490 312.110 3196.670 ;
        RECT 310.930 3017.090 312.110 3018.270 ;
        RECT 310.930 3015.490 312.110 3016.670 ;
        RECT 310.930 2837.090 312.110 2838.270 ;
        RECT 310.930 2835.490 312.110 2836.670 ;
        RECT 310.930 2657.090 312.110 2658.270 ;
        RECT 310.930 2655.490 312.110 2656.670 ;
        RECT 310.930 2477.090 312.110 2478.270 ;
        RECT 310.930 2475.490 312.110 2476.670 ;
        RECT 310.930 2297.090 312.110 2298.270 ;
        RECT 310.930 2295.490 312.110 2296.670 ;
        RECT 310.930 2117.090 312.110 2118.270 ;
        RECT 310.930 2115.490 312.110 2116.670 ;
        RECT 310.930 1937.090 312.110 1938.270 ;
        RECT 310.930 1935.490 312.110 1936.670 ;
        RECT 310.930 1757.090 312.110 1758.270 ;
        RECT 310.930 1755.490 312.110 1756.670 ;
        RECT 310.930 1577.090 312.110 1578.270 ;
        RECT 310.930 1575.490 312.110 1576.670 ;
        RECT 310.930 1397.090 312.110 1398.270 ;
        RECT 310.930 1395.490 312.110 1396.670 ;
        RECT 310.930 1217.090 312.110 1218.270 ;
        RECT 310.930 1215.490 312.110 1216.670 ;
        RECT 310.930 1037.090 312.110 1038.270 ;
        RECT 310.930 1035.490 312.110 1036.670 ;
        RECT 310.930 857.090 312.110 858.270 ;
        RECT 310.930 855.490 312.110 856.670 ;
        RECT 310.930 677.090 312.110 678.270 ;
        RECT 310.930 675.490 312.110 676.670 ;
        RECT 310.930 497.090 312.110 498.270 ;
        RECT 310.930 495.490 312.110 496.670 ;
        RECT 310.930 317.090 312.110 318.270 ;
        RECT 310.930 315.490 312.110 316.670 ;
        RECT 310.930 137.090 312.110 138.270 ;
        RECT 310.930 135.490 312.110 136.670 ;
        RECT 310.930 -25.910 312.110 -24.730 ;
        RECT 310.930 -27.510 312.110 -26.330 ;
        RECT 490.930 3546.010 492.110 3547.190 ;
        RECT 490.930 3544.410 492.110 3545.590 ;
        RECT 490.930 3377.090 492.110 3378.270 ;
        RECT 490.930 3375.490 492.110 3376.670 ;
        RECT 490.930 3197.090 492.110 3198.270 ;
        RECT 490.930 3195.490 492.110 3196.670 ;
        RECT 490.930 3017.090 492.110 3018.270 ;
        RECT 490.930 3015.490 492.110 3016.670 ;
        RECT 490.930 2837.090 492.110 2838.270 ;
        RECT 490.930 2835.490 492.110 2836.670 ;
        RECT 490.930 2657.090 492.110 2658.270 ;
        RECT 490.930 2655.490 492.110 2656.670 ;
        RECT 490.930 2477.090 492.110 2478.270 ;
        RECT 490.930 2475.490 492.110 2476.670 ;
        RECT 490.930 2297.090 492.110 2298.270 ;
        RECT 490.930 2295.490 492.110 2296.670 ;
        RECT 490.930 2117.090 492.110 2118.270 ;
        RECT 490.930 2115.490 492.110 2116.670 ;
        RECT 490.930 1937.090 492.110 1938.270 ;
        RECT 490.930 1935.490 492.110 1936.670 ;
        RECT 490.930 1757.090 492.110 1758.270 ;
        RECT 490.930 1755.490 492.110 1756.670 ;
        RECT 490.930 1577.090 492.110 1578.270 ;
        RECT 490.930 1575.490 492.110 1576.670 ;
        RECT 490.930 1397.090 492.110 1398.270 ;
        RECT 490.930 1395.490 492.110 1396.670 ;
        RECT 490.930 1217.090 492.110 1218.270 ;
        RECT 490.930 1215.490 492.110 1216.670 ;
        RECT 490.930 1037.090 492.110 1038.270 ;
        RECT 490.930 1035.490 492.110 1036.670 ;
        RECT 490.930 857.090 492.110 858.270 ;
        RECT 490.930 855.490 492.110 856.670 ;
        RECT 490.930 677.090 492.110 678.270 ;
        RECT 490.930 675.490 492.110 676.670 ;
        RECT 490.930 497.090 492.110 498.270 ;
        RECT 490.930 495.490 492.110 496.670 ;
        RECT 490.930 317.090 492.110 318.270 ;
        RECT 490.930 315.490 492.110 316.670 ;
        RECT 490.930 137.090 492.110 138.270 ;
        RECT 490.930 135.490 492.110 136.670 ;
        RECT 490.930 -25.910 492.110 -24.730 ;
        RECT 490.930 -27.510 492.110 -26.330 ;
        RECT 670.930 3546.010 672.110 3547.190 ;
        RECT 670.930 3544.410 672.110 3545.590 ;
        RECT 670.930 3377.090 672.110 3378.270 ;
        RECT 670.930 3375.490 672.110 3376.670 ;
        RECT 670.930 3197.090 672.110 3198.270 ;
        RECT 670.930 3195.490 672.110 3196.670 ;
        RECT 670.930 3017.090 672.110 3018.270 ;
        RECT 670.930 3015.490 672.110 3016.670 ;
        RECT 670.930 2837.090 672.110 2838.270 ;
        RECT 670.930 2835.490 672.110 2836.670 ;
        RECT 670.930 2657.090 672.110 2658.270 ;
        RECT 670.930 2655.490 672.110 2656.670 ;
        RECT 670.930 2477.090 672.110 2478.270 ;
        RECT 670.930 2475.490 672.110 2476.670 ;
        RECT 670.930 2297.090 672.110 2298.270 ;
        RECT 670.930 2295.490 672.110 2296.670 ;
        RECT 670.930 2117.090 672.110 2118.270 ;
        RECT 670.930 2115.490 672.110 2116.670 ;
        RECT 670.930 1937.090 672.110 1938.270 ;
        RECT 670.930 1935.490 672.110 1936.670 ;
        RECT 670.930 1757.090 672.110 1758.270 ;
        RECT 670.930 1755.490 672.110 1756.670 ;
        RECT 670.930 1577.090 672.110 1578.270 ;
        RECT 670.930 1575.490 672.110 1576.670 ;
        RECT 670.930 1397.090 672.110 1398.270 ;
        RECT 670.930 1395.490 672.110 1396.670 ;
        RECT 670.930 1217.090 672.110 1218.270 ;
        RECT 670.930 1215.490 672.110 1216.670 ;
        RECT 670.930 1037.090 672.110 1038.270 ;
        RECT 670.930 1035.490 672.110 1036.670 ;
        RECT 670.930 857.090 672.110 858.270 ;
        RECT 670.930 855.490 672.110 856.670 ;
        RECT 670.930 677.090 672.110 678.270 ;
        RECT 670.930 675.490 672.110 676.670 ;
        RECT 670.930 497.090 672.110 498.270 ;
        RECT 670.930 495.490 672.110 496.670 ;
        RECT 670.930 317.090 672.110 318.270 ;
        RECT 670.930 315.490 672.110 316.670 ;
        RECT 670.930 137.090 672.110 138.270 ;
        RECT 670.930 135.490 672.110 136.670 ;
        RECT 670.930 -25.910 672.110 -24.730 ;
        RECT 670.930 -27.510 672.110 -26.330 ;
        RECT 850.930 3546.010 852.110 3547.190 ;
        RECT 850.930 3544.410 852.110 3545.590 ;
        RECT 850.930 3377.090 852.110 3378.270 ;
        RECT 850.930 3375.490 852.110 3376.670 ;
        RECT 850.930 3197.090 852.110 3198.270 ;
        RECT 850.930 3195.490 852.110 3196.670 ;
        RECT 850.930 3017.090 852.110 3018.270 ;
        RECT 850.930 3015.490 852.110 3016.670 ;
        RECT 850.930 2837.090 852.110 2838.270 ;
        RECT 850.930 2835.490 852.110 2836.670 ;
        RECT 850.930 2657.090 852.110 2658.270 ;
        RECT 850.930 2655.490 852.110 2656.670 ;
        RECT 850.930 2477.090 852.110 2478.270 ;
        RECT 850.930 2475.490 852.110 2476.670 ;
        RECT 850.930 2297.090 852.110 2298.270 ;
        RECT 850.930 2295.490 852.110 2296.670 ;
        RECT 850.930 2117.090 852.110 2118.270 ;
        RECT 850.930 2115.490 852.110 2116.670 ;
        RECT 850.930 1937.090 852.110 1938.270 ;
        RECT 850.930 1935.490 852.110 1936.670 ;
        RECT 850.930 1757.090 852.110 1758.270 ;
        RECT 850.930 1755.490 852.110 1756.670 ;
        RECT 850.930 1577.090 852.110 1578.270 ;
        RECT 850.930 1575.490 852.110 1576.670 ;
        RECT 850.930 1397.090 852.110 1398.270 ;
        RECT 850.930 1395.490 852.110 1396.670 ;
        RECT 850.930 1217.090 852.110 1218.270 ;
        RECT 850.930 1215.490 852.110 1216.670 ;
        RECT 850.930 1037.090 852.110 1038.270 ;
        RECT 850.930 1035.490 852.110 1036.670 ;
        RECT 850.930 857.090 852.110 858.270 ;
        RECT 850.930 855.490 852.110 856.670 ;
        RECT 850.930 677.090 852.110 678.270 ;
        RECT 850.930 675.490 852.110 676.670 ;
        RECT 850.930 497.090 852.110 498.270 ;
        RECT 850.930 495.490 852.110 496.670 ;
        RECT 850.930 317.090 852.110 318.270 ;
        RECT 850.930 315.490 852.110 316.670 ;
        RECT 850.930 137.090 852.110 138.270 ;
        RECT 850.930 135.490 852.110 136.670 ;
        RECT 850.930 -25.910 852.110 -24.730 ;
        RECT 850.930 -27.510 852.110 -26.330 ;
        RECT 1030.930 3546.010 1032.110 3547.190 ;
        RECT 1030.930 3544.410 1032.110 3545.590 ;
        RECT 1030.930 3377.090 1032.110 3378.270 ;
        RECT 1030.930 3375.490 1032.110 3376.670 ;
        RECT 1030.930 3197.090 1032.110 3198.270 ;
        RECT 1030.930 3195.490 1032.110 3196.670 ;
        RECT 1030.930 3017.090 1032.110 3018.270 ;
        RECT 1030.930 3015.490 1032.110 3016.670 ;
        RECT 1030.930 2837.090 1032.110 2838.270 ;
        RECT 1030.930 2835.490 1032.110 2836.670 ;
        RECT 1030.930 2657.090 1032.110 2658.270 ;
        RECT 1030.930 2655.490 1032.110 2656.670 ;
        RECT 1030.930 2477.090 1032.110 2478.270 ;
        RECT 1030.930 2475.490 1032.110 2476.670 ;
        RECT 1030.930 2297.090 1032.110 2298.270 ;
        RECT 1030.930 2295.490 1032.110 2296.670 ;
        RECT 1030.930 2117.090 1032.110 2118.270 ;
        RECT 1030.930 2115.490 1032.110 2116.670 ;
        RECT 1030.930 1937.090 1032.110 1938.270 ;
        RECT 1030.930 1935.490 1032.110 1936.670 ;
        RECT 1030.930 1757.090 1032.110 1758.270 ;
        RECT 1030.930 1755.490 1032.110 1756.670 ;
        RECT 1030.930 1577.090 1032.110 1578.270 ;
        RECT 1030.930 1575.490 1032.110 1576.670 ;
        RECT 1030.930 1397.090 1032.110 1398.270 ;
        RECT 1030.930 1395.490 1032.110 1396.670 ;
        RECT 1030.930 1217.090 1032.110 1218.270 ;
        RECT 1030.930 1215.490 1032.110 1216.670 ;
        RECT 1030.930 1037.090 1032.110 1038.270 ;
        RECT 1030.930 1035.490 1032.110 1036.670 ;
        RECT 1030.930 857.090 1032.110 858.270 ;
        RECT 1030.930 855.490 1032.110 856.670 ;
        RECT 1030.930 677.090 1032.110 678.270 ;
        RECT 1030.930 675.490 1032.110 676.670 ;
        RECT 1030.930 497.090 1032.110 498.270 ;
        RECT 1030.930 495.490 1032.110 496.670 ;
        RECT 1030.930 317.090 1032.110 318.270 ;
        RECT 1030.930 315.490 1032.110 316.670 ;
        RECT 1030.930 137.090 1032.110 138.270 ;
        RECT 1030.930 135.490 1032.110 136.670 ;
        RECT 1030.930 -25.910 1032.110 -24.730 ;
        RECT 1030.930 -27.510 1032.110 -26.330 ;
        RECT 1210.930 3546.010 1212.110 3547.190 ;
        RECT 1210.930 3544.410 1212.110 3545.590 ;
        RECT 1210.930 3377.090 1212.110 3378.270 ;
        RECT 1210.930 3375.490 1212.110 3376.670 ;
        RECT 1210.930 3197.090 1212.110 3198.270 ;
        RECT 1210.930 3195.490 1212.110 3196.670 ;
        RECT 1210.930 3017.090 1212.110 3018.270 ;
        RECT 1210.930 3015.490 1212.110 3016.670 ;
        RECT 1210.930 2837.090 1212.110 2838.270 ;
        RECT 1210.930 2835.490 1212.110 2836.670 ;
        RECT 1210.930 2657.090 1212.110 2658.270 ;
        RECT 1210.930 2655.490 1212.110 2656.670 ;
        RECT 1210.930 2477.090 1212.110 2478.270 ;
        RECT 1210.930 2475.490 1212.110 2476.670 ;
        RECT 1210.930 2297.090 1212.110 2298.270 ;
        RECT 1210.930 2295.490 1212.110 2296.670 ;
        RECT 1210.930 2117.090 1212.110 2118.270 ;
        RECT 1210.930 2115.490 1212.110 2116.670 ;
        RECT 1210.930 1937.090 1212.110 1938.270 ;
        RECT 1210.930 1935.490 1212.110 1936.670 ;
        RECT 1210.930 1757.090 1212.110 1758.270 ;
        RECT 1210.930 1755.490 1212.110 1756.670 ;
        RECT 1210.930 1577.090 1212.110 1578.270 ;
        RECT 1210.930 1575.490 1212.110 1576.670 ;
        RECT 1210.930 1397.090 1212.110 1398.270 ;
        RECT 1210.930 1395.490 1212.110 1396.670 ;
        RECT 1210.930 1217.090 1212.110 1218.270 ;
        RECT 1210.930 1215.490 1212.110 1216.670 ;
        RECT 1210.930 1037.090 1212.110 1038.270 ;
        RECT 1210.930 1035.490 1212.110 1036.670 ;
        RECT 1210.930 857.090 1212.110 858.270 ;
        RECT 1210.930 855.490 1212.110 856.670 ;
        RECT 1210.930 677.090 1212.110 678.270 ;
        RECT 1210.930 675.490 1212.110 676.670 ;
        RECT 1210.930 497.090 1212.110 498.270 ;
        RECT 1210.930 495.490 1212.110 496.670 ;
        RECT 1210.930 317.090 1212.110 318.270 ;
        RECT 1210.930 315.490 1212.110 316.670 ;
        RECT 1210.930 137.090 1212.110 138.270 ;
        RECT 1210.930 135.490 1212.110 136.670 ;
        RECT 1210.930 -25.910 1212.110 -24.730 ;
        RECT 1210.930 -27.510 1212.110 -26.330 ;
        RECT 1390.930 3546.010 1392.110 3547.190 ;
        RECT 1390.930 3544.410 1392.110 3545.590 ;
        RECT 1390.930 3377.090 1392.110 3378.270 ;
        RECT 1390.930 3375.490 1392.110 3376.670 ;
        RECT 1390.930 3197.090 1392.110 3198.270 ;
        RECT 1390.930 3195.490 1392.110 3196.670 ;
        RECT 1390.930 3017.090 1392.110 3018.270 ;
        RECT 1390.930 3015.490 1392.110 3016.670 ;
        RECT 1390.930 2837.090 1392.110 2838.270 ;
        RECT 1390.930 2835.490 1392.110 2836.670 ;
        RECT 1390.930 2657.090 1392.110 2658.270 ;
        RECT 1390.930 2655.490 1392.110 2656.670 ;
        RECT 1390.930 2477.090 1392.110 2478.270 ;
        RECT 1390.930 2475.490 1392.110 2476.670 ;
        RECT 1390.930 2297.090 1392.110 2298.270 ;
        RECT 1390.930 2295.490 1392.110 2296.670 ;
        RECT 1390.930 2117.090 1392.110 2118.270 ;
        RECT 1390.930 2115.490 1392.110 2116.670 ;
        RECT 1390.930 1937.090 1392.110 1938.270 ;
        RECT 1390.930 1935.490 1392.110 1936.670 ;
        RECT 1390.930 1757.090 1392.110 1758.270 ;
        RECT 1390.930 1755.490 1392.110 1756.670 ;
        RECT 1390.930 1577.090 1392.110 1578.270 ;
        RECT 1390.930 1575.490 1392.110 1576.670 ;
        RECT 1390.930 1397.090 1392.110 1398.270 ;
        RECT 1390.930 1395.490 1392.110 1396.670 ;
        RECT 1390.930 1217.090 1392.110 1218.270 ;
        RECT 1390.930 1215.490 1392.110 1216.670 ;
        RECT 1390.930 1037.090 1392.110 1038.270 ;
        RECT 1390.930 1035.490 1392.110 1036.670 ;
        RECT 1390.930 857.090 1392.110 858.270 ;
        RECT 1390.930 855.490 1392.110 856.670 ;
        RECT 1390.930 677.090 1392.110 678.270 ;
        RECT 1390.930 675.490 1392.110 676.670 ;
        RECT 1390.930 497.090 1392.110 498.270 ;
        RECT 1390.930 495.490 1392.110 496.670 ;
        RECT 1390.930 317.090 1392.110 318.270 ;
        RECT 1390.930 315.490 1392.110 316.670 ;
        RECT 1390.930 137.090 1392.110 138.270 ;
        RECT 1390.930 135.490 1392.110 136.670 ;
        RECT 1390.930 -25.910 1392.110 -24.730 ;
        RECT 1390.930 -27.510 1392.110 -26.330 ;
        RECT 1570.930 3546.010 1572.110 3547.190 ;
        RECT 1570.930 3544.410 1572.110 3545.590 ;
        RECT 1570.930 3377.090 1572.110 3378.270 ;
        RECT 1570.930 3375.490 1572.110 3376.670 ;
        RECT 1570.930 3197.090 1572.110 3198.270 ;
        RECT 1570.930 3195.490 1572.110 3196.670 ;
        RECT 1570.930 3017.090 1572.110 3018.270 ;
        RECT 1570.930 3015.490 1572.110 3016.670 ;
        RECT 1570.930 2837.090 1572.110 2838.270 ;
        RECT 1570.930 2835.490 1572.110 2836.670 ;
        RECT 1570.930 2657.090 1572.110 2658.270 ;
        RECT 1570.930 2655.490 1572.110 2656.670 ;
        RECT 1570.930 2477.090 1572.110 2478.270 ;
        RECT 1570.930 2475.490 1572.110 2476.670 ;
        RECT 1570.930 2297.090 1572.110 2298.270 ;
        RECT 1570.930 2295.490 1572.110 2296.670 ;
        RECT 1570.930 2117.090 1572.110 2118.270 ;
        RECT 1570.930 2115.490 1572.110 2116.670 ;
        RECT 1570.930 1937.090 1572.110 1938.270 ;
        RECT 1570.930 1935.490 1572.110 1936.670 ;
        RECT 1570.930 1757.090 1572.110 1758.270 ;
        RECT 1570.930 1755.490 1572.110 1756.670 ;
        RECT 1570.930 1577.090 1572.110 1578.270 ;
        RECT 1570.930 1575.490 1572.110 1576.670 ;
        RECT 1570.930 1397.090 1572.110 1398.270 ;
        RECT 1570.930 1395.490 1572.110 1396.670 ;
        RECT 1570.930 1217.090 1572.110 1218.270 ;
        RECT 1570.930 1215.490 1572.110 1216.670 ;
        RECT 1570.930 1037.090 1572.110 1038.270 ;
        RECT 1570.930 1035.490 1572.110 1036.670 ;
        RECT 1570.930 857.090 1572.110 858.270 ;
        RECT 1570.930 855.490 1572.110 856.670 ;
        RECT 1570.930 677.090 1572.110 678.270 ;
        RECT 1570.930 675.490 1572.110 676.670 ;
        RECT 1570.930 497.090 1572.110 498.270 ;
        RECT 1570.930 495.490 1572.110 496.670 ;
        RECT 1570.930 317.090 1572.110 318.270 ;
        RECT 1570.930 315.490 1572.110 316.670 ;
        RECT 1570.930 137.090 1572.110 138.270 ;
        RECT 1570.930 135.490 1572.110 136.670 ;
        RECT 1570.930 -25.910 1572.110 -24.730 ;
        RECT 1570.930 -27.510 1572.110 -26.330 ;
        RECT 1750.930 3546.010 1752.110 3547.190 ;
        RECT 1750.930 3544.410 1752.110 3545.590 ;
        RECT 1750.930 3377.090 1752.110 3378.270 ;
        RECT 1750.930 3375.490 1752.110 3376.670 ;
        RECT 1750.930 3197.090 1752.110 3198.270 ;
        RECT 1750.930 3195.490 1752.110 3196.670 ;
        RECT 1750.930 3017.090 1752.110 3018.270 ;
        RECT 1750.930 3015.490 1752.110 3016.670 ;
        RECT 1750.930 2837.090 1752.110 2838.270 ;
        RECT 1750.930 2835.490 1752.110 2836.670 ;
        RECT 1750.930 2657.090 1752.110 2658.270 ;
        RECT 1750.930 2655.490 1752.110 2656.670 ;
        RECT 1750.930 2477.090 1752.110 2478.270 ;
        RECT 1750.930 2475.490 1752.110 2476.670 ;
        RECT 1750.930 2297.090 1752.110 2298.270 ;
        RECT 1750.930 2295.490 1752.110 2296.670 ;
        RECT 1750.930 2117.090 1752.110 2118.270 ;
        RECT 1750.930 2115.490 1752.110 2116.670 ;
        RECT 1750.930 1937.090 1752.110 1938.270 ;
        RECT 1750.930 1935.490 1752.110 1936.670 ;
        RECT 1750.930 1757.090 1752.110 1758.270 ;
        RECT 1750.930 1755.490 1752.110 1756.670 ;
        RECT 1750.930 1577.090 1752.110 1578.270 ;
        RECT 1750.930 1575.490 1752.110 1576.670 ;
        RECT 1750.930 1397.090 1752.110 1398.270 ;
        RECT 1750.930 1395.490 1752.110 1396.670 ;
        RECT 1750.930 1217.090 1752.110 1218.270 ;
        RECT 1750.930 1215.490 1752.110 1216.670 ;
        RECT 1750.930 1037.090 1752.110 1038.270 ;
        RECT 1750.930 1035.490 1752.110 1036.670 ;
        RECT 1750.930 857.090 1752.110 858.270 ;
        RECT 1750.930 855.490 1752.110 856.670 ;
        RECT 1750.930 677.090 1752.110 678.270 ;
        RECT 1750.930 675.490 1752.110 676.670 ;
        RECT 1750.930 497.090 1752.110 498.270 ;
        RECT 1750.930 495.490 1752.110 496.670 ;
        RECT 1750.930 317.090 1752.110 318.270 ;
        RECT 1750.930 315.490 1752.110 316.670 ;
        RECT 1750.930 137.090 1752.110 138.270 ;
        RECT 1750.930 135.490 1752.110 136.670 ;
        RECT 1750.930 -25.910 1752.110 -24.730 ;
        RECT 1750.930 -27.510 1752.110 -26.330 ;
        RECT 1930.930 3546.010 1932.110 3547.190 ;
        RECT 1930.930 3544.410 1932.110 3545.590 ;
        RECT 1930.930 3377.090 1932.110 3378.270 ;
        RECT 1930.930 3375.490 1932.110 3376.670 ;
        RECT 1930.930 3197.090 1932.110 3198.270 ;
        RECT 1930.930 3195.490 1932.110 3196.670 ;
        RECT 1930.930 3017.090 1932.110 3018.270 ;
        RECT 1930.930 3015.490 1932.110 3016.670 ;
        RECT 1930.930 2837.090 1932.110 2838.270 ;
        RECT 1930.930 2835.490 1932.110 2836.670 ;
        RECT 1930.930 2657.090 1932.110 2658.270 ;
        RECT 1930.930 2655.490 1932.110 2656.670 ;
        RECT 1930.930 2477.090 1932.110 2478.270 ;
        RECT 1930.930 2475.490 1932.110 2476.670 ;
        RECT 1930.930 2297.090 1932.110 2298.270 ;
        RECT 1930.930 2295.490 1932.110 2296.670 ;
        RECT 1930.930 2117.090 1932.110 2118.270 ;
        RECT 1930.930 2115.490 1932.110 2116.670 ;
        RECT 1930.930 1937.090 1932.110 1938.270 ;
        RECT 1930.930 1935.490 1932.110 1936.670 ;
        RECT 1930.930 1757.090 1932.110 1758.270 ;
        RECT 1930.930 1755.490 1932.110 1756.670 ;
        RECT 1930.930 1577.090 1932.110 1578.270 ;
        RECT 1930.930 1575.490 1932.110 1576.670 ;
        RECT 1930.930 1397.090 1932.110 1398.270 ;
        RECT 1930.930 1395.490 1932.110 1396.670 ;
        RECT 1930.930 1217.090 1932.110 1218.270 ;
        RECT 1930.930 1215.490 1932.110 1216.670 ;
        RECT 1930.930 1037.090 1932.110 1038.270 ;
        RECT 1930.930 1035.490 1932.110 1036.670 ;
        RECT 1930.930 857.090 1932.110 858.270 ;
        RECT 1930.930 855.490 1932.110 856.670 ;
        RECT 1930.930 677.090 1932.110 678.270 ;
        RECT 1930.930 675.490 1932.110 676.670 ;
        RECT 1930.930 497.090 1932.110 498.270 ;
        RECT 1930.930 495.490 1932.110 496.670 ;
        RECT 1930.930 317.090 1932.110 318.270 ;
        RECT 1930.930 315.490 1932.110 316.670 ;
        RECT 1930.930 137.090 1932.110 138.270 ;
        RECT 1930.930 135.490 1932.110 136.670 ;
        RECT 1930.930 -25.910 1932.110 -24.730 ;
        RECT 1930.930 -27.510 1932.110 -26.330 ;
        RECT 2110.930 3546.010 2112.110 3547.190 ;
        RECT 2110.930 3544.410 2112.110 3545.590 ;
        RECT 2110.930 3377.090 2112.110 3378.270 ;
        RECT 2110.930 3375.490 2112.110 3376.670 ;
        RECT 2110.930 3197.090 2112.110 3198.270 ;
        RECT 2110.930 3195.490 2112.110 3196.670 ;
        RECT 2110.930 3017.090 2112.110 3018.270 ;
        RECT 2110.930 3015.490 2112.110 3016.670 ;
        RECT 2110.930 2837.090 2112.110 2838.270 ;
        RECT 2110.930 2835.490 2112.110 2836.670 ;
        RECT 2110.930 2657.090 2112.110 2658.270 ;
        RECT 2110.930 2655.490 2112.110 2656.670 ;
        RECT 2110.930 2477.090 2112.110 2478.270 ;
        RECT 2110.930 2475.490 2112.110 2476.670 ;
        RECT 2110.930 2297.090 2112.110 2298.270 ;
        RECT 2110.930 2295.490 2112.110 2296.670 ;
        RECT 2110.930 2117.090 2112.110 2118.270 ;
        RECT 2110.930 2115.490 2112.110 2116.670 ;
        RECT 2110.930 1937.090 2112.110 1938.270 ;
        RECT 2110.930 1935.490 2112.110 1936.670 ;
        RECT 2110.930 1757.090 2112.110 1758.270 ;
        RECT 2110.930 1755.490 2112.110 1756.670 ;
        RECT 2110.930 1577.090 2112.110 1578.270 ;
        RECT 2110.930 1575.490 2112.110 1576.670 ;
        RECT 2110.930 1397.090 2112.110 1398.270 ;
        RECT 2110.930 1395.490 2112.110 1396.670 ;
        RECT 2110.930 1217.090 2112.110 1218.270 ;
        RECT 2110.930 1215.490 2112.110 1216.670 ;
        RECT 2110.930 1037.090 2112.110 1038.270 ;
        RECT 2110.930 1035.490 2112.110 1036.670 ;
        RECT 2110.930 857.090 2112.110 858.270 ;
        RECT 2110.930 855.490 2112.110 856.670 ;
        RECT 2110.930 677.090 2112.110 678.270 ;
        RECT 2110.930 675.490 2112.110 676.670 ;
        RECT 2110.930 497.090 2112.110 498.270 ;
        RECT 2110.930 495.490 2112.110 496.670 ;
        RECT 2110.930 317.090 2112.110 318.270 ;
        RECT 2110.930 315.490 2112.110 316.670 ;
        RECT 2110.930 137.090 2112.110 138.270 ;
        RECT 2110.930 135.490 2112.110 136.670 ;
        RECT 2110.930 -25.910 2112.110 -24.730 ;
        RECT 2110.930 -27.510 2112.110 -26.330 ;
        RECT 2290.930 3546.010 2292.110 3547.190 ;
        RECT 2290.930 3544.410 2292.110 3545.590 ;
        RECT 2290.930 3377.090 2292.110 3378.270 ;
        RECT 2290.930 3375.490 2292.110 3376.670 ;
        RECT 2290.930 3197.090 2292.110 3198.270 ;
        RECT 2290.930 3195.490 2292.110 3196.670 ;
        RECT 2290.930 3017.090 2292.110 3018.270 ;
        RECT 2290.930 3015.490 2292.110 3016.670 ;
        RECT 2290.930 2837.090 2292.110 2838.270 ;
        RECT 2290.930 2835.490 2292.110 2836.670 ;
        RECT 2290.930 2657.090 2292.110 2658.270 ;
        RECT 2290.930 2655.490 2292.110 2656.670 ;
        RECT 2290.930 2477.090 2292.110 2478.270 ;
        RECT 2290.930 2475.490 2292.110 2476.670 ;
        RECT 2290.930 2297.090 2292.110 2298.270 ;
        RECT 2290.930 2295.490 2292.110 2296.670 ;
        RECT 2290.930 2117.090 2292.110 2118.270 ;
        RECT 2290.930 2115.490 2292.110 2116.670 ;
        RECT 2290.930 1937.090 2292.110 1938.270 ;
        RECT 2290.930 1935.490 2292.110 1936.670 ;
        RECT 2290.930 1757.090 2292.110 1758.270 ;
        RECT 2290.930 1755.490 2292.110 1756.670 ;
        RECT 2290.930 1577.090 2292.110 1578.270 ;
        RECT 2290.930 1575.490 2292.110 1576.670 ;
        RECT 2290.930 1397.090 2292.110 1398.270 ;
        RECT 2290.930 1395.490 2292.110 1396.670 ;
        RECT 2290.930 1217.090 2292.110 1218.270 ;
        RECT 2290.930 1215.490 2292.110 1216.670 ;
        RECT 2290.930 1037.090 2292.110 1038.270 ;
        RECT 2290.930 1035.490 2292.110 1036.670 ;
        RECT 2290.930 857.090 2292.110 858.270 ;
        RECT 2290.930 855.490 2292.110 856.670 ;
        RECT 2290.930 677.090 2292.110 678.270 ;
        RECT 2290.930 675.490 2292.110 676.670 ;
        RECT 2290.930 497.090 2292.110 498.270 ;
        RECT 2290.930 495.490 2292.110 496.670 ;
        RECT 2290.930 317.090 2292.110 318.270 ;
        RECT 2290.930 315.490 2292.110 316.670 ;
        RECT 2290.930 137.090 2292.110 138.270 ;
        RECT 2290.930 135.490 2292.110 136.670 ;
        RECT 2290.930 -25.910 2292.110 -24.730 ;
        RECT 2290.930 -27.510 2292.110 -26.330 ;
        RECT 2470.930 3546.010 2472.110 3547.190 ;
        RECT 2470.930 3544.410 2472.110 3545.590 ;
        RECT 2470.930 3377.090 2472.110 3378.270 ;
        RECT 2470.930 3375.490 2472.110 3376.670 ;
        RECT 2470.930 3197.090 2472.110 3198.270 ;
        RECT 2470.930 3195.490 2472.110 3196.670 ;
        RECT 2470.930 3017.090 2472.110 3018.270 ;
        RECT 2470.930 3015.490 2472.110 3016.670 ;
        RECT 2470.930 2837.090 2472.110 2838.270 ;
        RECT 2470.930 2835.490 2472.110 2836.670 ;
        RECT 2470.930 2657.090 2472.110 2658.270 ;
        RECT 2470.930 2655.490 2472.110 2656.670 ;
        RECT 2470.930 2477.090 2472.110 2478.270 ;
        RECT 2470.930 2475.490 2472.110 2476.670 ;
        RECT 2470.930 2297.090 2472.110 2298.270 ;
        RECT 2470.930 2295.490 2472.110 2296.670 ;
        RECT 2470.930 2117.090 2472.110 2118.270 ;
        RECT 2470.930 2115.490 2472.110 2116.670 ;
        RECT 2470.930 1937.090 2472.110 1938.270 ;
        RECT 2470.930 1935.490 2472.110 1936.670 ;
        RECT 2470.930 1757.090 2472.110 1758.270 ;
        RECT 2470.930 1755.490 2472.110 1756.670 ;
        RECT 2470.930 1577.090 2472.110 1578.270 ;
        RECT 2470.930 1575.490 2472.110 1576.670 ;
        RECT 2470.930 1397.090 2472.110 1398.270 ;
        RECT 2470.930 1395.490 2472.110 1396.670 ;
        RECT 2470.930 1217.090 2472.110 1218.270 ;
        RECT 2470.930 1215.490 2472.110 1216.670 ;
        RECT 2470.930 1037.090 2472.110 1038.270 ;
        RECT 2470.930 1035.490 2472.110 1036.670 ;
        RECT 2470.930 857.090 2472.110 858.270 ;
        RECT 2470.930 855.490 2472.110 856.670 ;
        RECT 2470.930 677.090 2472.110 678.270 ;
        RECT 2470.930 675.490 2472.110 676.670 ;
        RECT 2470.930 497.090 2472.110 498.270 ;
        RECT 2470.930 495.490 2472.110 496.670 ;
        RECT 2470.930 317.090 2472.110 318.270 ;
        RECT 2470.930 315.490 2472.110 316.670 ;
        RECT 2470.930 137.090 2472.110 138.270 ;
        RECT 2470.930 135.490 2472.110 136.670 ;
        RECT 2470.930 -25.910 2472.110 -24.730 ;
        RECT 2470.930 -27.510 2472.110 -26.330 ;
        RECT 2650.930 3546.010 2652.110 3547.190 ;
        RECT 2650.930 3544.410 2652.110 3545.590 ;
        RECT 2650.930 3377.090 2652.110 3378.270 ;
        RECT 2650.930 3375.490 2652.110 3376.670 ;
        RECT 2650.930 3197.090 2652.110 3198.270 ;
        RECT 2650.930 3195.490 2652.110 3196.670 ;
        RECT 2650.930 3017.090 2652.110 3018.270 ;
        RECT 2650.930 3015.490 2652.110 3016.670 ;
        RECT 2650.930 2837.090 2652.110 2838.270 ;
        RECT 2650.930 2835.490 2652.110 2836.670 ;
        RECT 2650.930 2657.090 2652.110 2658.270 ;
        RECT 2650.930 2655.490 2652.110 2656.670 ;
        RECT 2650.930 2477.090 2652.110 2478.270 ;
        RECT 2650.930 2475.490 2652.110 2476.670 ;
        RECT 2650.930 2297.090 2652.110 2298.270 ;
        RECT 2650.930 2295.490 2652.110 2296.670 ;
        RECT 2650.930 2117.090 2652.110 2118.270 ;
        RECT 2650.930 2115.490 2652.110 2116.670 ;
        RECT 2650.930 1937.090 2652.110 1938.270 ;
        RECT 2650.930 1935.490 2652.110 1936.670 ;
        RECT 2650.930 1757.090 2652.110 1758.270 ;
        RECT 2650.930 1755.490 2652.110 1756.670 ;
        RECT 2650.930 1577.090 2652.110 1578.270 ;
        RECT 2650.930 1575.490 2652.110 1576.670 ;
        RECT 2650.930 1397.090 2652.110 1398.270 ;
        RECT 2650.930 1395.490 2652.110 1396.670 ;
        RECT 2650.930 1217.090 2652.110 1218.270 ;
        RECT 2650.930 1215.490 2652.110 1216.670 ;
        RECT 2650.930 1037.090 2652.110 1038.270 ;
        RECT 2650.930 1035.490 2652.110 1036.670 ;
        RECT 2650.930 857.090 2652.110 858.270 ;
        RECT 2650.930 855.490 2652.110 856.670 ;
        RECT 2650.930 677.090 2652.110 678.270 ;
        RECT 2650.930 675.490 2652.110 676.670 ;
        RECT 2650.930 497.090 2652.110 498.270 ;
        RECT 2650.930 495.490 2652.110 496.670 ;
        RECT 2650.930 317.090 2652.110 318.270 ;
        RECT 2650.930 315.490 2652.110 316.670 ;
        RECT 2650.930 137.090 2652.110 138.270 ;
        RECT 2650.930 135.490 2652.110 136.670 ;
        RECT 2650.930 -25.910 2652.110 -24.730 ;
        RECT 2650.930 -27.510 2652.110 -26.330 ;
        RECT 2830.930 3546.010 2832.110 3547.190 ;
        RECT 2830.930 3544.410 2832.110 3545.590 ;
        RECT 2830.930 3377.090 2832.110 3378.270 ;
        RECT 2830.930 3375.490 2832.110 3376.670 ;
        RECT 2830.930 3197.090 2832.110 3198.270 ;
        RECT 2830.930 3195.490 2832.110 3196.670 ;
        RECT 2830.930 3017.090 2832.110 3018.270 ;
        RECT 2830.930 3015.490 2832.110 3016.670 ;
        RECT 2830.930 2837.090 2832.110 2838.270 ;
        RECT 2830.930 2835.490 2832.110 2836.670 ;
        RECT 2830.930 2657.090 2832.110 2658.270 ;
        RECT 2830.930 2655.490 2832.110 2656.670 ;
        RECT 2830.930 2477.090 2832.110 2478.270 ;
        RECT 2830.930 2475.490 2832.110 2476.670 ;
        RECT 2830.930 2297.090 2832.110 2298.270 ;
        RECT 2830.930 2295.490 2832.110 2296.670 ;
        RECT 2830.930 2117.090 2832.110 2118.270 ;
        RECT 2830.930 2115.490 2832.110 2116.670 ;
        RECT 2830.930 1937.090 2832.110 1938.270 ;
        RECT 2830.930 1935.490 2832.110 1936.670 ;
        RECT 2830.930 1757.090 2832.110 1758.270 ;
        RECT 2830.930 1755.490 2832.110 1756.670 ;
        RECT 2830.930 1577.090 2832.110 1578.270 ;
        RECT 2830.930 1575.490 2832.110 1576.670 ;
        RECT 2830.930 1397.090 2832.110 1398.270 ;
        RECT 2830.930 1395.490 2832.110 1396.670 ;
        RECT 2830.930 1217.090 2832.110 1218.270 ;
        RECT 2830.930 1215.490 2832.110 1216.670 ;
        RECT 2830.930 1037.090 2832.110 1038.270 ;
        RECT 2830.930 1035.490 2832.110 1036.670 ;
        RECT 2830.930 857.090 2832.110 858.270 ;
        RECT 2830.930 855.490 2832.110 856.670 ;
        RECT 2830.930 677.090 2832.110 678.270 ;
        RECT 2830.930 675.490 2832.110 676.670 ;
        RECT 2830.930 497.090 2832.110 498.270 ;
        RECT 2830.930 495.490 2832.110 496.670 ;
        RECT 2830.930 317.090 2832.110 318.270 ;
        RECT 2830.930 315.490 2832.110 316.670 ;
        RECT 2830.930 137.090 2832.110 138.270 ;
        RECT 2830.930 135.490 2832.110 136.670 ;
        RECT 2830.930 -25.910 2832.110 -24.730 ;
        RECT 2830.930 -27.510 2832.110 -26.330 ;
        RECT 2950.510 3546.010 2951.690 3547.190 ;
        RECT 2950.510 3544.410 2951.690 3545.590 ;
        RECT 2950.510 3377.090 2951.690 3378.270 ;
        RECT 2950.510 3375.490 2951.690 3376.670 ;
        RECT 2950.510 3197.090 2951.690 3198.270 ;
        RECT 2950.510 3195.490 2951.690 3196.670 ;
        RECT 2950.510 3017.090 2951.690 3018.270 ;
        RECT 2950.510 3015.490 2951.690 3016.670 ;
        RECT 2950.510 2837.090 2951.690 2838.270 ;
        RECT 2950.510 2835.490 2951.690 2836.670 ;
        RECT 2950.510 2657.090 2951.690 2658.270 ;
        RECT 2950.510 2655.490 2951.690 2656.670 ;
        RECT 2950.510 2477.090 2951.690 2478.270 ;
        RECT 2950.510 2475.490 2951.690 2476.670 ;
        RECT 2950.510 2297.090 2951.690 2298.270 ;
        RECT 2950.510 2295.490 2951.690 2296.670 ;
        RECT 2950.510 2117.090 2951.690 2118.270 ;
        RECT 2950.510 2115.490 2951.690 2116.670 ;
        RECT 2950.510 1937.090 2951.690 1938.270 ;
        RECT 2950.510 1935.490 2951.690 1936.670 ;
        RECT 2950.510 1757.090 2951.690 1758.270 ;
        RECT 2950.510 1755.490 2951.690 1756.670 ;
        RECT 2950.510 1577.090 2951.690 1578.270 ;
        RECT 2950.510 1575.490 2951.690 1576.670 ;
        RECT 2950.510 1397.090 2951.690 1398.270 ;
        RECT 2950.510 1395.490 2951.690 1396.670 ;
        RECT 2950.510 1217.090 2951.690 1218.270 ;
        RECT 2950.510 1215.490 2951.690 1216.670 ;
        RECT 2950.510 1037.090 2951.690 1038.270 ;
        RECT 2950.510 1035.490 2951.690 1036.670 ;
        RECT 2950.510 857.090 2951.690 858.270 ;
        RECT 2950.510 855.490 2951.690 856.670 ;
        RECT 2950.510 677.090 2951.690 678.270 ;
        RECT 2950.510 675.490 2951.690 676.670 ;
        RECT 2950.510 497.090 2951.690 498.270 ;
        RECT 2950.510 495.490 2951.690 496.670 ;
        RECT 2950.510 317.090 2951.690 318.270 ;
        RECT 2950.510 315.490 2951.690 316.670 ;
        RECT 2950.510 137.090 2951.690 138.270 ;
        RECT 2950.510 135.490 2951.690 136.670 ;
        RECT 2950.510 -25.910 2951.690 -24.730 ;
        RECT 2950.510 -27.510 2951.690 -26.330 ;
      LAYER met5 ;
        RECT -32.980 3547.300 -29.980 3547.310 ;
        RECT 130.020 3547.300 133.020 3547.310 ;
        RECT 310.020 3547.300 313.020 3547.310 ;
        RECT 490.020 3547.300 493.020 3547.310 ;
        RECT 670.020 3547.300 673.020 3547.310 ;
        RECT 850.020 3547.300 853.020 3547.310 ;
        RECT 1030.020 3547.300 1033.020 3547.310 ;
        RECT 1210.020 3547.300 1213.020 3547.310 ;
        RECT 1390.020 3547.300 1393.020 3547.310 ;
        RECT 1570.020 3547.300 1573.020 3547.310 ;
        RECT 1750.020 3547.300 1753.020 3547.310 ;
        RECT 1930.020 3547.300 1933.020 3547.310 ;
        RECT 2110.020 3547.300 2113.020 3547.310 ;
        RECT 2290.020 3547.300 2293.020 3547.310 ;
        RECT 2470.020 3547.300 2473.020 3547.310 ;
        RECT 2650.020 3547.300 2653.020 3547.310 ;
        RECT 2830.020 3547.300 2833.020 3547.310 ;
        RECT 2949.600 3547.300 2952.600 3547.310 ;
        RECT -32.980 3544.300 2952.600 3547.300 ;
        RECT -32.980 3544.290 -29.980 3544.300 ;
        RECT 130.020 3544.290 133.020 3544.300 ;
        RECT 310.020 3544.290 313.020 3544.300 ;
        RECT 490.020 3544.290 493.020 3544.300 ;
        RECT 670.020 3544.290 673.020 3544.300 ;
        RECT 850.020 3544.290 853.020 3544.300 ;
        RECT 1030.020 3544.290 1033.020 3544.300 ;
        RECT 1210.020 3544.290 1213.020 3544.300 ;
        RECT 1390.020 3544.290 1393.020 3544.300 ;
        RECT 1570.020 3544.290 1573.020 3544.300 ;
        RECT 1750.020 3544.290 1753.020 3544.300 ;
        RECT 1930.020 3544.290 1933.020 3544.300 ;
        RECT 2110.020 3544.290 2113.020 3544.300 ;
        RECT 2290.020 3544.290 2293.020 3544.300 ;
        RECT 2470.020 3544.290 2473.020 3544.300 ;
        RECT 2650.020 3544.290 2653.020 3544.300 ;
        RECT 2830.020 3544.290 2833.020 3544.300 ;
        RECT 2949.600 3544.290 2952.600 3544.300 ;
        RECT -32.980 3378.380 -29.980 3378.390 ;
        RECT 130.020 3378.380 133.020 3378.390 ;
        RECT 310.020 3378.380 313.020 3378.390 ;
        RECT 490.020 3378.380 493.020 3378.390 ;
        RECT 670.020 3378.380 673.020 3378.390 ;
        RECT 850.020 3378.380 853.020 3378.390 ;
        RECT 1030.020 3378.380 1033.020 3378.390 ;
        RECT 1210.020 3378.380 1213.020 3378.390 ;
        RECT 1390.020 3378.380 1393.020 3378.390 ;
        RECT 1570.020 3378.380 1573.020 3378.390 ;
        RECT 1750.020 3378.380 1753.020 3378.390 ;
        RECT 1930.020 3378.380 1933.020 3378.390 ;
        RECT 2110.020 3378.380 2113.020 3378.390 ;
        RECT 2290.020 3378.380 2293.020 3378.390 ;
        RECT 2470.020 3378.380 2473.020 3378.390 ;
        RECT 2650.020 3378.380 2653.020 3378.390 ;
        RECT 2830.020 3378.380 2833.020 3378.390 ;
        RECT 2949.600 3378.380 2952.600 3378.390 ;
        RECT -32.980 3375.380 2952.600 3378.380 ;
        RECT -32.980 3375.370 -29.980 3375.380 ;
        RECT 130.020 3375.370 133.020 3375.380 ;
        RECT 310.020 3375.370 313.020 3375.380 ;
        RECT 490.020 3375.370 493.020 3375.380 ;
        RECT 670.020 3375.370 673.020 3375.380 ;
        RECT 850.020 3375.370 853.020 3375.380 ;
        RECT 1030.020 3375.370 1033.020 3375.380 ;
        RECT 1210.020 3375.370 1213.020 3375.380 ;
        RECT 1390.020 3375.370 1393.020 3375.380 ;
        RECT 1570.020 3375.370 1573.020 3375.380 ;
        RECT 1750.020 3375.370 1753.020 3375.380 ;
        RECT 1930.020 3375.370 1933.020 3375.380 ;
        RECT 2110.020 3375.370 2113.020 3375.380 ;
        RECT 2290.020 3375.370 2293.020 3375.380 ;
        RECT 2470.020 3375.370 2473.020 3375.380 ;
        RECT 2650.020 3375.370 2653.020 3375.380 ;
        RECT 2830.020 3375.370 2833.020 3375.380 ;
        RECT 2949.600 3375.370 2952.600 3375.380 ;
        RECT -32.980 3198.380 -29.980 3198.390 ;
        RECT 130.020 3198.380 133.020 3198.390 ;
        RECT 310.020 3198.380 313.020 3198.390 ;
        RECT 490.020 3198.380 493.020 3198.390 ;
        RECT 670.020 3198.380 673.020 3198.390 ;
        RECT 850.020 3198.380 853.020 3198.390 ;
        RECT 1030.020 3198.380 1033.020 3198.390 ;
        RECT 1210.020 3198.380 1213.020 3198.390 ;
        RECT 1390.020 3198.380 1393.020 3198.390 ;
        RECT 1570.020 3198.380 1573.020 3198.390 ;
        RECT 1750.020 3198.380 1753.020 3198.390 ;
        RECT 1930.020 3198.380 1933.020 3198.390 ;
        RECT 2110.020 3198.380 2113.020 3198.390 ;
        RECT 2290.020 3198.380 2293.020 3198.390 ;
        RECT 2470.020 3198.380 2473.020 3198.390 ;
        RECT 2650.020 3198.380 2653.020 3198.390 ;
        RECT 2830.020 3198.380 2833.020 3198.390 ;
        RECT 2949.600 3198.380 2952.600 3198.390 ;
        RECT -32.980 3195.380 2952.600 3198.380 ;
        RECT -32.980 3195.370 -29.980 3195.380 ;
        RECT 130.020 3195.370 133.020 3195.380 ;
        RECT 310.020 3195.370 313.020 3195.380 ;
        RECT 490.020 3195.370 493.020 3195.380 ;
        RECT 670.020 3195.370 673.020 3195.380 ;
        RECT 850.020 3195.370 853.020 3195.380 ;
        RECT 1030.020 3195.370 1033.020 3195.380 ;
        RECT 1210.020 3195.370 1213.020 3195.380 ;
        RECT 1390.020 3195.370 1393.020 3195.380 ;
        RECT 1570.020 3195.370 1573.020 3195.380 ;
        RECT 1750.020 3195.370 1753.020 3195.380 ;
        RECT 1930.020 3195.370 1933.020 3195.380 ;
        RECT 2110.020 3195.370 2113.020 3195.380 ;
        RECT 2290.020 3195.370 2293.020 3195.380 ;
        RECT 2470.020 3195.370 2473.020 3195.380 ;
        RECT 2650.020 3195.370 2653.020 3195.380 ;
        RECT 2830.020 3195.370 2833.020 3195.380 ;
        RECT 2949.600 3195.370 2952.600 3195.380 ;
        RECT -32.980 3018.380 -29.980 3018.390 ;
        RECT 130.020 3018.380 133.020 3018.390 ;
        RECT 310.020 3018.380 313.020 3018.390 ;
        RECT 490.020 3018.380 493.020 3018.390 ;
        RECT 670.020 3018.380 673.020 3018.390 ;
        RECT 850.020 3018.380 853.020 3018.390 ;
        RECT 1030.020 3018.380 1033.020 3018.390 ;
        RECT 1210.020 3018.380 1213.020 3018.390 ;
        RECT 1390.020 3018.380 1393.020 3018.390 ;
        RECT 1570.020 3018.380 1573.020 3018.390 ;
        RECT 1750.020 3018.380 1753.020 3018.390 ;
        RECT 1930.020 3018.380 1933.020 3018.390 ;
        RECT 2110.020 3018.380 2113.020 3018.390 ;
        RECT 2290.020 3018.380 2293.020 3018.390 ;
        RECT 2470.020 3018.380 2473.020 3018.390 ;
        RECT 2650.020 3018.380 2653.020 3018.390 ;
        RECT 2830.020 3018.380 2833.020 3018.390 ;
        RECT 2949.600 3018.380 2952.600 3018.390 ;
        RECT -32.980 3015.380 2952.600 3018.380 ;
        RECT -32.980 3015.370 -29.980 3015.380 ;
        RECT 130.020 3015.370 133.020 3015.380 ;
        RECT 310.020 3015.370 313.020 3015.380 ;
        RECT 490.020 3015.370 493.020 3015.380 ;
        RECT 670.020 3015.370 673.020 3015.380 ;
        RECT 850.020 3015.370 853.020 3015.380 ;
        RECT 1030.020 3015.370 1033.020 3015.380 ;
        RECT 1210.020 3015.370 1213.020 3015.380 ;
        RECT 1390.020 3015.370 1393.020 3015.380 ;
        RECT 1570.020 3015.370 1573.020 3015.380 ;
        RECT 1750.020 3015.370 1753.020 3015.380 ;
        RECT 1930.020 3015.370 1933.020 3015.380 ;
        RECT 2110.020 3015.370 2113.020 3015.380 ;
        RECT 2290.020 3015.370 2293.020 3015.380 ;
        RECT 2470.020 3015.370 2473.020 3015.380 ;
        RECT 2650.020 3015.370 2653.020 3015.380 ;
        RECT 2830.020 3015.370 2833.020 3015.380 ;
        RECT 2949.600 3015.370 2952.600 3015.380 ;
        RECT -32.980 2838.380 -29.980 2838.390 ;
        RECT 130.020 2838.380 133.020 2838.390 ;
        RECT 310.020 2838.380 313.020 2838.390 ;
        RECT 490.020 2838.380 493.020 2838.390 ;
        RECT 670.020 2838.380 673.020 2838.390 ;
        RECT 850.020 2838.380 853.020 2838.390 ;
        RECT 1030.020 2838.380 1033.020 2838.390 ;
        RECT 1210.020 2838.380 1213.020 2838.390 ;
        RECT 1390.020 2838.380 1393.020 2838.390 ;
        RECT 1570.020 2838.380 1573.020 2838.390 ;
        RECT 1750.020 2838.380 1753.020 2838.390 ;
        RECT 1930.020 2838.380 1933.020 2838.390 ;
        RECT 2110.020 2838.380 2113.020 2838.390 ;
        RECT 2290.020 2838.380 2293.020 2838.390 ;
        RECT 2470.020 2838.380 2473.020 2838.390 ;
        RECT 2650.020 2838.380 2653.020 2838.390 ;
        RECT 2830.020 2838.380 2833.020 2838.390 ;
        RECT 2949.600 2838.380 2952.600 2838.390 ;
        RECT -32.980 2835.380 2952.600 2838.380 ;
        RECT -32.980 2835.370 -29.980 2835.380 ;
        RECT 130.020 2835.370 133.020 2835.380 ;
        RECT 310.020 2835.370 313.020 2835.380 ;
        RECT 490.020 2835.370 493.020 2835.380 ;
        RECT 670.020 2835.370 673.020 2835.380 ;
        RECT 850.020 2835.370 853.020 2835.380 ;
        RECT 1030.020 2835.370 1033.020 2835.380 ;
        RECT 1210.020 2835.370 1213.020 2835.380 ;
        RECT 1390.020 2835.370 1393.020 2835.380 ;
        RECT 1570.020 2835.370 1573.020 2835.380 ;
        RECT 1750.020 2835.370 1753.020 2835.380 ;
        RECT 1930.020 2835.370 1933.020 2835.380 ;
        RECT 2110.020 2835.370 2113.020 2835.380 ;
        RECT 2290.020 2835.370 2293.020 2835.380 ;
        RECT 2470.020 2835.370 2473.020 2835.380 ;
        RECT 2650.020 2835.370 2653.020 2835.380 ;
        RECT 2830.020 2835.370 2833.020 2835.380 ;
        RECT 2949.600 2835.370 2952.600 2835.380 ;
        RECT -32.980 2658.380 -29.980 2658.390 ;
        RECT 130.020 2658.380 133.020 2658.390 ;
        RECT 310.020 2658.380 313.020 2658.390 ;
        RECT 490.020 2658.380 493.020 2658.390 ;
        RECT 670.020 2658.380 673.020 2658.390 ;
        RECT 850.020 2658.380 853.020 2658.390 ;
        RECT 1030.020 2658.380 1033.020 2658.390 ;
        RECT 1210.020 2658.380 1213.020 2658.390 ;
        RECT 1390.020 2658.380 1393.020 2658.390 ;
        RECT 1570.020 2658.380 1573.020 2658.390 ;
        RECT 1750.020 2658.380 1753.020 2658.390 ;
        RECT 1930.020 2658.380 1933.020 2658.390 ;
        RECT 2110.020 2658.380 2113.020 2658.390 ;
        RECT 2290.020 2658.380 2293.020 2658.390 ;
        RECT 2470.020 2658.380 2473.020 2658.390 ;
        RECT 2650.020 2658.380 2653.020 2658.390 ;
        RECT 2830.020 2658.380 2833.020 2658.390 ;
        RECT 2949.600 2658.380 2952.600 2658.390 ;
        RECT -32.980 2655.380 2952.600 2658.380 ;
        RECT -32.980 2655.370 -29.980 2655.380 ;
        RECT 130.020 2655.370 133.020 2655.380 ;
        RECT 310.020 2655.370 313.020 2655.380 ;
        RECT 490.020 2655.370 493.020 2655.380 ;
        RECT 670.020 2655.370 673.020 2655.380 ;
        RECT 850.020 2655.370 853.020 2655.380 ;
        RECT 1030.020 2655.370 1033.020 2655.380 ;
        RECT 1210.020 2655.370 1213.020 2655.380 ;
        RECT 1390.020 2655.370 1393.020 2655.380 ;
        RECT 1570.020 2655.370 1573.020 2655.380 ;
        RECT 1750.020 2655.370 1753.020 2655.380 ;
        RECT 1930.020 2655.370 1933.020 2655.380 ;
        RECT 2110.020 2655.370 2113.020 2655.380 ;
        RECT 2290.020 2655.370 2293.020 2655.380 ;
        RECT 2470.020 2655.370 2473.020 2655.380 ;
        RECT 2650.020 2655.370 2653.020 2655.380 ;
        RECT 2830.020 2655.370 2833.020 2655.380 ;
        RECT 2949.600 2655.370 2952.600 2655.380 ;
        RECT -32.980 2478.380 -29.980 2478.390 ;
        RECT 130.020 2478.380 133.020 2478.390 ;
        RECT 310.020 2478.380 313.020 2478.390 ;
        RECT 490.020 2478.380 493.020 2478.390 ;
        RECT 670.020 2478.380 673.020 2478.390 ;
        RECT 850.020 2478.380 853.020 2478.390 ;
        RECT 1030.020 2478.380 1033.020 2478.390 ;
        RECT 1210.020 2478.380 1213.020 2478.390 ;
        RECT 1390.020 2478.380 1393.020 2478.390 ;
        RECT 1570.020 2478.380 1573.020 2478.390 ;
        RECT 1750.020 2478.380 1753.020 2478.390 ;
        RECT 1930.020 2478.380 1933.020 2478.390 ;
        RECT 2110.020 2478.380 2113.020 2478.390 ;
        RECT 2290.020 2478.380 2293.020 2478.390 ;
        RECT 2470.020 2478.380 2473.020 2478.390 ;
        RECT 2650.020 2478.380 2653.020 2478.390 ;
        RECT 2830.020 2478.380 2833.020 2478.390 ;
        RECT 2949.600 2478.380 2952.600 2478.390 ;
        RECT -32.980 2475.380 2952.600 2478.380 ;
        RECT -32.980 2475.370 -29.980 2475.380 ;
        RECT 130.020 2475.370 133.020 2475.380 ;
        RECT 310.020 2475.370 313.020 2475.380 ;
        RECT 490.020 2475.370 493.020 2475.380 ;
        RECT 670.020 2475.370 673.020 2475.380 ;
        RECT 850.020 2475.370 853.020 2475.380 ;
        RECT 1030.020 2475.370 1033.020 2475.380 ;
        RECT 1210.020 2475.370 1213.020 2475.380 ;
        RECT 1390.020 2475.370 1393.020 2475.380 ;
        RECT 1570.020 2475.370 1573.020 2475.380 ;
        RECT 1750.020 2475.370 1753.020 2475.380 ;
        RECT 1930.020 2475.370 1933.020 2475.380 ;
        RECT 2110.020 2475.370 2113.020 2475.380 ;
        RECT 2290.020 2475.370 2293.020 2475.380 ;
        RECT 2470.020 2475.370 2473.020 2475.380 ;
        RECT 2650.020 2475.370 2653.020 2475.380 ;
        RECT 2830.020 2475.370 2833.020 2475.380 ;
        RECT 2949.600 2475.370 2952.600 2475.380 ;
        RECT -32.980 2298.380 -29.980 2298.390 ;
        RECT 130.020 2298.380 133.020 2298.390 ;
        RECT 310.020 2298.380 313.020 2298.390 ;
        RECT 490.020 2298.380 493.020 2298.390 ;
        RECT 670.020 2298.380 673.020 2298.390 ;
        RECT 850.020 2298.380 853.020 2298.390 ;
        RECT 1030.020 2298.380 1033.020 2298.390 ;
        RECT 1210.020 2298.380 1213.020 2298.390 ;
        RECT 1390.020 2298.380 1393.020 2298.390 ;
        RECT 1570.020 2298.380 1573.020 2298.390 ;
        RECT 1750.020 2298.380 1753.020 2298.390 ;
        RECT 1930.020 2298.380 1933.020 2298.390 ;
        RECT 2110.020 2298.380 2113.020 2298.390 ;
        RECT 2290.020 2298.380 2293.020 2298.390 ;
        RECT 2470.020 2298.380 2473.020 2298.390 ;
        RECT 2650.020 2298.380 2653.020 2298.390 ;
        RECT 2830.020 2298.380 2833.020 2298.390 ;
        RECT 2949.600 2298.380 2952.600 2298.390 ;
        RECT -32.980 2295.380 2952.600 2298.380 ;
        RECT -32.980 2295.370 -29.980 2295.380 ;
        RECT 130.020 2295.370 133.020 2295.380 ;
        RECT 310.020 2295.370 313.020 2295.380 ;
        RECT 490.020 2295.370 493.020 2295.380 ;
        RECT 670.020 2295.370 673.020 2295.380 ;
        RECT 850.020 2295.370 853.020 2295.380 ;
        RECT 1030.020 2295.370 1033.020 2295.380 ;
        RECT 1210.020 2295.370 1213.020 2295.380 ;
        RECT 1390.020 2295.370 1393.020 2295.380 ;
        RECT 1570.020 2295.370 1573.020 2295.380 ;
        RECT 1750.020 2295.370 1753.020 2295.380 ;
        RECT 1930.020 2295.370 1933.020 2295.380 ;
        RECT 2110.020 2295.370 2113.020 2295.380 ;
        RECT 2290.020 2295.370 2293.020 2295.380 ;
        RECT 2470.020 2295.370 2473.020 2295.380 ;
        RECT 2650.020 2295.370 2653.020 2295.380 ;
        RECT 2830.020 2295.370 2833.020 2295.380 ;
        RECT 2949.600 2295.370 2952.600 2295.380 ;
        RECT -32.980 2118.380 -29.980 2118.390 ;
        RECT 130.020 2118.380 133.020 2118.390 ;
        RECT 310.020 2118.380 313.020 2118.390 ;
        RECT 490.020 2118.380 493.020 2118.390 ;
        RECT 670.020 2118.380 673.020 2118.390 ;
        RECT 850.020 2118.380 853.020 2118.390 ;
        RECT 1030.020 2118.380 1033.020 2118.390 ;
        RECT 1210.020 2118.380 1213.020 2118.390 ;
        RECT 1390.020 2118.380 1393.020 2118.390 ;
        RECT 1570.020 2118.380 1573.020 2118.390 ;
        RECT 1750.020 2118.380 1753.020 2118.390 ;
        RECT 1930.020 2118.380 1933.020 2118.390 ;
        RECT 2110.020 2118.380 2113.020 2118.390 ;
        RECT 2290.020 2118.380 2293.020 2118.390 ;
        RECT 2470.020 2118.380 2473.020 2118.390 ;
        RECT 2650.020 2118.380 2653.020 2118.390 ;
        RECT 2830.020 2118.380 2833.020 2118.390 ;
        RECT 2949.600 2118.380 2952.600 2118.390 ;
        RECT -32.980 2115.380 2952.600 2118.380 ;
        RECT -32.980 2115.370 -29.980 2115.380 ;
        RECT 130.020 2115.370 133.020 2115.380 ;
        RECT 310.020 2115.370 313.020 2115.380 ;
        RECT 490.020 2115.370 493.020 2115.380 ;
        RECT 670.020 2115.370 673.020 2115.380 ;
        RECT 850.020 2115.370 853.020 2115.380 ;
        RECT 1030.020 2115.370 1033.020 2115.380 ;
        RECT 1210.020 2115.370 1213.020 2115.380 ;
        RECT 1390.020 2115.370 1393.020 2115.380 ;
        RECT 1570.020 2115.370 1573.020 2115.380 ;
        RECT 1750.020 2115.370 1753.020 2115.380 ;
        RECT 1930.020 2115.370 1933.020 2115.380 ;
        RECT 2110.020 2115.370 2113.020 2115.380 ;
        RECT 2290.020 2115.370 2293.020 2115.380 ;
        RECT 2470.020 2115.370 2473.020 2115.380 ;
        RECT 2650.020 2115.370 2653.020 2115.380 ;
        RECT 2830.020 2115.370 2833.020 2115.380 ;
        RECT 2949.600 2115.370 2952.600 2115.380 ;
        RECT -32.980 1938.380 -29.980 1938.390 ;
        RECT 130.020 1938.380 133.020 1938.390 ;
        RECT 310.020 1938.380 313.020 1938.390 ;
        RECT 490.020 1938.380 493.020 1938.390 ;
        RECT 670.020 1938.380 673.020 1938.390 ;
        RECT 850.020 1938.380 853.020 1938.390 ;
        RECT 1030.020 1938.380 1033.020 1938.390 ;
        RECT 1210.020 1938.380 1213.020 1938.390 ;
        RECT 1390.020 1938.380 1393.020 1938.390 ;
        RECT 1570.020 1938.380 1573.020 1938.390 ;
        RECT 1750.020 1938.380 1753.020 1938.390 ;
        RECT 1930.020 1938.380 1933.020 1938.390 ;
        RECT 2110.020 1938.380 2113.020 1938.390 ;
        RECT 2290.020 1938.380 2293.020 1938.390 ;
        RECT 2470.020 1938.380 2473.020 1938.390 ;
        RECT 2650.020 1938.380 2653.020 1938.390 ;
        RECT 2830.020 1938.380 2833.020 1938.390 ;
        RECT 2949.600 1938.380 2952.600 1938.390 ;
        RECT -32.980 1935.380 2952.600 1938.380 ;
        RECT -32.980 1935.370 -29.980 1935.380 ;
        RECT 130.020 1935.370 133.020 1935.380 ;
        RECT 310.020 1935.370 313.020 1935.380 ;
        RECT 490.020 1935.370 493.020 1935.380 ;
        RECT 670.020 1935.370 673.020 1935.380 ;
        RECT 850.020 1935.370 853.020 1935.380 ;
        RECT 1030.020 1935.370 1033.020 1935.380 ;
        RECT 1210.020 1935.370 1213.020 1935.380 ;
        RECT 1390.020 1935.370 1393.020 1935.380 ;
        RECT 1570.020 1935.370 1573.020 1935.380 ;
        RECT 1750.020 1935.370 1753.020 1935.380 ;
        RECT 1930.020 1935.370 1933.020 1935.380 ;
        RECT 2110.020 1935.370 2113.020 1935.380 ;
        RECT 2290.020 1935.370 2293.020 1935.380 ;
        RECT 2470.020 1935.370 2473.020 1935.380 ;
        RECT 2650.020 1935.370 2653.020 1935.380 ;
        RECT 2830.020 1935.370 2833.020 1935.380 ;
        RECT 2949.600 1935.370 2952.600 1935.380 ;
        RECT -32.980 1758.380 -29.980 1758.390 ;
        RECT 130.020 1758.380 133.020 1758.390 ;
        RECT 310.020 1758.380 313.020 1758.390 ;
        RECT 490.020 1758.380 493.020 1758.390 ;
        RECT 670.020 1758.380 673.020 1758.390 ;
        RECT 850.020 1758.380 853.020 1758.390 ;
        RECT 1030.020 1758.380 1033.020 1758.390 ;
        RECT 1210.020 1758.380 1213.020 1758.390 ;
        RECT 1390.020 1758.380 1393.020 1758.390 ;
        RECT 1570.020 1758.380 1573.020 1758.390 ;
        RECT 1750.020 1758.380 1753.020 1758.390 ;
        RECT 1930.020 1758.380 1933.020 1758.390 ;
        RECT 2110.020 1758.380 2113.020 1758.390 ;
        RECT 2290.020 1758.380 2293.020 1758.390 ;
        RECT 2470.020 1758.380 2473.020 1758.390 ;
        RECT 2650.020 1758.380 2653.020 1758.390 ;
        RECT 2830.020 1758.380 2833.020 1758.390 ;
        RECT 2949.600 1758.380 2952.600 1758.390 ;
        RECT -32.980 1755.380 2952.600 1758.380 ;
        RECT -32.980 1755.370 -29.980 1755.380 ;
        RECT 130.020 1755.370 133.020 1755.380 ;
        RECT 310.020 1755.370 313.020 1755.380 ;
        RECT 490.020 1755.370 493.020 1755.380 ;
        RECT 670.020 1755.370 673.020 1755.380 ;
        RECT 850.020 1755.370 853.020 1755.380 ;
        RECT 1030.020 1755.370 1033.020 1755.380 ;
        RECT 1210.020 1755.370 1213.020 1755.380 ;
        RECT 1390.020 1755.370 1393.020 1755.380 ;
        RECT 1570.020 1755.370 1573.020 1755.380 ;
        RECT 1750.020 1755.370 1753.020 1755.380 ;
        RECT 1930.020 1755.370 1933.020 1755.380 ;
        RECT 2110.020 1755.370 2113.020 1755.380 ;
        RECT 2290.020 1755.370 2293.020 1755.380 ;
        RECT 2470.020 1755.370 2473.020 1755.380 ;
        RECT 2650.020 1755.370 2653.020 1755.380 ;
        RECT 2830.020 1755.370 2833.020 1755.380 ;
        RECT 2949.600 1755.370 2952.600 1755.380 ;
        RECT -32.980 1578.380 -29.980 1578.390 ;
        RECT 130.020 1578.380 133.020 1578.390 ;
        RECT 310.020 1578.380 313.020 1578.390 ;
        RECT 490.020 1578.380 493.020 1578.390 ;
        RECT 670.020 1578.380 673.020 1578.390 ;
        RECT 850.020 1578.380 853.020 1578.390 ;
        RECT 1030.020 1578.380 1033.020 1578.390 ;
        RECT 1210.020 1578.380 1213.020 1578.390 ;
        RECT 1390.020 1578.380 1393.020 1578.390 ;
        RECT 1570.020 1578.380 1573.020 1578.390 ;
        RECT 1750.020 1578.380 1753.020 1578.390 ;
        RECT 1930.020 1578.380 1933.020 1578.390 ;
        RECT 2110.020 1578.380 2113.020 1578.390 ;
        RECT 2290.020 1578.380 2293.020 1578.390 ;
        RECT 2470.020 1578.380 2473.020 1578.390 ;
        RECT 2650.020 1578.380 2653.020 1578.390 ;
        RECT 2830.020 1578.380 2833.020 1578.390 ;
        RECT 2949.600 1578.380 2952.600 1578.390 ;
        RECT -32.980 1575.380 2952.600 1578.380 ;
        RECT -32.980 1575.370 -29.980 1575.380 ;
        RECT 130.020 1575.370 133.020 1575.380 ;
        RECT 310.020 1575.370 313.020 1575.380 ;
        RECT 490.020 1575.370 493.020 1575.380 ;
        RECT 670.020 1575.370 673.020 1575.380 ;
        RECT 850.020 1575.370 853.020 1575.380 ;
        RECT 1030.020 1575.370 1033.020 1575.380 ;
        RECT 1210.020 1575.370 1213.020 1575.380 ;
        RECT 1390.020 1575.370 1393.020 1575.380 ;
        RECT 1570.020 1575.370 1573.020 1575.380 ;
        RECT 1750.020 1575.370 1753.020 1575.380 ;
        RECT 1930.020 1575.370 1933.020 1575.380 ;
        RECT 2110.020 1575.370 2113.020 1575.380 ;
        RECT 2290.020 1575.370 2293.020 1575.380 ;
        RECT 2470.020 1575.370 2473.020 1575.380 ;
        RECT 2650.020 1575.370 2653.020 1575.380 ;
        RECT 2830.020 1575.370 2833.020 1575.380 ;
        RECT 2949.600 1575.370 2952.600 1575.380 ;
        RECT -32.980 1398.380 -29.980 1398.390 ;
        RECT 130.020 1398.380 133.020 1398.390 ;
        RECT 310.020 1398.380 313.020 1398.390 ;
        RECT 490.020 1398.380 493.020 1398.390 ;
        RECT 670.020 1398.380 673.020 1398.390 ;
        RECT 850.020 1398.380 853.020 1398.390 ;
        RECT 1030.020 1398.380 1033.020 1398.390 ;
        RECT 1210.020 1398.380 1213.020 1398.390 ;
        RECT 1390.020 1398.380 1393.020 1398.390 ;
        RECT 1570.020 1398.380 1573.020 1398.390 ;
        RECT 1750.020 1398.380 1753.020 1398.390 ;
        RECT 1930.020 1398.380 1933.020 1398.390 ;
        RECT 2110.020 1398.380 2113.020 1398.390 ;
        RECT 2290.020 1398.380 2293.020 1398.390 ;
        RECT 2470.020 1398.380 2473.020 1398.390 ;
        RECT 2650.020 1398.380 2653.020 1398.390 ;
        RECT 2830.020 1398.380 2833.020 1398.390 ;
        RECT 2949.600 1398.380 2952.600 1398.390 ;
        RECT -32.980 1395.380 2952.600 1398.380 ;
        RECT -32.980 1395.370 -29.980 1395.380 ;
        RECT 130.020 1395.370 133.020 1395.380 ;
        RECT 310.020 1395.370 313.020 1395.380 ;
        RECT 490.020 1395.370 493.020 1395.380 ;
        RECT 670.020 1395.370 673.020 1395.380 ;
        RECT 850.020 1395.370 853.020 1395.380 ;
        RECT 1030.020 1395.370 1033.020 1395.380 ;
        RECT 1210.020 1395.370 1213.020 1395.380 ;
        RECT 1390.020 1395.370 1393.020 1395.380 ;
        RECT 1570.020 1395.370 1573.020 1395.380 ;
        RECT 1750.020 1395.370 1753.020 1395.380 ;
        RECT 1930.020 1395.370 1933.020 1395.380 ;
        RECT 2110.020 1395.370 2113.020 1395.380 ;
        RECT 2290.020 1395.370 2293.020 1395.380 ;
        RECT 2470.020 1395.370 2473.020 1395.380 ;
        RECT 2650.020 1395.370 2653.020 1395.380 ;
        RECT 2830.020 1395.370 2833.020 1395.380 ;
        RECT 2949.600 1395.370 2952.600 1395.380 ;
        RECT -32.980 1218.380 -29.980 1218.390 ;
        RECT 130.020 1218.380 133.020 1218.390 ;
        RECT 310.020 1218.380 313.020 1218.390 ;
        RECT 490.020 1218.380 493.020 1218.390 ;
        RECT 670.020 1218.380 673.020 1218.390 ;
        RECT 850.020 1218.380 853.020 1218.390 ;
        RECT 1030.020 1218.380 1033.020 1218.390 ;
        RECT 1210.020 1218.380 1213.020 1218.390 ;
        RECT 1390.020 1218.380 1393.020 1218.390 ;
        RECT 1570.020 1218.380 1573.020 1218.390 ;
        RECT 1750.020 1218.380 1753.020 1218.390 ;
        RECT 1930.020 1218.380 1933.020 1218.390 ;
        RECT 2110.020 1218.380 2113.020 1218.390 ;
        RECT 2290.020 1218.380 2293.020 1218.390 ;
        RECT 2470.020 1218.380 2473.020 1218.390 ;
        RECT 2650.020 1218.380 2653.020 1218.390 ;
        RECT 2830.020 1218.380 2833.020 1218.390 ;
        RECT 2949.600 1218.380 2952.600 1218.390 ;
        RECT -32.980 1215.380 2952.600 1218.380 ;
        RECT -32.980 1215.370 -29.980 1215.380 ;
        RECT 130.020 1215.370 133.020 1215.380 ;
        RECT 310.020 1215.370 313.020 1215.380 ;
        RECT 490.020 1215.370 493.020 1215.380 ;
        RECT 670.020 1215.370 673.020 1215.380 ;
        RECT 850.020 1215.370 853.020 1215.380 ;
        RECT 1030.020 1215.370 1033.020 1215.380 ;
        RECT 1210.020 1215.370 1213.020 1215.380 ;
        RECT 1390.020 1215.370 1393.020 1215.380 ;
        RECT 1570.020 1215.370 1573.020 1215.380 ;
        RECT 1750.020 1215.370 1753.020 1215.380 ;
        RECT 1930.020 1215.370 1933.020 1215.380 ;
        RECT 2110.020 1215.370 2113.020 1215.380 ;
        RECT 2290.020 1215.370 2293.020 1215.380 ;
        RECT 2470.020 1215.370 2473.020 1215.380 ;
        RECT 2650.020 1215.370 2653.020 1215.380 ;
        RECT 2830.020 1215.370 2833.020 1215.380 ;
        RECT 2949.600 1215.370 2952.600 1215.380 ;
        RECT -32.980 1038.380 -29.980 1038.390 ;
        RECT 130.020 1038.380 133.020 1038.390 ;
        RECT 310.020 1038.380 313.020 1038.390 ;
        RECT 490.020 1038.380 493.020 1038.390 ;
        RECT 670.020 1038.380 673.020 1038.390 ;
        RECT 850.020 1038.380 853.020 1038.390 ;
        RECT 1030.020 1038.380 1033.020 1038.390 ;
        RECT 1210.020 1038.380 1213.020 1038.390 ;
        RECT 1390.020 1038.380 1393.020 1038.390 ;
        RECT 1570.020 1038.380 1573.020 1038.390 ;
        RECT 1750.020 1038.380 1753.020 1038.390 ;
        RECT 1930.020 1038.380 1933.020 1038.390 ;
        RECT 2110.020 1038.380 2113.020 1038.390 ;
        RECT 2290.020 1038.380 2293.020 1038.390 ;
        RECT 2470.020 1038.380 2473.020 1038.390 ;
        RECT 2650.020 1038.380 2653.020 1038.390 ;
        RECT 2830.020 1038.380 2833.020 1038.390 ;
        RECT 2949.600 1038.380 2952.600 1038.390 ;
        RECT -32.980 1035.380 2952.600 1038.380 ;
        RECT -32.980 1035.370 -29.980 1035.380 ;
        RECT 130.020 1035.370 133.020 1035.380 ;
        RECT 310.020 1035.370 313.020 1035.380 ;
        RECT 490.020 1035.370 493.020 1035.380 ;
        RECT 670.020 1035.370 673.020 1035.380 ;
        RECT 850.020 1035.370 853.020 1035.380 ;
        RECT 1030.020 1035.370 1033.020 1035.380 ;
        RECT 1210.020 1035.370 1213.020 1035.380 ;
        RECT 1390.020 1035.370 1393.020 1035.380 ;
        RECT 1570.020 1035.370 1573.020 1035.380 ;
        RECT 1750.020 1035.370 1753.020 1035.380 ;
        RECT 1930.020 1035.370 1933.020 1035.380 ;
        RECT 2110.020 1035.370 2113.020 1035.380 ;
        RECT 2290.020 1035.370 2293.020 1035.380 ;
        RECT 2470.020 1035.370 2473.020 1035.380 ;
        RECT 2650.020 1035.370 2653.020 1035.380 ;
        RECT 2830.020 1035.370 2833.020 1035.380 ;
        RECT 2949.600 1035.370 2952.600 1035.380 ;
        RECT -32.980 858.380 -29.980 858.390 ;
        RECT 130.020 858.380 133.020 858.390 ;
        RECT 310.020 858.380 313.020 858.390 ;
        RECT 490.020 858.380 493.020 858.390 ;
        RECT 670.020 858.380 673.020 858.390 ;
        RECT 850.020 858.380 853.020 858.390 ;
        RECT 1030.020 858.380 1033.020 858.390 ;
        RECT 1210.020 858.380 1213.020 858.390 ;
        RECT 1390.020 858.380 1393.020 858.390 ;
        RECT 1570.020 858.380 1573.020 858.390 ;
        RECT 1750.020 858.380 1753.020 858.390 ;
        RECT 1930.020 858.380 1933.020 858.390 ;
        RECT 2110.020 858.380 2113.020 858.390 ;
        RECT 2290.020 858.380 2293.020 858.390 ;
        RECT 2470.020 858.380 2473.020 858.390 ;
        RECT 2650.020 858.380 2653.020 858.390 ;
        RECT 2830.020 858.380 2833.020 858.390 ;
        RECT 2949.600 858.380 2952.600 858.390 ;
        RECT -32.980 855.380 2952.600 858.380 ;
        RECT -32.980 855.370 -29.980 855.380 ;
        RECT 130.020 855.370 133.020 855.380 ;
        RECT 310.020 855.370 313.020 855.380 ;
        RECT 490.020 855.370 493.020 855.380 ;
        RECT 670.020 855.370 673.020 855.380 ;
        RECT 850.020 855.370 853.020 855.380 ;
        RECT 1030.020 855.370 1033.020 855.380 ;
        RECT 1210.020 855.370 1213.020 855.380 ;
        RECT 1390.020 855.370 1393.020 855.380 ;
        RECT 1570.020 855.370 1573.020 855.380 ;
        RECT 1750.020 855.370 1753.020 855.380 ;
        RECT 1930.020 855.370 1933.020 855.380 ;
        RECT 2110.020 855.370 2113.020 855.380 ;
        RECT 2290.020 855.370 2293.020 855.380 ;
        RECT 2470.020 855.370 2473.020 855.380 ;
        RECT 2650.020 855.370 2653.020 855.380 ;
        RECT 2830.020 855.370 2833.020 855.380 ;
        RECT 2949.600 855.370 2952.600 855.380 ;
        RECT -32.980 678.380 -29.980 678.390 ;
        RECT 130.020 678.380 133.020 678.390 ;
        RECT 310.020 678.380 313.020 678.390 ;
        RECT 490.020 678.380 493.020 678.390 ;
        RECT 670.020 678.380 673.020 678.390 ;
        RECT 850.020 678.380 853.020 678.390 ;
        RECT 1030.020 678.380 1033.020 678.390 ;
        RECT 1210.020 678.380 1213.020 678.390 ;
        RECT 1390.020 678.380 1393.020 678.390 ;
        RECT 1570.020 678.380 1573.020 678.390 ;
        RECT 1750.020 678.380 1753.020 678.390 ;
        RECT 1930.020 678.380 1933.020 678.390 ;
        RECT 2110.020 678.380 2113.020 678.390 ;
        RECT 2290.020 678.380 2293.020 678.390 ;
        RECT 2470.020 678.380 2473.020 678.390 ;
        RECT 2650.020 678.380 2653.020 678.390 ;
        RECT 2830.020 678.380 2833.020 678.390 ;
        RECT 2949.600 678.380 2952.600 678.390 ;
        RECT -32.980 675.380 2952.600 678.380 ;
        RECT -32.980 675.370 -29.980 675.380 ;
        RECT 130.020 675.370 133.020 675.380 ;
        RECT 310.020 675.370 313.020 675.380 ;
        RECT 490.020 675.370 493.020 675.380 ;
        RECT 670.020 675.370 673.020 675.380 ;
        RECT 850.020 675.370 853.020 675.380 ;
        RECT 1030.020 675.370 1033.020 675.380 ;
        RECT 1210.020 675.370 1213.020 675.380 ;
        RECT 1390.020 675.370 1393.020 675.380 ;
        RECT 1570.020 675.370 1573.020 675.380 ;
        RECT 1750.020 675.370 1753.020 675.380 ;
        RECT 1930.020 675.370 1933.020 675.380 ;
        RECT 2110.020 675.370 2113.020 675.380 ;
        RECT 2290.020 675.370 2293.020 675.380 ;
        RECT 2470.020 675.370 2473.020 675.380 ;
        RECT 2650.020 675.370 2653.020 675.380 ;
        RECT 2830.020 675.370 2833.020 675.380 ;
        RECT 2949.600 675.370 2952.600 675.380 ;
        RECT -32.980 498.380 -29.980 498.390 ;
        RECT 130.020 498.380 133.020 498.390 ;
        RECT 310.020 498.380 313.020 498.390 ;
        RECT 490.020 498.380 493.020 498.390 ;
        RECT 670.020 498.380 673.020 498.390 ;
        RECT 850.020 498.380 853.020 498.390 ;
        RECT 1030.020 498.380 1033.020 498.390 ;
        RECT 1210.020 498.380 1213.020 498.390 ;
        RECT 1390.020 498.380 1393.020 498.390 ;
        RECT 1570.020 498.380 1573.020 498.390 ;
        RECT 1750.020 498.380 1753.020 498.390 ;
        RECT 1930.020 498.380 1933.020 498.390 ;
        RECT 2110.020 498.380 2113.020 498.390 ;
        RECT 2290.020 498.380 2293.020 498.390 ;
        RECT 2470.020 498.380 2473.020 498.390 ;
        RECT 2650.020 498.380 2653.020 498.390 ;
        RECT 2830.020 498.380 2833.020 498.390 ;
        RECT 2949.600 498.380 2952.600 498.390 ;
        RECT -32.980 495.380 2952.600 498.380 ;
        RECT -32.980 495.370 -29.980 495.380 ;
        RECT 130.020 495.370 133.020 495.380 ;
        RECT 310.020 495.370 313.020 495.380 ;
        RECT 490.020 495.370 493.020 495.380 ;
        RECT 670.020 495.370 673.020 495.380 ;
        RECT 850.020 495.370 853.020 495.380 ;
        RECT 1030.020 495.370 1033.020 495.380 ;
        RECT 1210.020 495.370 1213.020 495.380 ;
        RECT 1390.020 495.370 1393.020 495.380 ;
        RECT 1570.020 495.370 1573.020 495.380 ;
        RECT 1750.020 495.370 1753.020 495.380 ;
        RECT 1930.020 495.370 1933.020 495.380 ;
        RECT 2110.020 495.370 2113.020 495.380 ;
        RECT 2290.020 495.370 2293.020 495.380 ;
        RECT 2470.020 495.370 2473.020 495.380 ;
        RECT 2650.020 495.370 2653.020 495.380 ;
        RECT 2830.020 495.370 2833.020 495.380 ;
        RECT 2949.600 495.370 2952.600 495.380 ;
        RECT -32.980 318.380 -29.980 318.390 ;
        RECT 130.020 318.380 133.020 318.390 ;
        RECT 310.020 318.380 313.020 318.390 ;
        RECT 490.020 318.380 493.020 318.390 ;
        RECT 670.020 318.380 673.020 318.390 ;
        RECT 850.020 318.380 853.020 318.390 ;
        RECT 1030.020 318.380 1033.020 318.390 ;
        RECT 1210.020 318.380 1213.020 318.390 ;
        RECT 1390.020 318.380 1393.020 318.390 ;
        RECT 1570.020 318.380 1573.020 318.390 ;
        RECT 1750.020 318.380 1753.020 318.390 ;
        RECT 1930.020 318.380 1933.020 318.390 ;
        RECT 2110.020 318.380 2113.020 318.390 ;
        RECT 2290.020 318.380 2293.020 318.390 ;
        RECT 2470.020 318.380 2473.020 318.390 ;
        RECT 2650.020 318.380 2653.020 318.390 ;
        RECT 2830.020 318.380 2833.020 318.390 ;
        RECT 2949.600 318.380 2952.600 318.390 ;
        RECT -32.980 315.380 2952.600 318.380 ;
        RECT -32.980 315.370 -29.980 315.380 ;
        RECT 130.020 315.370 133.020 315.380 ;
        RECT 310.020 315.370 313.020 315.380 ;
        RECT 490.020 315.370 493.020 315.380 ;
        RECT 670.020 315.370 673.020 315.380 ;
        RECT 850.020 315.370 853.020 315.380 ;
        RECT 1030.020 315.370 1033.020 315.380 ;
        RECT 1210.020 315.370 1213.020 315.380 ;
        RECT 1390.020 315.370 1393.020 315.380 ;
        RECT 1570.020 315.370 1573.020 315.380 ;
        RECT 1750.020 315.370 1753.020 315.380 ;
        RECT 1930.020 315.370 1933.020 315.380 ;
        RECT 2110.020 315.370 2113.020 315.380 ;
        RECT 2290.020 315.370 2293.020 315.380 ;
        RECT 2470.020 315.370 2473.020 315.380 ;
        RECT 2650.020 315.370 2653.020 315.380 ;
        RECT 2830.020 315.370 2833.020 315.380 ;
        RECT 2949.600 315.370 2952.600 315.380 ;
        RECT -32.980 138.380 -29.980 138.390 ;
        RECT 130.020 138.380 133.020 138.390 ;
        RECT 310.020 138.380 313.020 138.390 ;
        RECT 490.020 138.380 493.020 138.390 ;
        RECT 670.020 138.380 673.020 138.390 ;
        RECT 850.020 138.380 853.020 138.390 ;
        RECT 1030.020 138.380 1033.020 138.390 ;
        RECT 1210.020 138.380 1213.020 138.390 ;
        RECT 1390.020 138.380 1393.020 138.390 ;
        RECT 1570.020 138.380 1573.020 138.390 ;
        RECT 1750.020 138.380 1753.020 138.390 ;
        RECT 1930.020 138.380 1933.020 138.390 ;
        RECT 2110.020 138.380 2113.020 138.390 ;
        RECT 2290.020 138.380 2293.020 138.390 ;
        RECT 2470.020 138.380 2473.020 138.390 ;
        RECT 2650.020 138.380 2653.020 138.390 ;
        RECT 2830.020 138.380 2833.020 138.390 ;
        RECT 2949.600 138.380 2952.600 138.390 ;
        RECT -32.980 135.380 2952.600 138.380 ;
        RECT -32.980 135.370 -29.980 135.380 ;
        RECT 130.020 135.370 133.020 135.380 ;
        RECT 310.020 135.370 313.020 135.380 ;
        RECT 490.020 135.370 493.020 135.380 ;
        RECT 670.020 135.370 673.020 135.380 ;
        RECT 850.020 135.370 853.020 135.380 ;
        RECT 1030.020 135.370 1033.020 135.380 ;
        RECT 1210.020 135.370 1213.020 135.380 ;
        RECT 1390.020 135.370 1393.020 135.380 ;
        RECT 1570.020 135.370 1573.020 135.380 ;
        RECT 1750.020 135.370 1753.020 135.380 ;
        RECT 1930.020 135.370 1933.020 135.380 ;
        RECT 2110.020 135.370 2113.020 135.380 ;
        RECT 2290.020 135.370 2293.020 135.380 ;
        RECT 2470.020 135.370 2473.020 135.380 ;
        RECT 2650.020 135.370 2653.020 135.380 ;
        RECT 2830.020 135.370 2833.020 135.380 ;
        RECT 2949.600 135.370 2952.600 135.380 ;
        RECT -32.980 -24.620 -29.980 -24.610 ;
        RECT 130.020 -24.620 133.020 -24.610 ;
        RECT 310.020 -24.620 313.020 -24.610 ;
        RECT 490.020 -24.620 493.020 -24.610 ;
        RECT 670.020 -24.620 673.020 -24.610 ;
        RECT 850.020 -24.620 853.020 -24.610 ;
        RECT 1030.020 -24.620 1033.020 -24.610 ;
        RECT 1210.020 -24.620 1213.020 -24.610 ;
        RECT 1390.020 -24.620 1393.020 -24.610 ;
        RECT 1570.020 -24.620 1573.020 -24.610 ;
        RECT 1750.020 -24.620 1753.020 -24.610 ;
        RECT 1930.020 -24.620 1933.020 -24.610 ;
        RECT 2110.020 -24.620 2113.020 -24.610 ;
        RECT 2290.020 -24.620 2293.020 -24.610 ;
        RECT 2470.020 -24.620 2473.020 -24.610 ;
        RECT 2650.020 -24.620 2653.020 -24.610 ;
        RECT 2830.020 -24.620 2833.020 -24.610 ;
        RECT 2949.600 -24.620 2952.600 -24.610 ;
        RECT -32.980 -27.620 2952.600 -24.620 ;
        RECT -32.980 -27.630 -29.980 -27.620 ;
        RECT 130.020 -27.630 133.020 -27.620 ;
        RECT 310.020 -27.630 313.020 -27.620 ;
        RECT 490.020 -27.630 493.020 -27.620 ;
        RECT 670.020 -27.630 673.020 -27.620 ;
        RECT 850.020 -27.630 853.020 -27.620 ;
        RECT 1030.020 -27.630 1033.020 -27.620 ;
        RECT 1210.020 -27.630 1213.020 -27.620 ;
        RECT 1390.020 -27.630 1393.020 -27.620 ;
        RECT 1570.020 -27.630 1573.020 -27.620 ;
        RECT 1750.020 -27.630 1753.020 -27.620 ;
        RECT 1930.020 -27.630 1933.020 -27.620 ;
        RECT 2110.020 -27.630 2113.020 -27.620 ;
        RECT 2290.020 -27.630 2293.020 -27.620 ;
        RECT 2470.020 -27.630 2473.020 -27.620 ;
        RECT 2650.020 -27.630 2653.020 -27.620 ;
        RECT 2830.020 -27.630 2833.020 -27.620 ;
        RECT 2949.600 -27.630 2952.600 -27.620 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -37.580 -32.220 -34.580 3551.900 ;
        RECT 58.020 -36.820 61.020 3556.500 ;
        RECT 238.020 -36.820 241.020 3556.500 ;
        RECT 418.020 -36.820 421.020 3556.500 ;
        RECT 598.020 -36.820 601.020 3556.500 ;
        RECT 778.020 -36.820 781.020 3556.500 ;
        RECT 958.020 -36.820 961.020 3556.500 ;
        RECT 1138.020 -36.820 1141.020 3556.500 ;
        RECT 1318.020 -36.820 1321.020 3556.500 ;
        RECT 1498.020 -36.820 1501.020 3556.500 ;
        RECT 1678.020 -36.820 1681.020 3556.500 ;
        RECT 1858.020 -36.820 1861.020 3556.500 ;
        RECT 2038.020 -36.820 2041.020 3556.500 ;
        RECT 2218.020 -36.820 2221.020 3556.500 ;
        RECT 2398.020 -36.820 2401.020 3556.500 ;
        RECT 2578.020 -36.820 2581.020 3556.500 ;
        RECT 2758.020 -36.820 2761.020 3556.500 ;
        RECT 2954.200 -32.220 2957.200 3551.900 ;
      LAYER via4 ;
        RECT -36.670 3550.610 -35.490 3551.790 ;
        RECT -36.670 3549.010 -35.490 3550.190 ;
        RECT -36.670 3485.090 -35.490 3486.270 ;
        RECT -36.670 3483.490 -35.490 3484.670 ;
        RECT -36.670 3305.090 -35.490 3306.270 ;
        RECT -36.670 3303.490 -35.490 3304.670 ;
        RECT -36.670 3125.090 -35.490 3126.270 ;
        RECT -36.670 3123.490 -35.490 3124.670 ;
        RECT -36.670 2945.090 -35.490 2946.270 ;
        RECT -36.670 2943.490 -35.490 2944.670 ;
        RECT -36.670 2765.090 -35.490 2766.270 ;
        RECT -36.670 2763.490 -35.490 2764.670 ;
        RECT -36.670 2585.090 -35.490 2586.270 ;
        RECT -36.670 2583.490 -35.490 2584.670 ;
        RECT -36.670 2405.090 -35.490 2406.270 ;
        RECT -36.670 2403.490 -35.490 2404.670 ;
        RECT -36.670 2225.090 -35.490 2226.270 ;
        RECT -36.670 2223.490 -35.490 2224.670 ;
        RECT -36.670 2045.090 -35.490 2046.270 ;
        RECT -36.670 2043.490 -35.490 2044.670 ;
        RECT -36.670 1865.090 -35.490 1866.270 ;
        RECT -36.670 1863.490 -35.490 1864.670 ;
        RECT -36.670 1685.090 -35.490 1686.270 ;
        RECT -36.670 1683.490 -35.490 1684.670 ;
        RECT -36.670 1505.090 -35.490 1506.270 ;
        RECT -36.670 1503.490 -35.490 1504.670 ;
        RECT -36.670 1325.090 -35.490 1326.270 ;
        RECT -36.670 1323.490 -35.490 1324.670 ;
        RECT -36.670 1145.090 -35.490 1146.270 ;
        RECT -36.670 1143.490 -35.490 1144.670 ;
        RECT -36.670 965.090 -35.490 966.270 ;
        RECT -36.670 963.490 -35.490 964.670 ;
        RECT -36.670 785.090 -35.490 786.270 ;
        RECT -36.670 783.490 -35.490 784.670 ;
        RECT -36.670 605.090 -35.490 606.270 ;
        RECT -36.670 603.490 -35.490 604.670 ;
        RECT -36.670 425.090 -35.490 426.270 ;
        RECT -36.670 423.490 -35.490 424.670 ;
        RECT -36.670 245.090 -35.490 246.270 ;
        RECT -36.670 243.490 -35.490 244.670 ;
        RECT -36.670 65.090 -35.490 66.270 ;
        RECT -36.670 63.490 -35.490 64.670 ;
        RECT -36.670 -30.510 -35.490 -29.330 ;
        RECT -36.670 -32.110 -35.490 -30.930 ;
        RECT 58.930 3550.610 60.110 3551.790 ;
        RECT 58.930 3549.010 60.110 3550.190 ;
        RECT 58.930 3485.090 60.110 3486.270 ;
        RECT 58.930 3483.490 60.110 3484.670 ;
        RECT 58.930 3305.090 60.110 3306.270 ;
        RECT 58.930 3303.490 60.110 3304.670 ;
        RECT 58.930 3125.090 60.110 3126.270 ;
        RECT 58.930 3123.490 60.110 3124.670 ;
        RECT 58.930 2945.090 60.110 2946.270 ;
        RECT 58.930 2943.490 60.110 2944.670 ;
        RECT 58.930 2765.090 60.110 2766.270 ;
        RECT 58.930 2763.490 60.110 2764.670 ;
        RECT 58.930 2585.090 60.110 2586.270 ;
        RECT 58.930 2583.490 60.110 2584.670 ;
        RECT 58.930 2405.090 60.110 2406.270 ;
        RECT 58.930 2403.490 60.110 2404.670 ;
        RECT 58.930 2225.090 60.110 2226.270 ;
        RECT 58.930 2223.490 60.110 2224.670 ;
        RECT 58.930 2045.090 60.110 2046.270 ;
        RECT 58.930 2043.490 60.110 2044.670 ;
        RECT 58.930 1865.090 60.110 1866.270 ;
        RECT 58.930 1863.490 60.110 1864.670 ;
        RECT 58.930 1685.090 60.110 1686.270 ;
        RECT 58.930 1683.490 60.110 1684.670 ;
        RECT 58.930 1505.090 60.110 1506.270 ;
        RECT 58.930 1503.490 60.110 1504.670 ;
        RECT 58.930 1325.090 60.110 1326.270 ;
        RECT 58.930 1323.490 60.110 1324.670 ;
        RECT 58.930 1145.090 60.110 1146.270 ;
        RECT 58.930 1143.490 60.110 1144.670 ;
        RECT 58.930 965.090 60.110 966.270 ;
        RECT 58.930 963.490 60.110 964.670 ;
        RECT 58.930 785.090 60.110 786.270 ;
        RECT 58.930 783.490 60.110 784.670 ;
        RECT 58.930 605.090 60.110 606.270 ;
        RECT 58.930 603.490 60.110 604.670 ;
        RECT 58.930 425.090 60.110 426.270 ;
        RECT 58.930 423.490 60.110 424.670 ;
        RECT 58.930 245.090 60.110 246.270 ;
        RECT 58.930 243.490 60.110 244.670 ;
        RECT 58.930 65.090 60.110 66.270 ;
        RECT 58.930 63.490 60.110 64.670 ;
        RECT 58.930 -30.510 60.110 -29.330 ;
        RECT 58.930 -32.110 60.110 -30.930 ;
        RECT 238.930 3550.610 240.110 3551.790 ;
        RECT 238.930 3549.010 240.110 3550.190 ;
        RECT 238.930 3485.090 240.110 3486.270 ;
        RECT 238.930 3483.490 240.110 3484.670 ;
        RECT 238.930 3305.090 240.110 3306.270 ;
        RECT 238.930 3303.490 240.110 3304.670 ;
        RECT 238.930 3125.090 240.110 3126.270 ;
        RECT 238.930 3123.490 240.110 3124.670 ;
        RECT 238.930 2945.090 240.110 2946.270 ;
        RECT 238.930 2943.490 240.110 2944.670 ;
        RECT 238.930 2765.090 240.110 2766.270 ;
        RECT 238.930 2763.490 240.110 2764.670 ;
        RECT 238.930 2585.090 240.110 2586.270 ;
        RECT 238.930 2583.490 240.110 2584.670 ;
        RECT 238.930 2405.090 240.110 2406.270 ;
        RECT 238.930 2403.490 240.110 2404.670 ;
        RECT 238.930 2225.090 240.110 2226.270 ;
        RECT 238.930 2223.490 240.110 2224.670 ;
        RECT 238.930 2045.090 240.110 2046.270 ;
        RECT 238.930 2043.490 240.110 2044.670 ;
        RECT 238.930 1865.090 240.110 1866.270 ;
        RECT 238.930 1863.490 240.110 1864.670 ;
        RECT 238.930 1685.090 240.110 1686.270 ;
        RECT 238.930 1683.490 240.110 1684.670 ;
        RECT 238.930 1505.090 240.110 1506.270 ;
        RECT 238.930 1503.490 240.110 1504.670 ;
        RECT 238.930 1325.090 240.110 1326.270 ;
        RECT 238.930 1323.490 240.110 1324.670 ;
        RECT 238.930 1145.090 240.110 1146.270 ;
        RECT 238.930 1143.490 240.110 1144.670 ;
        RECT 238.930 965.090 240.110 966.270 ;
        RECT 238.930 963.490 240.110 964.670 ;
        RECT 238.930 785.090 240.110 786.270 ;
        RECT 238.930 783.490 240.110 784.670 ;
        RECT 238.930 605.090 240.110 606.270 ;
        RECT 238.930 603.490 240.110 604.670 ;
        RECT 238.930 425.090 240.110 426.270 ;
        RECT 238.930 423.490 240.110 424.670 ;
        RECT 238.930 245.090 240.110 246.270 ;
        RECT 238.930 243.490 240.110 244.670 ;
        RECT 238.930 65.090 240.110 66.270 ;
        RECT 238.930 63.490 240.110 64.670 ;
        RECT 238.930 -30.510 240.110 -29.330 ;
        RECT 238.930 -32.110 240.110 -30.930 ;
        RECT 418.930 3550.610 420.110 3551.790 ;
        RECT 418.930 3549.010 420.110 3550.190 ;
        RECT 418.930 3485.090 420.110 3486.270 ;
        RECT 418.930 3483.490 420.110 3484.670 ;
        RECT 418.930 3305.090 420.110 3306.270 ;
        RECT 418.930 3303.490 420.110 3304.670 ;
        RECT 418.930 3125.090 420.110 3126.270 ;
        RECT 418.930 3123.490 420.110 3124.670 ;
        RECT 418.930 2945.090 420.110 2946.270 ;
        RECT 418.930 2943.490 420.110 2944.670 ;
        RECT 418.930 2765.090 420.110 2766.270 ;
        RECT 418.930 2763.490 420.110 2764.670 ;
        RECT 418.930 2585.090 420.110 2586.270 ;
        RECT 418.930 2583.490 420.110 2584.670 ;
        RECT 418.930 2405.090 420.110 2406.270 ;
        RECT 418.930 2403.490 420.110 2404.670 ;
        RECT 418.930 2225.090 420.110 2226.270 ;
        RECT 418.930 2223.490 420.110 2224.670 ;
        RECT 418.930 2045.090 420.110 2046.270 ;
        RECT 418.930 2043.490 420.110 2044.670 ;
        RECT 418.930 1865.090 420.110 1866.270 ;
        RECT 418.930 1863.490 420.110 1864.670 ;
        RECT 418.930 1685.090 420.110 1686.270 ;
        RECT 418.930 1683.490 420.110 1684.670 ;
        RECT 418.930 1505.090 420.110 1506.270 ;
        RECT 418.930 1503.490 420.110 1504.670 ;
        RECT 418.930 1325.090 420.110 1326.270 ;
        RECT 418.930 1323.490 420.110 1324.670 ;
        RECT 418.930 1145.090 420.110 1146.270 ;
        RECT 418.930 1143.490 420.110 1144.670 ;
        RECT 418.930 965.090 420.110 966.270 ;
        RECT 418.930 963.490 420.110 964.670 ;
        RECT 418.930 785.090 420.110 786.270 ;
        RECT 418.930 783.490 420.110 784.670 ;
        RECT 418.930 605.090 420.110 606.270 ;
        RECT 418.930 603.490 420.110 604.670 ;
        RECT 418.930 425.090 420.110 426.270 ;
        RECT 418.930 423.490 420.110 424.670 ;
        RECT 418.930 245.090 420.110 246.270 ;
        RECT 418.930 243.490 420.110 244.670 ;
        RECT 418.930 65.090 420.110 66.270 ;
        RECT 418.930 63.490 420.110 64.670 ;
        RECT 418.930 -30.510 420.110 -29.330 ;
        RECT 418.930 -32.110 420.110 -30.930 ;
        RECT 598.930 3550.610 600.110 3551.790 ;
        RECT 598.930 3549.010 600.110 3550.190 ;
        RECT 598.930 3485.090 600.110 3486.270 ;
        RECT 598.930 3483.490 600.110 3484.670 ;
        RECT 598.930 3305.090 600.110 3306.270 ;
        RECT 598.930 3303.490 600.110 3304.670 ;
        RECT 598.930 3125.090 600.110 3126.270 ;
        RECT 598.930 3123.490 600.110 3124.670 ;
        RECT 598.930 2945.090 600.110 2946.270 ;
        RECT 598.930 2943.490 600.110 2944.670 ;
        RECT 598.930 2765.090 600.110 2766.270 ;
        RECT 598.930 2763.490 600.110 2764.670 ;
        RECT 598.930 2585.090 600.110 2586.270 ;
        RECT 598.930 2583.490 600.110 2584.670 ;
        RECT 598.930 2405.090 600.110 2406.270 ;
        RECT 598.930 2403.490 600.110 2404.670 ;
        RECT 598.930 2225.090 600.110 2226.270 ;
        RECT 598.930 2223.490 600.110 2224.670 ;
        RECT 598.930 2045.090 600.110 2046.270 ;
        RECT 598.930 2043.490 600.110 2044.670 ;
        RECT 598.930 1865.090 600.110 1866.270 ;
        RECT 598.930 1863.490 600.110 1864.670 ;
        RECT 598.930 1685.090 600.110 1686.270 ;
        RECT 598.930 1683.490 600.110 1684.670 ;
        RECT 598.930 1505.090 600.110 1506.270 ;
        RECT 598.930 1503.490 600.110 1504.670 ;
        RECT 598.930 1325.090 600.110 1326.270 ;
        RECT 598.930 1323.490 600.110 1324.670 ;
        RECT 598.930 1145.090 600.110 1146.270 ;
        RECT 598.930 1143.490 600.110 1144.670 ;
        RECT 598.930 965.090 600.110 966.270 ;
        RECT 598.930 963.490 600.110 964.670 ;
        RECT 598.930 785.090 600.110 786.270 ;
        RECT 598.930 783.490 600.110 784.670 ;
        RECT 598.930 605.090 600.110 606.270 ;
        RECT 598.930 603.490 600.110 604.670 ;
        RECT 598.930 425.090 600.110 426.270 ;
        RECT 598.930 423.490 600.110 424.670 ;
        RECT 598.930 245.090 600.110 246.270 ;
        RECT 598.930 243.490 600.110 244.670 ;
        RECT 598.930 65.090 600.110 66.270 ;
        RECT 598.930 63.490 600.110 64.670 ;
        RECT 598.930 -30.510 600.110 -29.330 ;
        RECT 598.930 -32.110 600.110 -30.930 ;
        RECT 778.930 3550.610 780.110 3551.790 ;
        RECT 778.930 3549.010 780.110 3550.190 ;
        RECT 778.930 3485.090 780.110 3486.270 ;
        RECT 778.930 3483.490 780.110 3484.670 ;
        RECT 778.930 3305.090 780.110 3306.270 ;
        RECT 778.930 3303.490 780.110 3304.670 ;
        RECT 778.930 3125.090 780.110 3126.270 ;
        RECT 778.930 3123.490 780.110 3124.670 ;
        RECT 778.930 2945.090 780.110 2946.270 ;
        RECT 778.930 2943.490 780.110 2944.670 ;
        RECT 778.930 2765.090 780.110 2766.270 ;
        RECT 778.930 2763.490 780.110 2764.670 ;
        RECT 778.930 2585.090 780.110 2586.270 ;
        RECT 778.930 2583.490 780.110 2584.670 ;
        RECT 778.930 2405.090 780.110 2406.270 ;
        RECT 778.930 2403.490 780.110 2404.670 ;
        RECT 778.930 2225.090 780.110 2226.270 ;
        RECT 778.930 2223.490 780.110 2224.670 ;
        RECT 778.930 2045.090 780.110 2046.270 ;
        RECT 778.930 2043.490 780.110 2044.670 ;
        RECT 778.930 1865.090 780.110 1866.270 ;
        RECT 778.930 1863.490 780.110 1864.670 ;
        RECT 778.930 1685.090 780.110 1686.270 ;
        RECT 778.930 1683.490 780.110 1684.670 ;
        RECT 778.930 1505.090 780.110 1506.270 ;
        RECT 778.930 1503.490 780.110 1504.670 ;
        RECT 778.930 1325.090 780.110 1326.270 ;
        RECT 778.930 1323.490 780.110 1324.670 ;
        RECT 778.930 1145.090 780.110 1146.270 ;
        RECT 778.930 1143.490 780.110 1144.670 ;
        RECT 778.930 965.090 780.110 966.270 ;
        RECT 778.930 963.490 780.110 964.670 ;
        RECT 778.930 785.090 780.110 786.270 ;
        RECT 778.930 783.490 780.110 784.670 ;
        RECT 778.930 605.090 780.110 606.270 ;
        RECT 778.930 603.490 780.110 604.670 ;
        RECT 778.930 425.090 780.110 426.270 ;
        RECT 778.930 423.490 780.110 424.670 ;
        RECT 778.930 245.090 780.110 246.270 ;
        RECT 778.930 243.490 780.110 244.670 ;
        RECT 778.930 65.090 780.110 66.270 ;
        RECT 778.930 63.490 780.110 64.670 ;
        RECT 778.930 -30.510 780.110 -29.330 ;
        RECT 778.930 -32.110 780.110 -30.930 ;
        RECT 958.930 3550.610 960.110 3551.790 ;
        RECT 958.930 3549.010 960.110 3550.190 ;
        RECT 958.930 3485.090 960.110 3486.270 ;
        RECT 958.930 3483.490 960.110 3484.670 ;
        RECT 958.930 3305.090 960.110 3306.270 ;
        RECT 958.930 3303.490 960.110 3304.670 ;
        RECT 958.930 3125.090 960.110 3126.270 ;
        RECT 958.930 3123.490 960.110 3124.670 ;
        RECT 958.930 2945.090 960.110 2946.270 ;
        RECT 958.930 2943.490 960.110 2944.670 ;
        RECT 958.930 2765.090 960.110 2766.270 ;
        RECT 958.930 2763.490 960.110 2764.670 ;
        RECT 958.930 2585.090 960.110 2586.270 ;
        RECT 958.930 2583.490 960.110 2584.670 ;
        RECT 958.930 2405.090 960.110 2406.270 ;
        RECT 958.930 2403.490 960.110 2404.670 ;
        RECT 958.930 2225.090 960.110 2226.270 ;
        RECT 958.930 2223.490 960.110 2224.670 ;
        RECT 958.930 2045.090 960.110 2046.270 ;
        RECT 958.930 2043.490 960.110 2044.670 ;
        RECT 958.930 1865.090 960.110 1866.270 ;
        RECT 958.930 1863.490 960.110 1864.670 ;
        RECT 958.930 1685.090 960.110 1686.270 ;
        RECT 958.930 1683.490 960.110 1684.670 ;
        RECT 958.930 1505.090 960.110 1506.270 ;
        RECT 958.930 1503.490 960.110 1504.670 ;
        RECT 958.930 1325.090 960.110 1326.270 ;
        RECT 958.930 1323.490 960.110 1324.670 ;
        RECT 958.930 1145.090 960.110 1146.270 ;
        RECT 958.930 1143.490 960.110 1144.670 ;
        RECT 958.930 965.090 960.110 966.270 ;
        RECT 958.930 963.490 960.110 964.670 ;
        RECT 958.930 785.090 960.110 786.270 ;
        RECT 958.930 783.490 960.110 784.670 ;
        RECT 958.930 605.090 960.110 606.270 ;
        RECT 958.930 603.490 960.110 604.670 ;
        RECT 958.930 425.090 960.110 426.270 ;
        RECT 958.930 423.490 960.110 424.670 ;
        RECT 958.930 245.090 960.110 246.270 ;
        RECT 958.930 243.490 960.110 244.670 ;
        RECT 958.930 65.090 960.110 66.270 ;
        RECT 958.930 63.490 960.110 64.670 ;
        RECT 958.930 -30.510 960.110 -29.330 ;
        RECT 958.930 -32.110 960.110 -30.930 ;
        RECT 1138.930 3550.610 1140.110 3551.790 ;
        RECT 1138.930 3549.010 1140.110 3550.190 ;
        RECT 1138.930 3485.090 1140.110 3486.270 ;
        RECT 1138.930 3483.490 1140.110 3484.670 ;
        RECT 1138.930 3305.090 1140.110 3306.270 ;
        RECT 1138.930 3303.490 1140.110 3304.670 ;
        RECT 1138.930 3125.090 1140.110 3126.270 ;
        RECT 1138.930 3123.490 1140.110 3124.670 ;
        RECT 1138.930 2945.090 1140.110 2946.270 ;
        RECT 1138.930 2943.490 1140.110 2944.670 ;
        RECT 1138.930 2765.090 1140.110 2766.270 ;
        RECT 1138.930 2763.490 1140.110 2764.670 ;
        RECT 1138.930 2585.090 1140.110 2586.270 ;
        RECT 1138.930 2583.490 1140.110 2584.670 ;
        RECT 1138.930 2405.090 1140.110 2406.270 ;
        RECT 1138.930 2403.490 1140.110 2404.670 ;
        RECT 1138.930 2225.090 1140.110 2226.270 ;
        RECT 1138.930 2223.490 1140.110 2224.670 ;
        RECT 1138.930 2045.090 1140.110 2046.270 ;
        RECT 1138.930 2043.490 1140.110 2044.670 ;
        RECT 1138.930 1865.090 1140.110 1866.270 ;
        RECT 1138.930 1863.490 1140.110 1864.670 ;
        RECT 1138.930 1685.090 1140.110 1686.270 ;
        RECT 1138.930 1683.490 1140.110 1684.670 ;
        RECT 1138.930 1505.090 1140.110 1506.270 ;
        RECT 1138.930 1503.490 1140.110 1504.670 ;
        RECT 1138.930 1325.090 1140.110 1326.270 ;
        RECT 1138.930 1323.490 1140.110 1324.670 ;
        RECT 1138.930 1145.090 1140.110 1146.270 ;
        RECT 1138.930 1143.490 1140.110 1144.670 ;
        RECT 1138.930 965.090 1140.110 966.270 ;
        RECT 1138.930 963.490 1140.110 964.670 ;
        RECT 1138.930 785.090 1140.110 786.270 ;
        RECT 1138.930 783.490 1140.110 784.670 ;
        RECT 1138.930 605.090 1140.110 606.270 ;
        RECT 1138.930 603.490 1140.110 604.670 ;
        RECT 1138.930 425.090 1140.110 426.270 ;
        RECT 1138.930 423.490 1140.110 424.670 ;
        RECT 1138.930 245.090 1140.110 246.270 ;
        RECT 1138.930 243.490 1140.110 244.670 ;
        RECT 1138.930 65.090 1140.110 66.270 ;
        RECT 1138.930 63.490 1140.110 64.670 ;
        RECT 1138.930 -30.510 1140.110 -29.330 ;
        RECT 1138.930 -32.110 1140.110 -30.930 ;
        RECT 1318.930 3550.610 1320.110 3551.790 ;
        RECT 1318.930 3549.010 1320.110 3550.190 ;
        RECT 1318.930 3485.090 1320.110 3486.270 ;
        RECT 1318.930 3483.490 1320.110 3484.670 ;
        RECT 1318.930 3305.090 1320.110 3306.270 ;
        RECT 1318.930 3303.490 1320.110 3304.670 ;
        RECT 1318.930 3125.090 1320.110 3126.270 ;
        RECT 1318.930 3123.490 1320.110 3124.670 ;
        RECT 1318.930 2945.090 1320.110 2946.270 ;
        RECT 1318.930 2943.490 1320.110 2944.670 ;
        RECT 1318.930 2765.090 1320.110 2766.270 ;
        RECT 1318.930 2763.490 1320.110 2764.670 ;
        RECT 1318.930 2585.090 1320.110 2586.270 ;
        RECT 1318.930 2583.490 1320.110 2584.670 ;
        RECT 1318.930 2405.090 1320.110 2406.270 ;
        RECT 1318.930 2403.490 1320.110 2404.670 ;
        RECT 1318.930 2225.090 1320.110 2226.270 ;
        RECT 1318.930 2223.490 1320.110 2224.670 ;
        RECT 1318.930 2045.090 1320.110 2046.270 ;
        RECT 1318.930 2043.490 1320.110 2044.670 ;
        RECT 1318.930 1865.090 1320.110 1866.270 ;
        RECT 1318.930 1863.490 1320.110 1864.670 ;
        RECT 1318.930 1685.090 1320.110 1686.270 ;
        RECT 1318.930 1683.490 1320.110 1684.670 ;
        RECT 1318.930 1505.090 1320.110 1506.270 ;
        RECT 1318.930 1503.490 1320.110 1504.670 ;
        RECT 1318.930 1325.090 1320.110 1326.270 ;
        RECT 1318.930 1323.490 1320.110 1324.670 ;
        RECT 1318.930 1145.090 1320.110 1146.270 ;
        RECT 1318.930 1143.490 1320.110 1144.670 ;
        RECT 1318.930 965.090 1320.110 966.270 ;
        RECT 1318.930 963.490 1320.110 964.670 ;
        RECT 1318.930 785.090 1320.110 786.270 ;
        RECT 1318.930 783.490 1320.110 784.670 ;
        RECT 1318.930 605.090 1320.110 606.270 ;
        RECT 1318.930 603.490 1320.110 604.670 ;
        RECT 1318.930 425.090 1320.110 426.270 ;
        RECT 1318.930 423.490 1320.110 424.670 ;
        RECT 1318.930 245.090 1320.110 246.270 ;
        RECT 1318.930 243.490 1320.110 244.670 ;
        RECT 1318.930 65.090 1320.110 66.270 ;
        RECT 1318.930 63.490 1320.110 64.670 ;
        RECT 1318.930 -30.510 1320.110 -29.330 ;
        RECT 1318.930 -32.110 1320.110 -30.930 ;
        RECT 1498.930 3550.610 1500.110 3551.790 ;
        RECT 1498.930 3549.010 1500.110 3550.190 ;
        RECT 1498.930 3485.090 1500.110 3486.270 ;
        RECT 1498.930 3483.490 1500.110 3484.670 ;
        RECT 1498.930 3305.090 1500.110 3306.270 ;
        RECT 1498.930 3303.490 1500.110 3304.670 ;
        RECT 1498.930 3125.090 1500.110 3126.270 ;
        RECT 1498.930 3123.490 1500.110 3124.670 ;
        RECT 1498.930 2945.090 1500.110 2946.270 ;
        RECT 1498.930 2943.490 1500.110 2944.670 ;
        RECT 1498.930 2765.090 1500.110 2766.270 ;
        RECT 1498.930 2763.490 1500.110 2764.670 ;
        RECT 1498.930 2585.090 1500.110 2586.270 ;
        RECT 1498.930 2583.490 1500.110 2584.670 ;
        RECT 1498.930 2405.090 1500.110 2406.270 ;
        RECT 1498.930 2403.490 1500.110 2404.670 ;
        RECT 1498.930 2225.090 1500.110 2226.270 ;
        RECT 1498.930 2223.490 1500.110 2224.670 ;
        RECT 1498.930 2045.090 1500.110 2046.270 ;
        RECT 1498.930 2043.490 1500.110 2044.670 ;
        RECT 1498.930 1865.090 1500.110 1866.270 ;
        RECT 1498.930 1863.490 1500.110 1864.670 ;
        RECT 1498.930 1685.090 1500.110 1686.270 ;
        RECT 1498.930 1683.490 1500.110 1684.670 ;
        RECT 1498.930 1505.090 1500.110 1506.270 ;
        RECT 1498.930 1503.490 1500.110 1504.670 ;
        RECT 1498.930 1325.090 1500.110 1326.270 ;
        RECT 1498.930 1323.490 1500.110 1324.670 ;
        RECT 1498.930 1145.090 1500.110 1146.270 ;
        RECT 1498.930 1143.490 1500.110 1144.670 ;
        RECT 1498.930 965.090 1500.110 966.270 ;
        RECT 1498.930 963.490 1500.110 964.670 ;
        RECT 1498.930 785.090 1500.110 786.270 ;
        RECT 1498.930 783.490 1500.110 784.670 ;
        RECT 1498.930 605.090 1500.110 606.270 ;
        RECT 1498.930 603.490 1500.110 604.670 ;
        RECT 1498.930 425.090 1500.110 426.270 ;
        RECT 1498.930 423.490 1500.110 424.670 ;
        RECT 1498.930 245.090 1500.110 246.270 ;
        RECT 1498.930 243.490 1500.110 244.670 ;
        RECT 1498.930 65.090 1500.110 66.270 ;
        RECT 1498.930 63.490 1500.110 64.670 ;
        RECT 1498.930 -30.510 1500.110 -29.330 ;
        RECT 1498.930 -32.110 1500.110 -30.930 ;
        RECT 1678.930 3550.610 1680.110 3551.790 ;
        RECT 1678.930 3549.010 1680.110 3550.190 ;
        RECT 1678.930 3485.090 1680.110 3486.270 ;
        RECT 1678.930 3483.490 1680.110 3484.670 ;
        RECT 1678.930 3305.090 1680.110 3306.270 ;
        RECT 1678.930 3303.490 1680.110 3304.670 ;
        RECT 1678.930 3125.090 1680.110 3126.270 ;
        RECT 1678.930 3123.490 1680.110 3124.670 ;
        RECT 1678.930 2945.090 1680.110 2946.270 ;
        RECT 1678.930 2943.490 1680.110 2944.670 ;
        RECT 1678.930 2765.090 1680.110 2766.270 ;
        RECT 1678.930 2763.490 1680.110 2764.670 ;
        RECT 1678.930 2585.090 1680.110 2586.270 ;
        RECT 1678.930 2583.490 1680.110 2584.670 ;
        RECT 1678.930 2405.090 1680.110 2406.270 ;
        RECT 1678.930 2403.490 1680.110 2404.670 ;
        RECT 1678.930 2225.090 1680.110 2226.270 ;
        RECT 1678.930 2223.490 1680.110 2224.670 ;
        RECT 1678.930 2045.090 1680.110 2046.270 ;
        RECT 1678.930 2043.490 1680.110 2044.670 ;
        RECT 1678.930 1865.090 1680.110 1866.270 ;
        RECT 1678.930 1863.490 1680.110 1864.670 ;
        RECT 1678.930 1685.090 1680.110 1686.270 ;
        RECT 1678.930 1683.490 1680.110 1684.670 ;
        RECT 1678.930 1505.090 1680.110 1506.270 ;
        RECT 1678.930 1503.490 1680.110 1504.670 ;
        RECT 1678.930 1325.090 1680.110 1326.270 ;
        RECT 1678.930 1323.490 1680.110 1324.670 ;
        RECT 1678.930 1145.090 1680.110 1146.270 ;
        RECT 1678.930 1143.490 1680.110 1144.670 ;
        RECT 1678.930 965.090 1680.110 966.270 ;
        RECT 1678.930 963.490 1680.110 964.670 ;
        RECT 1678.930 785.090 1680.110 786.270 ;
        RECT 1678.930 783.490 1680.110 784.670 ;
        RECT 1678.930 605.090 1680.110 606.270 ;
        RECT 1678.930 603.490 1680.110 604.670 ;
        RECT 1678.930 425.090 1680.110 426.270 ;
        RECT 1678.930 423.490 1680.110 424.670 ;
        RECT 1678.930 245.090 1680.110 246.270 ;
        RECT 1678.930 243.490 1680.110 244.670 ;
        RECT 1678.930 65.090 1680.110 66.270 ;
        RECT 1678.930 63.490 1680.110 64.670 ;
        RECT 1678.930 -30.510 1680.110 -29.330 ;
        RECT 1678.930 -32.110 1680.110 -30.930 ;
        RECT 1858.930 3550.610 1860.110 3551.790 ;
        RECT 1858.930 3549.010 1860.110 3550.190 ;
        RECT 1858.930 3485.090 1860.110 3486.270 ;
        RECT 1858.930 3483.490 1860.110 3484.670 ;
        RECT 1858.930 3305.090 1860.110 3306.270 ;
        RECT 1858.930 3303.490 1860.110 3304.670 ;
        RECT 1858.930 3125.090 1860.110 3126.270 ;
        RECT 1858.930 3123.490 1860.110 3124.670 ;
        RECT 1858.930 2945.090 1860.110 2946.270 ;
        RECT 1858.930 2943.490 1860.110 2944.670 ;
        RECT 1858.930 2765.090 1860.110 2766.270 ;
        RECT 1858.930 2763.490 1860.110 2764.670 ;
        RECT 1858.930 2585.090 1860.110 2586.270 ;
        RECT 1858.930 2583.490 1860.110 2584.670 ;
        RECT 1858.930 2405.090 1860.110 2406.270 ;
        RECT 1858.930 2403.490 1860.110 2404.670 ;
        RECT 1858.930 2225.090 1860.110 2226.270 ;
        RECT 1858.930 2223.490 1860.110 2224.670 ;
        RECT 1858.930 2045.090 1860.110 2046.270 ;
        RECT 1858.930 2043.490 1860.110 2044.670 ;
        RECT 1858.930 1865.090 1860.110 1866.270 ;
        RECT 1858.930 1863.490 1860.110 1864.670 ;
        RECT 1858.930 1685.090 1860.110 1686.270 ;
        RECT 1858.930 1683.490 1860.110 1684.670 ;
        RECT 1858.930 1505.090 1860.110 1506.270 ;
        RECT 1858.930 1503.490 1860.110 1504.670 ;
        RECT 1858.930 1325.090 1860.110 1326.270 ;
        RECT 1858.930 1323.490 1860.110 1324.670 ;
        RECT 1858.930 1145.090 1860.110 1146.270 ;
        RECT 1858.930 1143.490 1860.110 1144.670 ;
        RECT 1858.930 965.090 1860.110 966.270 ;
        RECT 1858.930 963.490 1860.110 964.670 ;
        RECT 1858.930 785.090 1860.110 786.270 ;
        RECT 1858.930 783.490 1860.110 784.670 ;
        RECT 1858.930 605.090 1860.110 606.270 ;
        RECT 1858.930 603.490 1860.110 604.670 ;
        RECT 1858.930 425.090 1860.110 426.270 ;
        RECT 1858.930 423.490 1860.110 424.670 ;
        RECT 1858.930 245.090 1860.110 246.270 ;
        RECT 1858.930 243.490 1860.110 244.670 ;
        RECT 1858.930 65.090 1860.110 66.270 ;
        RECT 1858.930 63.490 1860.110 64.670 ;
        RECT 1858.930 -30.510 1860.110 -29.330 ;
        RECT 1858.930 -32.110 1860.110 -30.930 ;
        RECT 2038.930 3550.610 2040.110 3551.790 ;
        RECT 2038.930 3549.010 2040.110 3550.190 ;
        RECT 2038.930 3485.090 2040.110 3486.270 ;
        RECT 2038.930 3483.490 2040.110 3484.670 ;
        RECT 2038.930 3305.090 2040.110 3306.270 ;
        RECT 2038.930 3303.490 2040.110 3304.670 ;
        RECT 2038.930 3125.090 2040.110 3126.270 ;
        RECT 2038.930 3123.490 2040.110 3124.670 ;
        RECT 2038.930 2945.090 2040.110 2946.270 ;
        RECT 2038.930 2943.490 2040.110 2944.670 ;
        RECT 2038.930 2765.090 2040.110 2766.270 ;
        RECT 2038.930 2763.490 2040.110 2764.670 ;
        RECT 2038.930 2585.090 2040.110 2586.270 ;
        RECT 2038.930 2583.490 2040.110 2584.670 ;
        RECT 2038.930 2405.090 2040.110 2406.270 ;
        RECT 2038.930 2403.490 2040.110 2404.670 ;
        RECT 2038.930 2225.090 2040.110 2226.270 ;
        RECT 2038.930 2223.490 2040.110 2224.670 ;
        RECT 2038.930 2045.090 2040.110 2046.270 ;
        RECT 2038.930 2043.490 2040.110 2044.670 ;
        RECT 2038.930 1865.090 2040.110 1866.270 ;
        RECT 2038.930 1863.490 2040.110 1864.670 ;
        RECT 2038.930 1685.090 2040.110 1686.270 ;
        RECT 2038.930 1683.490 2040.110 1684.670 ;
        RECT 2038.930 1505.090 2040.110 1506.270 ;
        RECT 2038.930 1503.490 2040.110 1504.670 ;
        RECT 2038.930 1325.090 2040.110 1326.270 ;
        RECT 2038.930 1323.490 2040.110 1324.670 ;
        RECT 2038.930 1145.090 2040.110 1146.270 ;
        RECT 2038.930 1143.490 2040.110 1144.670 ;
        RECT 2038.930 965.090 2040.110 966.270 ;
        RECT 2038.930 963.490 2040.110 964.670 ;
        RECT 2038.930 785.090 2040.110 786.270 ;
        RECT 2038.930 783.490 2040.110 784.670 ;
        RECT 2038.930 605.090 2040.110 606.270 ;
        RECT 2038.930 603.490 2040.110 604.670 ;
        RECT 2038.930 425.090 2040.110 426.270 ;
        RECT 2038.930 423.490 2040.110 424.670 ;
        RECT 2038.930 245.090 2040.110 246.270 ;
        RECT 2038.930 243.490 2040.110 244.670 ;
        RECT 2038.930 65.090 2040.110 66.270 ;
        RECT 2038.930 63.490 2040.110 64.670 ;
        RECT 2038.930 -30.510 2040.110 -29.330 ;
        RECT 2038.930 -32.110 2040.110 -30.930 ;
        RECT 2218.930 3550.610 2220.110 3551.790 ;
        RECT 2218.930 3549.010 2220.110 3550.190 ;
        RECT 2218.930 3485.090 2220.110 3486.270 ;
        RECT 2218.930 3483.490 2220.110 3484.670 ;
        RECT 2218.930 3305.090 2220.110 3306.270 ;
        RECT 2218.930 3303.490 2220.110 3304.670 ;
        RECT 2218.930 3125.090 2220.110 3126.270 ;
        RECT 2218.930 3123.490 2220.110 3124.670 ;
        RECT 2218.930 2945.090 2220.110 2946.270 ;
        RECT 2218.930 2943.490 2220.110 2944.670 ;
        RECT 2218.930 2765.090 2220.110 2766.270 ;
        RECT 2218.930 2763.490 2220.110 2764.670 ;
        RECT 2218.930 2585.090 2220.110 2586.270 ;
        RECT 2218.930 2583.490 2220.110 2584.670 ;
        RECT 2218.930 2405.090 2220.110 2406.270 ;
        RECT 2218.930 2403.490 2220.110 2404.670 ;
        RECT 2218.930 2225.090 2220.110 2226.270 ;
        RECT 2218.930 2223.490 2220.110 2224.670 ;
        RECT 2218.930 2045.090 2220.110 2046.270 ;
        RECT 2218.930 2043.490 2220.110 2044.670 ;
        RECT 2218.930 1865.090 2220.110 1866.270 ;
        RECT 2218.930 1863.490 2220.110 1864.670 ;
        RECT 2218.930 1685.090 2220.110 1686.270 ;
        RECT 2218.930 1683.490 2220.110 1684.670 ;
        RECT 2218.930 1505.090 2220.110 1506.270 ;
        RECT 2218.930 1503.490 2220.110 1504.670 ;
        RECT 2218.930 1325.090 2220.110 1326.270 ;
        RECT 2218.930 1323.490 2220.110 1324.670 ;
        RECT 2218.930 1145.090 2220.110 1146.270 ;
        RECT 2218.930 1143.490 2220.110 1144.670 ;
        RECT 2218.930 965.090 2220.110 966.270 ;
        RECT 2218.930 963.490 2220.110 964.670 ;
        RECT 2218.930 785.090 2220.110 786.270 ;
        RECT 2218.930 783.490 2220.110 784.670 ;
        RECT 2218.930 605.090 2220.110 606.270 ;
        RECT 2218.930 603.490 2220.110 604.670 ;
        RECT 2218.930 425.090 2220.110 426.270 ;
        RECT 2218.930 423.490 2220.110 424.670 ;
        RECT 2218.930 245.090 2220.110 246.270 ;
        RECT 2218.930 243.490 2220.110 244.670 ;
        RECT 2218.930 65.090 2220.110 66.270 ;
        RECT 2218.930 63.490 2220.110 64.670 ;
        RECT 2218.930 -30.510 2220.110 -29.330 ;
        RECT 2218.930 -32.110 2220.110 -30.930 ;
        RECT 2398.930 3550.610 2400.110 3551.790 ;
        RECT 2398.930 3549.010 2400.110 3550.190 ;
        RECT 2398.930 3485.090 2400.110 3486.270 ;
        RECT 2398.930 3483.490 2400.110 3484.670 ;
        RECT 2398.930 3305.090 2400.110 3306.270 ;
        RECT 2398.930 3303.490 2400.110 3304.670 ;
        RECT 2398.930 3125.090 2400.110 3126.270 ;
        RECT 2398.930 3123.490 2400.110 3124.670 ;
        RECT 2398.930 2945.090 2400.110 2946.270 ;
        RECT 2398.930 2943.490 2400.110 2944.670 ;
        RECT 2398.930 2765.090 2400.110 2766.270 ;
        RECT 2398.930 2763.490 2400.110 2764.670 ;
        RECT 2398.930 2585.090 2400.110 2586.270 ;
        RECT 2398.930 2583.490 2400.110 2584.670 ;
        RECT 2398.930 2405.090 2400.110 2406.270 ;
        RECT 2398.930 2403.490 2400.110 2404.670 ;
        RECT 2398.930 2225.090 2400.110 2226.270 ;
        RECT 2398.930 2223.490 2400.110 2224.670 ;
        RECT 2398.930 2045.090 2400.110 2046.270 ;
        RECT 2398.930 2043.490 2400.110 2044.670 ;
        RECT 2398.930 1865.090 2400.110 1866.270 ;
        RECT 2398.930 1863.490 2400.110 1864.670 ;
        RECT 2398.930 1685.090 2400.110 1686.270 ;
        RECT 2398.930 1683.490 2400.110 1684.670 ;
        RECT 2398.930 1505.090 2400.110 1506.270 ;
        RECT 2398.930 1503.490 2400.110 1504.670 ;
        RECT 2398.930 1325.090 2400.110 1326.270 ;
        RECT 2398.930 1323.490 2400.110 1324.670 ;
        RECT 2398.930 1145.090 2400.110 1146.270 ;
        RECT 2398.930 1143.490 2400.110 1144.670 ;
        RECT 2398.930 965.090 2400.110 966.270 ;
        RECT 2398.930 963.490 2400.110 964.670 ;
        RECT 2398.930 785.090 2400.110 786.270 ;
        RECT 2398.930 783.490 2400.110 784.670 ;
        RECT 2398.930 605.090 2400.110 606.270 ;
        RECT 2398.930 603.490 2400.110 604.670 ;
        RECT 2398.930 425.090 2400.110 426.270 ;
        RECT 2398.930 423.490 2400.110 424.670 ;
        RECT 2398.930 245.090 2400.110 246.270 ;
        RECT 2398.930 243.490 2400.110 244.670 ;
        RECT 2398.930 65.090 2400.110 66.270 ;
        RECT 2398.930 63.490 2400.110 64.670 ;
        RECT 2398.930 -30.510 2400.110 -29.330 ;
        RECT 2398.930 -32.110 2400.110 -30.930 ;
        RECT 2578.930 3550.610 2580.110 3551.790 ;
        RECT 2578.930 3549.010 2580.110 3550.190 ;
        RECT 2578.930 3485.090 2580.110 3486.270 ;
        RECT 2578.930 3483.490 2580.110 3484.670 ;
        RECT 2578.930 3305.090 2580.110 3306.270 ;
        RECT 2578.930 3303.490 2580.110 3304.670 ;
        RECT 2578.930 3125.090 2580.110 3126.270 ;
        RECT 2578.930 3123.490 2580.110 3124.670 ;
        RECT 2578.930 2945.090 2580.110 2946.270 ;
        RECT 2578.930 2943.490 2580.110 2944.670 ;
        RECT 2578.930 2765.090 2580.110 2766.270 ;
        RECT 2578.930 2763.490 2580.110 2764.670 ;
        RECT 2578.930 2585.090 2580.110 2586.270 ;
        RECT 2578.930 2583.490 2580.110 2584.670 ;
        RECT 2578.930 2405.090 2580.110 2406.270 ;
        RECT 2578.930 2403.490 2580.110 2404.670 ;
        RECT 2578.930 2225.090 2580.110 2226.270 ;
        RECT 2578.930 2223.490 2580.110 2224.670 ;
        RECT 2578.930 2045.090 2580.110 2046.270 ;
        RECT 2578.930 2043.490 2580.110 2044.670 ;
        RECT 2578.930 1865.090 2580.110 1866.270 ;
        RECT 2578.930 1863.490 2580.110 1864.670 ;
        RECT 2578.930 1685.090 2580.110 1686.270 ;
        RECT 2578.930 1683.490 2580.110 1684.670 ;
        RECT 2578.930 1505.090 2580.110 1506.270 ;
        RECT 2578.930 1503.490 2580.110 1504.670 ;
        RECT 2578.930 1325.090 2580.110 1326.270 ;
        RECT 2578.930 1323.490 2580.110 1324.670 ;
        RECT 2578.930 1145.090 2580.110 1146.270 ;
        RECT 2578.930 1143.490 2580.110 1144.670 ;
        RECT 2578.930 965.090 2580.110 966.270 ;
        RECT 2578.930 963.490 2580.110 964.670 ;
        RECT 2578.930 785.090 2580.110 786.270 ;
        RECT 2578.930 783.490 2580.110 784.670 ;
        RECT 2578.930 605.090 2580.110 606.270 ;
        RECT 2578.930 603.490 2580.110 604.670 ;
        RECT 2578.930 425.090 2580.110 426.270 ;
        RECT 2578.930 423.490 2580.110 424.670 ;
        RECT 2578.930 245.090 2580.110 246.270 ;
        RECT 2578.930 243.490 2580.110 244.670 ;
        RECT 2578.930 65.090 2580.110 66.270 ;
        RECT 2578.930 63.490 2580.110 64.670 ;
        RECT 2578.930 -30.510 2580.110 -29.330 ;
        RECT 2578.930 -32.110 2580.110 -30.930 ;
        RECT 2758.930 3550.610 2760.110 3551.790 ;
        RECT 2758.930 3549.010 2760.110 3550.190 ;
        RECT 2758.930 3485.090 2760.110 3486.270 ;
        RECT 2758.930 3483.490 2760.110 3484.670 ;
        RECT 2758.930 3305.090 2760.110 3306.270 ;
        RECT 2758.930 3303.490 2760.110 3304.670 ;
        RECT 2758.930 3125.090 2760.110 3126.270 ;
        RECT 2758.930 3123.490 2760.110 3124.670 ;
        RECT 2758.930 2945.090 2760.110 2946.270 ;
        RECT 2758.930 2943.490 2760.110 2944.670 ;
        RECT 2758.930 2765.090 2760.110 2766.270 ;
        RECT 2758.930 2763.490 2760.110 2764.670 ;
        RECT 2758.930 2585.090 2760.110 2586.270 ;
        RECT 2758.930 2583.490 2760.110 2584.670 ;
        RECT 2758.930 2405.090 2760.110 2406.270 ;
        RECT 2758.930 2403.490 2760.110 2404.670 ;
        RECT 2758.930 2225.090 2760.110 2226.270 ;
        RECT 2758.930 2223.490 2760.110 2224.670 ;
        RECT 2758.930 2045.090 2760.110 2046.270 ;
        RECT 2758.930 2043.490 2760.110 2044.670 ;
        RECT 2758.930 1865.090 2760.110 1866.270 ;
        RECT 2758.930 1863.490 2760.110 1864.670 ;
        RECT 2758.930 1685.090 2760.110 1686.270 ;
        RECT 2758.930 1683.490 2760.110 1684.670 ;
        RECT 2758.930 1505.090 2760.110 1506.270 ;
        RECT 2758.930 1503.490 2760.110 1504.670 ;
        RECT 2758.930 1325.090 2760.110 1326.270 ;
        RECT 2758.930 1323.490 2760.110 1324.670 ;
        RECT 2758.930 1145.090 2760.110 1146.270 ;
        RECT 2758.930 1143.490 2760.110 1144.670 ;
        RECT 2758.930 965.090 2760.110 966.270 ;
        RECT 2758.930 963.490 2760.110 964.670 ;
        RECT 2758.930 785.090 2760.110 786.270 ;
        RECT 2758.930 783.490 2760.110 784.670 ;
        RECT 2758.930 605.090 2760.110 606.270 ;
        RECT 2758.930 603.490 2760.110 604.670 ;
        RECT 2758.930 425.090 2760.110 426.270 ;
        RECT 2758.930 423.490 2760.110 424.670 ;
        RECT 2758.930 245.090 2760.110 246.270 ;
        RECT 2758.930 243.490 2760.110 244.670 ;
        RECT 2758.930 65.090 2760.110 66.270 ;
        RECT 2758.930 63.490 2760.110 64.670 ;
        RECT 2758.930 -30.510 2760.110 -29.330 ;
        RECT 2758.930 -32.110 2760.110 -30.930 ;
        RECT 2955.110 3550.610 2956.290 3551.790 ;
        RECT 2955.110 3549.010 2956.290 3550.190 ;
        RECT 2955.110 3485.090 2956.290 3486.270 ;
        RECT 2955.110 3483.490 2956.290 3484.670 ;
        RECT 2955.110 3305.090 2956.290 3306.270 ;
        RECT 2955.110 3303.490 2956.290 3304.670 ;
        RECT 2955.110 3125.090 2956.290 3126.270 ;
        RECT 2955.110 3123.490 2956.290 3124.670 ;
        RECT 2955.110 2945.090 2956.290 2946.270 ;
        RECT 2955.110 2943.490 2956.290 2944.670 ;
        RECT 2955.110 2765.090 2956.290 2766.270 ;
        RECT 2955.110 2763.490 2956.290 2764.670 ;
        RECT 2955.110 2585.090 2956.290 2586.270 ;
        RECT 2955.110 2583.490 2956.290 2584.670 ;
        RECT 2955.110 2405.090 2956.290 2406.270 ;
        RECT 2955.110 2403.490 2956.290 2404.670 ;
        RECT 2955.110 2225.090 2956.290 2226.270 ;
        RECT 2955.110 2223.490 2956.290 2224.670 ;
        RECT 2955.110 2045.090 2956.290 2046.270 ;
        RECT 2955.110 2043.490 2956.290 2044.670 ;
        RECT 2955.110 1865.090 2956.290 1866.270 ;
        RECT 2955.110 1863.490 2956.290 1864.670 ;
        RECT 2955.110 1685.090 2956.290 1686.270 ;
        RECT 2955.110 1683.490 2956.290 1684.670 ;
        RECT 2955.110 1505.090 2956.290 1506.270 ;
        RECT 2955.110 1503.490 2956.290 1504.670 ;
        RECT 2955.110 1325.090 2956.290 1326.270 ;
        RECT 2955.110 1323.490 2956.290 1324.670 ;
        RECT 2955.110 1145.090 2956.290 1146.270 ;
        RECT 2955.110 1143.490 2956.290 1144.670 ;
        RECT 2955.110 965.090 2956.290 966.270 ;
        RECT 2955.110 963.490 2956.290 964.670 ;
        RECT 2955.110 785.090 2956.290 786.270 ;
        RECT 2955.110 783.490 2956.290 784.670 ;
        RECT 2955.110 605.090 2956.290 606.270 ;
        RECT 2955.110 603.490 2956.290 604.670 ;
        RECT 2955.110 425.090 2956.290 426.270 ;
        RECT 2955.110 423.490 2956.290 424.670 ;
        RECT 2955.110 245.090 2956.290 246.270 ;
        RECT 2955.110 243.490 2956.290 244.670 ;
        RECT 2955.110 65.090 2956.290 66.270 ;
        RECT 2955.110 63.490 2956.290 64.670 ;
        RECT 2955.110 -30.510 2956.290 -29.330 ;
        RECT 2955.110 -32.110 2956.290 -30.930 ;
      LAYER met5 ;
        RECT -37.580 3551.900 -34.580 3551.910 ;
        RECT 58.020 3551.900 61.020 3551.910 ;
        RECT 238.020 3551.900 241.020 3551.910 ;
        RECT 418.020 3551.900 421.020 3551.910 ;
        RECT 598.020 3551.900 601.020 3551.910 ;
        RECT 778.020 3551.900 781.020 3551.910 ;
        RECT 958.020 3551.900 961.020 3551.910 ;
        RECT 1138.020 3551.900 1141.020 3551.910 ;
        RECT 1318.020 3551.900 1321.020 3551.910 ;
        RECT 1498.020 3551.900 1501.020 3551.910 ;
        RECT 1678.020 3551.900 1681.020 3551.910 ;
        RECT 1858.020 3551.900 1861.020 3551.910 ;
        RECT 2038.020 3551.900 2041.020 3551.910 ;
        RECT 2218.020 3551.900 2221.020 3551.910 ;
        RECT 2398.020 3551.900 2401.020 3551.910 ;
        RECT 2578.020 3551.900 2581.020 3551.910 ;
        RECT 2758.020 3551.900 2761.020 3551.910 ;
        RECT 2954.200 3551.900 2957.200 3551.910 ;
        RECT -37.580 3548.900 2957.200 3551.900 ;
        RECT -37.580 3548.890 -34.580 3548.900 ;
        RECT 58.020 3548.890 61.020 3548.900 ;
        RECT 238.020 3548.890 241.020 3548.900 ;
        RECT 418.020 3548.890 421.020 3548.900 ;
        RECT 598.020 3548.890 601.020 3548.900 ;
        RECT 778.020 3548.890 781.020 3548.900 ;
        RECT 958.020 3548.890 961.020 3548.900 ;
        RECT 1138.020 3548.890 1141.020 3548.900 ;
        RECT 1318.020 3548.890 1321.020 3548.900 ;
        RECT 1498.020 3548.890 1501.020 3548.900 ;
        RECT 1678.020 3548.890 1681.020 3548.900 ;
        RECT 1858.020 3548.890 1861.020 3548.900 ;
        RECT 2038.020 3548.890 2041.020 3548.900 ;
        RECT 2218.020 3548.890 2221.020 3548.900 ;
        RECT 2398.020 3548.890 2401.020 3548.900 ;
        RECT 2578.020 3548.890 2581.020 3548.900 ;
        RECT 2758.020 3548.890 2761.020 3548.900 ;
        RECT 2954.200 3548.890 2957.200 3548.900 ;
        RECT -37.580 3486.380 -34.580 3486.390 ;
        RECT 58.020 3486.380 61.020 3486.390 ;
        RECT 238.020 3486.380 241.020 3486.390 ;
        RECT 418.020 3486.380 421.020 3486.390 ;
        RECT 598.020 3486.380 601.020 3486.390 ;
        RECT 778.020 3486.380 781.020 3486.390 ;
        RECT 958.020 3486.380 961.020 3486.390 ;
        RECT 1138.020 3486.380 1141.020 3486.390 ;
        RECT 1318.020 3486.380 1321.020 3486.390 ;
        RECT 1498.020 3486.380 1501.020 3486.390 ;
        RECT 1678.020 3486.380 1681.020 3486.390 ;
        RECT 1858.020 3486.380 1861.020 3486.390 ;
        RECT 2038.020 3486.380 2041.020 3486.390 ;
        RECT 2218.020 3486.380 2221.020 3486.390 ;
        RECT 2398.020 3486.380 2401.020 3486.390 ;
        RECT 2578.020 3486.380 2581.020 3486.390 ;
        RECT 2758.020 3486.380 2761.020 3486.390 ;
        RECT 2954.200 3486.380 2957.200 3486.390 ;
        RECT -42.180 3483.380 2961.800 3486.380 ;
        RECT -37.580 3483.370 -34.580 3483.380 ;
        RECT 58.020 3483.370 61.020 3483.380 ;
        RECT 238.020 3483.370 241.020 3483.380 ;
        RECT 418.020 3483.370 421.020 3483.380 ;
        RECT 598.020 3483.370 601.020 3483.380 ;
        RECT 778.020 3483.370 781.020 3483.380 ;
        RECT 958.020 3483.370 961.020 3483.380 ;
        RECT 1138.020 3483.370 1141.020 3483.380 ;
        RECT 1318.020 3483.370 1321.020 3483.380 ;
        RECT 1498.020 3483.370 1501.020 3483.380 ;
        RECT 1678.020 3483.370 1681.020 3483.380 ;
        RECT 1858.020 3483.370 1861.020 3483.380 ;
        RECT 2038.020 3483.370 2041.020 3483.380 ;
        RECT 2218.020 3483.370 2221.020 3483.380 ;
        RECT 2398.020 3483.370 2401.020 3483.380 ;
        RECT 2578.020 3483.370 2581.020 3483.380 ;
        RECT 2758.020 3483.370 2761.020 3483.380 ;
        RECT 2954.200 3483.370 2957.200 3483.380 ;
        RECT -37.580 3306.380 -34.580 3306.390 ;
        RECT 58.020 3306.380 61.020 3306.390 ;
        RECT 238.020 3306.380 241.020 3306.390 ;
        RECT 418.020 3306.380 421.020 3306.390 ;
        RECT 598.020 3306.380 601.020 3306.390 ;
        RECT 778.020 3306.380 781.020 3306.390 ;
        RECT 958.020 3306.380 961.020 3306.390 ;
        RECT 1138.020 3306.380 1141.020 3306.390 ;
        RECT 1318.020 3306.380 1321.020 3306.390 ;
        RECT 1498.020 3306.380 1501.020 3306.390 ;
        RECT 1678.020 3306.380 1681.020 3306.390 ;
        RECT 1858.020 3306.380 1861.020 3306.390 ;
        RECT 2038.020 3306.380 2041.020 3306.390 ;
        RECT 2218.020 3306.380 2221.020 3306.390 ;
        RECT 2398.020 3306.380 2401.020 3306.390 ;
        RECT 2578.020 3306.380 2581.020 3306.390 ;
        RECT 2758.020 3306.380 2761.020 3306.390 ;
        RECT 2954.200 3306.380 2957.200 3306.390 ;
        RECT -42.180 3303.380 2961.800 3306.380 ;
        RECT -37.580 3303.370 -34.580 3303.380 ;
        RECT 58.020 3303.370 61.020 3303.380 ;
        RECT 238.020 3303.370 241.020 3303.380 ;
        RECT 418.020 3303.370 421.020 3303.380 ;
        RECT 598.020 3303.370 601.020 3303.380 ;
        RECT 778.020 3303.370 781.020 3303.380 ;
        RECT 958.020 3303.370 961.020 3303.380 ;
        RECT 1138.020 3303.370 1141.020 3303.380 ;
        RECT 1318.020 3303.370 1321.020 3303.380 ;
        RECT 1498.020 3303.370 1501.020 3303.380 ;
        RECT 1678.020 3303.370 1681.020 3303.380 ;
        RECT 1858.020 3303.370 1861.020 3303.380 ;
        RECT 2038.020 3303.370 2041.020 3303.380 ;
        RECT 2218.020 3303.370 2221.020 3303.380 ;
        RECT 2398.020 3303.370 2401.020 3303.380 ;
        RECT 2578.020 3303.370 2581.020 3303.380 ;
        RECT 2758.020 3303.370 2761.020 3303.380 ;
        RECT 2954.200 3303.370 2957.200 3303.380 ;
        RECT -37.580 3126.380 -34.580 3126.390 ;
        RECT 58.020 3126.380 61.020 3126.390 ;
        RECT 238.020 3126.380 241.020 3126.390 ;
        RECT 418.020 3126.380 421.020 3126.390 ;
        RECT 598.020 3126.380 601.020 3126.390 ;
        RECT 778.020 3126.380 781.020 3126.390 ;
        RECT 958.020 3126.380 961.020 3126.390 ;
        RECT 1138.020 3126.380 1141.020 3126.390 ;
        RECT 1318.020 3126.380 1321.020 3126.390 ;
        RECT 1498.020 3126.380 1501.020 3126.390 ;
        RECT 1678.020 3126.380 1681.020 3126.390 ;
        RECT 1858.020 3126.380 1861.020 3126.390 ;
        RECT 2038.020 3126.380 2041.020 3126.390 ;
        RECT 2218.020 3126.380 2221.020 3126.390 ;
        RECT 2398.020 3126.380 2401.020 3126.390 ;
        RECT 2578.020 3126.380 2581.020 3126.390 ;
        RECT 2758.020 3126.380 2761.020 3126.390 ;
        RECT 2954.200 3126.380 2957.200 3126.390 ;
        RECT -42.180 3123.380 2961.800 3126.380 ;
        RECT -37.580 3123.370 -34.580 3123.380 ;
        RECT 58.020 3123.370 61.020 3123.380 ;
        RECT 238.020 3123.370 241.020 3123.380 ;
        RECT 418.020 3123.370 421.020 3123.380 ;
        RECT 598.020 3123.370 601.020 3123.380 ;
        RECT 778.020 3123.370 781.020 3123.380 ;
        RECT 958.020 3123.370 961.020 3123.380 ;
        RECT 1138.020 3123.370 1141.020 3123.380 ;
        RECT 1318.020 3123.370 1321.020 3123.380 ;
        RECT 1498.020 3123.370 1501.020 3123.380 ;
        RECT 1678.020 3123.370 1681.020 3123.380 ;
        RECT 1858.020 3123.370 1861.020 3123.380 ;
        RECT 2038.020 3123.370 2041.020 3123.380 ;
        RECT 2218.020 3123.370 2221.020 3123.380 ;
        RECT 2398.020 3123.370 2401.020 3123.380 ;
        RECT 2578.020 3123.370 2581.020 3123.380 ;
        RECT 2758.020 3123.370 2761.020 3123.380 ;
        RECT 2954.200 3123.370 2957.200 3123.380 ;
        RECT -37.580 2946.380 -34.580 2946.390 ;
        RECT 58.020 2946.380 61.020 2946.390 ;
        RECT 238.020 2946.380 241.020 2946.390 ;
        RECT 418.020 2946.380 421.020 2946.390 ;
        RECT 598.020 2946.380 601.020 2946.390 ;
        RECT 778.020 2946.380 781.020 2946.390 ;
        RECT 958.020 2946.380 961.020 2946.390 ;
        RECT 1138.020 2946.380 1141.020 2946.390 ;
        RECT 1318.020 2946.380 1321.020 2946.390 ;
        RECT 1498.020 2946.380 1501.020 2946.390 ;
        RECT 1678.020 2946.380 1681.020 2946.390 ;
        RECT 1858.020 2946.380 1861.020 2946.390 ;
        RECT 2038.020 2946.380 2041.020 2946.390 ;
        RECT 2218.020 2946.380 2221.020 2946.390 ;
        RECT 2398.020 2946.380 2401.020 2946.390 ;
        RECT 2578.020 2946.380 2581.020 2946.390 ;
        RECT 2758.020 2946.380 2761.020 2946.390 ;
        RECT 2954.200 2946.380 2957.200 2946.390 ;
        RECT -42.180 2943.380 2961.800 2946.380 ;
        RECT -37.580 2943.370 -34.580 2943.380 ;
        RECT 58.020 2943.370 61.020 2943.380 ;
        RECT 238.020 2943.370 241.020 2943.380 ;
        RECT 418.020 2943.370 421.020 2943.380 ;
        RECT 598.020 2943.370 601.020 2943.380 ;
        RECT 778.020 2943.370 781.020 2943.380 ;
        RECT 958.020 2943.370 961.020 2943.380 ;
        RECT 1138.020 2943.370 1141.020 2943.380 ;
        RECT 1318.020 2943.370 1321.020 2943.380 ;
        RECT 1498.020 2943.370 1501.020 2943.380 ;
        RECT 1678.020 2943.370 1681.020 2943.380 ;
        RECT 1858.020 2943.370 1861.020 2943.380 ;
        RECT 2038.020 2943.370 2041.020 2943.380 ;
        RECT 2218.020 2943.370 2221.020 2943.380 ;
        RECT 2398.020 2943.370 2401.020 2943.380 ;
        RECT 2578.020 2943.370 2581.020 2943.380 ;
        RECT 2758.020 2943.370 2761.020 2943.380 ;
        RECT 2954.200 2943.370 2957.200 2943.380 ;
        RECT -37.580 2766.380 -34.580 2766.390 ;
        RECT 58.020 2766.380 61.020 2766.390 ;
        RECT 238.020 2766.380 241.020 2766.390 ;
        RECT 418.020 2766.380 421.020 2766.390 ;
        RECT 598.020 2766.380 601.020 2766.390 ;
        RECT 778.020 2766.380 781.020 2766.390 ;
        RECT 958.020 2766.380 961.020 2766.390 ;
        RECT 1138.020 2766.380 1141.020 2766.390 ;
        RECT 1318.020 2766.380 1321.020 2766.390 ;
        RECT 1498.020 2766.380 1501.020 2766.390 ;
        RECT 1678.020 2766.380 1681.020 2766.390 ;
        RECT 1858.020 2766.380 1861.020 2766.390 ;
        RECT 2038.020 2766.380 2041.020 2766.390 ;
        RECT 2218.020 2766.380 2221.020 2766.390 ;
        RECT 2398.020 2766.380 2401.020 2766.390 ;
        RECT 2578.020 2766.380 2581.020 2766.390 ;
        RECT 2758.020 2766.380 2761.020 2766.390 ;
        RECT 2954.200 2766.380 2957.200 2766.390 ;
        RECT -42.180 2763.380 2961.800 2766.380 ;
        RECT -37.580 2763.370 -34.580 2763.380 ;
        RECT 58.020 2763.370 61.020 2763.380 ;
        RECT 238.020 2763.370 241.020 2763.380 ;
        RECT 418.020 2763.370 421.020 2763.380 ;
        RECT 598.020 2763.370 601.020 2763.380 ;
        RECT 778.020 2763.370 781.020 2763.380 ;
        RECT 958.020 2763.370 961.020 2763.380 ;
        RECT 1138.020 2763.370 1141.020 2763.380 ;
        RECT 1318.020 2763.370 1321.020 2763.380 ;
        RECT 1498.020 2763.370 1501.020 2763.380 ;
        RECT 1678.020 2763.370 1681.020 2763.380 ;
        RECT 1858.020 2763.370 1861.020 2763.380 ;
        RECT 2038.020 2763.370 2041.020 2763.380 ;
        RECT 2218.020 2763.370 2221.020 2763.380 ;
        RECT 2398.020 2763.370 2401.020 2763.380 ;
        RECT 2578.020 2763.370 2581.020 2763.380 ;
        RECT 2758.020 2763.370 2761.020 2763.380 ;
        RECT 2954.200 2763.370 2957.200 2763.380 ;
        RECT -37.580 2586.380 -34.580 2586.390 ;
        RECT 58.020 2586.380 61.020 2586.390 ;
        RECT 238.020 2586.380 241.020 2586.390 ;
        RECT 418.020 2586.380 421.020 2586.390 ;
        RECT 598.020 2586.380 601.020 2586.390 ;
        RECT 778.020 2586.380 781.020 2586.390 ;
        RECT 958.020 2586.380 961.020 2586.390 ;
        RECT 1138.020 2586.380 1141.020 2586.390 ;
        RECT 1318.020 2586.380 1321.020 2586.390 ;
        RECT 1498.020 2586.380 1501.020 2586.390 ;
        RECT 1678.020 2586.380 1681.020 2586.390 ;
        RECT 1858.020 2586.380 1861.020 2586.390 ;
        RECT 2038.020 2586.380 2041.020 2586.390 ;
        RECT 2218.020 2586.380 2221.020 2586.390 ;
        RECT 2398.020 2586.380 2401.020 2586.390 ;
        RECT 2578.020 2586.380 2581.020 2586.390 ;
        RECT 2758.020 2586.380 2761.020 2586.390 ;
        RECT 2954.200 2586.380 2957.200 2586.390 ;
        RECT -42.180 2583.380 2961.800 2586.380 ;
        RECT -37.580 2583.370 -34.580 2583.380 ;
        RECT 58.020 2583.370 61.020 2583.380 ;
        RECT 238.020 2583.370 241.020 2583.380 ;
        RECT 418.020 2583.370 421.020 2583.380 ;
        RECT 598.020 2583.370 601.020 2583.380 ;
        RECT 778.020 2583.370 781.020 2583.380 ;
        RECT 958.020 2583.370 961.020 2583.380 ;
        RECT 1138.020 2583.370 1141.020 2583.380 ;
        RECT 1318.020 2583.370 1321.020 2583.380 ;
        RECT 1498.020 2583.370 1501.020 2583.380 ;
        RECT 1678.020 2583.370 1681.020 2583.380 ;
        RECT 1858.020 2583.370 1861.020 2583.380 ;
        RECT 2038.020 2583.370 2041.020 2583.380 ;
        RECT 2218.020 2583.370 2221.020 2583.380 ;
        RECT 2398.020 2583.370 2401.020 2583.380 ;
        RECT 2578.020 2583.370 2581.020 2583.380 ;
        RECT 2758.020 2583.370 2761.020 2583.380 ;
        RECT 2954.200 2583.370 2957.200 2583.380 ;
        RECT -37.580 2406.380 -34.580 2406.390 ;
        RECT 58.020 2406.380 61.020 2406.390 ;
        RECT 238.020 2406.380 241.020 2406.390 ;
        RECT 418.020 2406.380 421.020 2406.390 ;
        RECT 598.020 2406.380 601.020 2406.390 ;
        RECT 778.020 2406.380 781.020 2406.390 ;
        RECT 958.020 2406.380 961.020 2406.390 ;
        RECT 1138.020 2406.380 1141.020 2406.390 ;
        RECT 1318.020 2406.380 1321.020 2406.390 ;
        RECT 1498.020 2406.380 1501.020 2406.390 ;
        RECT 1678.020 2406.380 1681.020 2406.390 ;
        RECT 1858.020 2406.380 1861.020 2406.390 ;
        RECT 2038.020 2406.380 2041.020 2406.390 ;
        RECT 2218.020 2406.380 2221.020 2406.390 ;
        RECT 2398.020 2406.380 2401.020 2406.390 ;
        RECT 2578.020 2406.380 2581.020 2406.390 ;
        RECT 2758.020 2406.380 2761.020 2406.390 ;
        RECT 2954.200 2406.380 2957.200 2406.390 ;
        RECT -42.180 2403.380 2961.800 2406.380 ;
        RECT -37.580 2403.370 -34.580 2403.380 ;
        RECT 58.020 2403.370 61.020 2403.380 ;
        RECT 238.020 2403.370 241.020 2403.380 ;
        RECT 418.020 2403.370 421.020 2403.380 ;
        RECT 598.020 2403.370 601.020 2403.380 ;
        RECT 778.020 2403.370 781.020 2403.380 ;
        RECT 958.020 2403.370 961.020 2403.380 ;
        RECT 1138.020 2403.370 1141.020 2403.380 ;
        RECT 1318.020 2403.370 1321.020 2403.380 ;
        RECT 1498.020 2403.370 1501.020 2403.380 ;
        RECT 1678.020 2403.370 1681.020 2403.380 ;
        RECT 1858.020 2403.370 1861.020 2403.380 ;
        RECT 2038.020 2403.370 2041.020 2403.380 ;
        RECT 2218.020 2403.370 2221.020 2403.380 ;
        RECT 2398.020 2403.370 2401.020 2403.380 ;
        RECT 2578.020 2403.370 2581.020 2403.380 ;
        RECT 2758.020 2403.370 2761.020 2403.380 ;
        RECT 2954.200 2403.370 2957.200 2403.380 ;
        RECT -37.580 2226.380 -34.580 2226.390 ;
        RECT 58.020 2226.380 61.020 2226.390 ;
        RECT 238.020 2226.380 241.020 2226.390 ;
        RECT 418.020 2226.380 421.020 2226.390 ;
        RECT 598.020 2226.380 601.020 2226.390 ;
        RECT 778.020 2226.380 781.020 2226.390 ;
        RECT 958.020 2226.380 961.020 2226.390 ;
        RECT 1138.020 2226.380 1141.020 2226.390 ;
        RECT 1318.020 2226.380 1321.020 2226.390 ;
        RECT 1498.020 2226.380 1501.020 2226.390 ;
        RECT 1678.020 2226.380 1681.020 2226.390 ;
        RECT 1858.020 2226.380 1861.020 2226.390 ;
        RECT 2038.020 2226.380 2041.020 2226.390 ;
        RECT 2218.020 2226.380 2221.020 2226.390 ;
        RECT 2398.020 2226.380 2401.020 2226.390 ;
        RECT 2578.020 2226.380 2581.020 2226.390 ;
        RECT 2758.020 2226.380 2761.020 2226.390 ;
        RECT 2954.200 2226.380 2957.200 2226.390 ;
        RECT -42.180 2223.380 2961.800 2226.380 ;
        RECT -37.580 2223.370 -34.580 2223.380 ;
        RECT 58.020 2223.370 61.020 2223.380 ;
        RECT 238.020 2223.370 241.020 2223.380 ;
        RECT 418.020 2223.370 421.020 2223.380 ;
        RECT 598.020 2223.370 601.020 2223.380 ;
        RECT 778.020 2223.370 781.020 2223.380 ;
        RECT 958.020 2223.370 961.020 2223.380 ;
        RECT 1138.020 2223.370 1141.020 2223.380 ;
        RECT 1318.020 2223.370 1321.020 2223.380 ;
        RECT 1498.020 2223.370 1501.020 2223.380 ;
        RECT 1678.020 2223.370 1681.020 2223.380 ;
        RECT 1858.020 2223.370 1861.020 2223.380 ;
        RECT 2038.020 2223.370 2041.020 2223.380 ;
        RECT 2218.020 2223.370 2221.020 2223.380 ;
        RECT 2398.020 2223.370 2401.020 2223.380 ;
        RECT 2578.020 2223.370 2581.020 2223.380 ;
        RECT 2758.020 2223.370 2761.020 2223.380 ;
        RECT 2954.200 2223.370 2957.200 2223.380 ;
        RECT -37.580 2046.380 -34.580 2046.390 ;
        RECT 58.020 2046.380 61.020 2046.390 ;
        RECT 238.020 2046.380 241.020 2046.390 ;
        RECT 418.020 2046.380 421.020 2046.390 ;
        RECT 598.020 2046.380 601.020 2046.390 ;
        RECT 778.020 2046.380 781.020 2046.390 ;
        RECT 958.020 2046.380 961.020 2046.390 ;
        RECT 1138.020 2046.380 1141.020 2046.390 ;
        RECT 1318.020 2046.380 1321.020 2046.390 ;
        RECT 1498.020 2046.380 1501.020 2046.390 ;
        RECT 1678.020 2046.380 1681.020 2046.390 ;
        RECT 1858.020 2046.380 1861.020 2046.390 ;
        RECT 2038.020 2046.380 2041.020 2046.390 ;
        RECT 2218.020 2046.380 2221.020 2046.390 ;
        RECT 2398.020 2046.380 2401.020 2046.390 ;
        RECT 2578.020 2046.380 2581.020 2046.390 ;
        RECT 2758.020 2046.380 2761.020 2046.390 ;
        RECT 2954.200 2046.380 2957.200 2046.390 ;
        RECT -42.180 2043.380 2961.800 2046.380 ;
        RECT -37.580 2043.370 -34.580 2043.380 ;
        RECT 58.020 2043.370 61.020 2043.380 ;
        RECT 238.020 2043.370 241.020 2043.380 ;
        RECT 418.020 2043.370 421.020 2043.380 ;
        RECT 598.020 2043.370 601.020 2043.380 ;
        RECT 778.020 2043.370 781.020 2043.380 ;
        RECT 958.020 2043.370 961.020 2043.380 ;
        RECT 1138.020 2043.370 1141.020 2043.380 ;
        RECT 1318.020 2043.370 1321.020 2043.380 ;
        RECT 1498.020 2043.370 1501.020 2043.380 ;
        RECT 1678.020 2043.370 1681.020 2043.380 ;
        RECT 1858.020 2043.370 1861.020 2043.380 ;
        RECT 2038.020 2043.370 2041.020 2043.380 ;
        RECT 2218.020 2043.370 2221.020 2043.380 ;
        RECT 2398.020 2043.370 2401.020 2043.380 ;
        RECT 2578.020 2043.370 2581.020 2043.380 ;
        RECT 2758.020 2043.370 2761.020 2043.380 ;
        RECT 2954.200 2043.370 2957.200 2043.380 ;
        RECT -37.580 1866.380 -34.580 1866.390 ;
        RECT 58.020 1866.380 61.020 1866.390 ;
        RECT 238.020 1866.380 241.020 1866.390 ;
        RECT 418.020 1866.380 421.020 1866.390 ;
        RECT 598.020 1866.380 601.020 1866.390 ;
        RECT 778.020 1866.380 781.020 1866.390 ;
        RECT 958.020 1866.380 961.020 1866.390 ;
        RECT 1138.020 1866.380 1141.020 1866.390 ;
        RECT 1318.020 1866.380 1321.020 1866.390 ;
        RECT 1498.020 1866.380 1501.020 1866.390 ;
        RECT 1678.020 1866.380 1681.020 1866.390 ;
        RECT 1858.020 1866.380 1861.020 1866.390 ;
        RECT 2038.020 1866.380 2041.020 1866.390 ;
        RECT 2218.020 1866.380 2221.020 1866.390 ;
        RECT 2398.020 1866.380 2401.020 1866.390 ;
        RECT 2578.020 1866.380 2581.020 1866.390 ;
        RECT 2758.020 1866.380 2761.020 1866.390 ;
        RECT 2954.200 1866.380 2957.200 1866.390 ;
        RECT -42.180 1863.380 2961.800 1866.380 ;
        RECT -37.580 1863.370 -34.580 1863.380 ;
        RECT 58.020 1863.370 61.020 1863.380 ;
        RECT 238.020 1863.370 241.020 1863.380 ;
        RECT 418.020 1863.370 421.020 1863.380 ;
        RECT 598.020 1863.370 601.020 1863.380 ;
        RECT 778.020 1863.370 781.020 1863.380 ;
        RECT 958.020 1863.370 961.020 1863.380 ;
        RECT 1138.020 1863.370 1141.020 1863.380 ;
        RECT 1318.020 1863.370 1321.020 1863.380 ;
        RECT 1498.020 1863.370 1501.020 1863.380 ;
        RECT 1678.020 1863.370 1681.020 1863.380 ;
        RECT 1858.020 1863.370 1861.020 1863.380 ;
        RECT 2038.020 1863.370 2041.020 1863.380 ;
        RECT 2218.020 1863.370 2221.020 1863.380 ;
        RECT 2398.020 1863.370 2401.020 1863.380 ;
        RECT 2578.020 1863.370 2581.020 1863.380 ;
        RECT 2758.020 1863.370 2761.020 1863.380 ;
        RECT 2954.200 1863.370 2957.200 1863.380 ;
        RECT -37.580 1686.380 -34.580 1686.390 ;
        RECT 58.020 1686.380 61.020 1686.390 ;
        RECT 238.020 1686.380 241.020 1686.390 ;
        RECT 418.020 1686.380 421.020 1686.390 ;
        RECT 598.020 1686.380 601.020 1686.390 ;
        RECT 778.020 1686.380 781.020 1686.390 ;
        RECT 958.020 1686.380 961.020 1686.390 ;
        RECT 1138.020 1686.380 1141.020 1686.390 ;
        RECT 1318.020 1686.380 1321.020 1686.390 ;
        RECT 1498.020 1686.380 1501.020 1686.390 ;
        RECT 1678.020 1686.380 1681.020 1686.390 ;
        RECT 1858.020 1686.380 1861.020 1686.390 ;
        RECT 2038.020 1686.380 2041.020 1686.390 ;
        RECT 2218.020 1686.380 2221.020 1686.390 ;
        RECT 2398.020 1686.380 2401.020 1686.390 ;
        RECT 2578.020 1686.380 2581.020 1686.390 ;
        RECT 2758.020 1686.380 2761.020 1686.390 ;
        RECT 2954.200 1686.380 2957.200 1686.390 ;
        RECT -42.180 1683.380 2961.800 1686.380 ;
        RECT -37.580 1683.370 -34.580 1683.380 ;
        RECT 58.020 1683.370 61.020 1683.380 ;
        RECT 238.020 1683.370 241.020 1683.380 ;
        RECT 418.020 1683.370 421.020 1683.380 ;
        RECT 598.020 1683.370 601.020 1683.380 ;
        RECT 778.020 1683.370 781.020 1683.380 ;
        RECT 958.020 1683.370 961.020 1683.380 ;
        RECT 1138.020 1683.370 1141.020 1683.380 ;
        RECT 1318.020 1683.370 1321.020 1683.380 ;
        RECT 1498.020 1683.370 1501.020 1683.380 ;
        RECT 1678.020 1683.370 1681.020 1683.380 ;
        RECT 1858.020 1683.370 1861.020 1683.380 ;
        RECT 2038.020 1683.370 2041.020 1683.380 ;
        RECT 2218.020 1683.370 2221.020 1683.380 ;
        RECT 2398.020 1683.370 2401.020 1683.380 ;
        RECT 2578.020 1683.370 2581.020 1683.380 ;
        RECT 2758.020 1683.370 2761.020 1683.380 ;
        RECT 2954.200 1683.370 2957.200 1683.380 ;
        RECT -37.580 1506.380 -34.580 1506.390 ;
        RECT 58.020 1506.380 61.020 1506.390 ;
        RECT 238.020 1506.380 241.020 1506.390 ;
        RECT 418.020 1506.380 421.020 1506.390 ;
        RECT 598.020 1506.380 601.020 1506.390 ;
        RECT 778.020 1506.380 781.020 1506.390 ;
        RECT 958.020 1506.380 961.020 1506.390 ;
        RECT 1138.020 1506.380 1141.020 1506.390 ;
        RECT 1318.020 1506.380 1321.020 1506.390 ;
        RECT 1498.020 1506.380 1501.020 1506.390 ;
        RECT 1678.020 1506.380 1681.020 1506.390 ;
        RECT 1858.020 1506.380 1861.020 1506.390 ;
        RECT 2038.020 1506.380 2041.020 1506.390 ;
        RECT 2218.020 1506.380 2221.020 1506.390 ;
        RECT 2398.020 1506.380 2401.020 1506.390 ;
        RECT 2578.020 1506.380 2581.020 1506.390 ;
        RECT 2758.020 1506.380 2761.020 1506.390 ;
        RECT 2954.200 1506.380 2957.200 1506.390 ;
        RECT -42.180 1503.380 2961.800 1506.380 ;
        RECT -37.580 1503.370 -34.580 1503.380 ;
        RECT 58.020 1503.370 61.020 1503.380 ;
        RECT 238.020 1503.370 241.020 1503.380 ;
        RECT 418.020 1503.370 421.020 1503.380 ;
        RECT 598.020 1503.370 601.020 1503.380 ;
        RECT 778.020 1503.370 781.020 1503.380 ;
        RECT 958.020 1503.370 961.020 1503.380 ;
        RECT 1138.020 1503.370 1141.020 1503.380 ;
        RECT 1318.020 1503.370 1321.020 1503.380 ;
        RECT 1498.020 1503.370 1501.020 1503.380 ;
        RECT 1678.020 1503.370 1681.020 1503.380 ;
        RECT 1858.020 1503.370 1861.020 1503.380 ;
        RECT 2038.020 1503.370 2041.020 1503.380 ;
        RECT 2218.020 1503.370 2221.020 1503.380 ;
        RECT 2398.020 1503.370 2401.020 1503.380 ;
        RECT 2578.020 1503.370 2581.020 1503.380 ;
        RECT 2758.020 1503.370 2761.020 1503.380 ;
        RECT 2954.200 1503.370 2957.200 1503.380 ;
        RECT -37.580 1326.380 -34.580 1326.390 ;
        RECT 58.020 1326.380 61.020 1326.390 ;
        RECT 238.020 1326.380 241.020 1326.390 ;
        RECT 418.020 1326.380 421.020 1326.390 ;
        RECT 598.020 1326.380 601.020 1326.390 ;
        RECT 778.020 1326.380 781.020 1326.390 ;
        RECT 958.020 1326.380 961.020 1326.390 ;
        RECT 1138.020 1326.380 1141.020 1326.390 ;
        RECT 1318.020 1326.380 1321.020 1326.390 ;
        RECT 1498.020 1326.380 1501.020 1326.390 ;
        RECT 1678.020 1326.380 1681.020 1326.390 ;
        RECT 1858.020 1326.380 1861.020 1326.390 ;
        RECT 2038.020 1326.380 2041.020 1326.390 ;
        RECT 2218.020 1326.380 2221.020 1326.390 ;
        RECT 2398.020 1326.380 2401.020 1326.390 ;
        RECT 2578.020 1326.380 2581.020 1326.390 ;
        RECT 2758.020 1326.380 2761.020 1326.390 ;
        RECT 2954.200 1326.380 2957.200 1326.390 ;
        RECT -42.180 1323.380 2961.800 1326.380 ;
        RECT -37.580 1323.370 -34.580 1323.380 ;
        RECT 58.020 1323.370 61.020 1323.380 ;
        RECT 238.020 1323.370 241.020 1323.380 ;
        RECT 418.020 1323.370 421.020 1323.380 ;
        RECT 598.020 1323.370 601.020 1323.380 ;
        RECT 778.020 1323.370 781.020 1323.380 ;
        RECT 958.020 1323.370 961.020 1323.380 ;
        RECT 1138.020 1323.370 1141.020 1323.380 ;
        RECT 1318.020 1323.370 1321.020 1323.380 ;
        RECT 1498.020 1323.370 1501.020 1323.380 ;
        RECT 1678.020 1323.370 1681.020 1323.380 ;
        RECT 1858.020 1323.370 1861.020 1323.380 ;
        RECT 2038.020 1323.370 2041.020 1323.380 ;
        RECT 2218.020 1323.370 2221.020 1323.380 ;
        RECT 2398.020 1323.370 2401.020 1323.380 ;
        RECT 2578.020 1323.370 2581.020 1323.380 ;
        RECT 2758.020 1323.370 2761.020 1323.380 ;
        RECT 2954.200 1323.370 2957.200 1323.380 ;
        RECT -37.580 1146.380 -34.580 1146.390 ;
        RECT 58.020 1146.380 61.020 1146.390 ;
        RECT 238.020 1146.380 241.020 1146.390 ;
        RECT 418.020 1146.380 421.020 1146.390 ;
        RECT 598.020 1146.380 601.020 1146.390 ;
        RECT 778.020 1146.380 781.020 1146.390 ;
        RECT 958.020 1146.380 961.020 1146.390 ;
        RECT 1138.020 1146.380 1141.020 1146.390 ;
        RECT 1318.020 1146.380 1321.020 1146.390 ;
        RECT 1498.020 1146.380 1501.020 1146.390 ;
        RECT 1678.020 1146.380 1681.020 1146.390 ;
        RECT 1858.020 1146.380 1861.020 1146.390 ;
        RECT 2038.020 1146.380 2041.020 1146.390 ;
        RECT 2218.020 1146.380 2221.020 1146.390 ;
        RECT 2398.020 1146.380 2401.020 1146.390 ;
        RECT 2578.020 1146.380 2581.020 1146.390 ;
        RECT 2758.020 1146.380 2761.020 1146.390 ;
        RECT 2954.200 1146.380 2957.200 1146.390 ;
        RECT -42.180 1143.380 2961.800 1146.380 ;
        RECT -37.580 1143.370 -34.580 1143.380 ;
        RECT 58.020 1143.370 61.020 1143.380 ;
        RECT 238.020 1143.370 241.020 1143.380 ;
        RECT 418.020 1143.370 421.020 1143.380 ;
        RECT 598.020 1143.370 601.020 1143.380 ;
        RECT 778.020 1143.370 781.020 1143.380 ;
        RECT 958.020 1143.370 961.020 1143.380 ;
        RECT 1138.020 1143.370 1141.020 1143.380 ;
        RECT 1318.020 1143.370 1321.020 1143.380 ;
        RECT 1498.020 1143.370 1501.020 1143.380 ;
        RECT 1678.020 1143.370 1681.020 1143.380 ;
        RECT 1858.020 1143.370 1861.020 1143.380 ;
        RECT 2038.020 1143.370 2041.020 1143.380 ;
        RECT 2218.020 1143.370 2221.020 1143.380 ;
        RECT 2398.020 1143.370 2401.020 1143.380 ;
        RECT 2578.020 1143.370 2581.020 1143.380 ;
        RECT 2758.020 1143.370 2761.020 1143.380 ;
        RECT 2954.200 1143.370 2957.200 1143.380 ;
        RECT -37.580 966.380 -34.580 966.390 ;
        RECT 58.020 966.380 61.020 966.390 ;
        RECT 238.020 966.380 241.020 966.390 ;
        RECT 418.020 966.380 421.020 966.390 ;
        RECT 598.020 966.380 601.020 966.390 ;
        RECT 778.020 966.380 781.020 966.390 ;
        RECT 958.020 966.380 961.020 966.390 ;
        RECT 1138.020 966.380 1141.020 966.390 ;
        RECT 1318.020 966.380 1321.020 966.390 ;
        RECT 1498.020 966.380 1501.020 966.390 ;
        RECT 1678.020 966.380 1681.020 966.390 ;
        RECT 1858.020 966.380 1861.020 966.390 ;
        RECT 2038.020 966.380 2041.020 966.390 ;
        RECT 2218.020 966.380 2221.020 966.390 ;
        RECT 2398.020 966.380 2401.020 966.390 ;
        RECT 2578.020 966.380 2581.020 966.390 ;
        RECT 2758.020 966.380 2761.020 966.390 ;
        RECT 2954.200 966.380 2957.200 966.390 ;
        RECT -42.180 963.380 2961.800 966.380 ;
        RECT -37.580 963.370 -34.580 963.380 ;
        RECT 58.020 963.370 61.020 963.380 ;
        RECT 238.020 963.370 241.020 963.380 ;
        RECT 418.020 963.370 421.020 963.380 ;
        RECT 598.020 963.370 601.020 963.380 ;
        RECT 778.020 963.370 781.020 963.380 ;
        RECT 958.020 963.370 961.020 963.380 ;
        RECT 1138.020 963.370 1141.020 963.380 ;
        RECT 1318.020 963.370 1321.020 963.380 ;
        RECT 1498.020 963.370 1501.020 963.380 ;
        RECT 1678.020 963.370 1681.020 963.380 ;
        RECT 1858.020 963.370 1861.020 963.380 ;
        RECT 2038.020 963.370 2041.020 963.380 ;
        RECT 2218.020 963.370 2221.020 963.380 ;
        RECT 2398.020 963.370 2401.020 963.380 ;
        RECT 2578.020 963.370 2581.020 963.380 ;
        RECT 2758.020 963.370 2761.020 963.380 ;
        RECT 2954.200 963.370 2957.200 963.380 ;
        RECT -37.580 786.380 -34.580 786.390 ;
        RECT 58.020 786.380 61.020 786.390 ;
        RECT 238.020 786.380 241.020 786.390 ;
        RECT 418.020 786.380 421.020 786.390 ;
        RECT 598.020 786.380 601.020 786.390 ;
        RECT 778.020 786.380 781.020 786.390 ;
        RECT 958.020 786.380 961.020 786.390 ;
        RECT 1138.020 786.380 1141.020 786.390 ;
        RECT 1318.020 786.380 1321.020 786.390 ;
        RECT 1498.020 786.380 1501.020 786.390 ;
        RECT 1678.020 786.380 1681.020 786.390 ;
        RECT 1858.020 786.380 1861.020 786.390 ;
        RECT 2038.020 786.380 2041.020 786.390 ;
        RECT 2218.020 786.380 2221.020 786.390 ;
        RECT 2398.020 786.380 2401.020 786.390 ;
        RECT 2578.020 786.380 2581.020 786.390 ;
        RECT 2758.020 786.380 2761.020 786.390 ;
        RECT 2954.200 786.380 2957.200 786.390 ;
        RECT -42.180 783.380 2961.800 786.380 ;
        RECT -37.580 783.370 -34.580 783.380 ;
        RECT 58.020 783.370 61.020 783.380 ;
        RECT 238.020 783.370 241.020 783.380 ;
        RECT 418.020 783.370 421.020 783.380 ;
        RECT 598.020 783.370 601.020 783.380 ;
        RECT 778.020 783.370 781.020 783.380 ;
        RECT 958.020 783.370 961.020 783.380 ;
        RECT 1138.020 783.370 1141.020 783.380 ;
        RECT 1318.020 783.370 1321.020 783.380 ;
        RECT 1498.020 783.370 1501.020 783.380 ;
        RECT 1678.020 783.370 1681.020 783.380 ;
        RECT 1858.020 783.370 1861.020 783.380 ;
        RECT 2038.020 783.370 2041.020 783.380 ;
        RECT 2218.020 783.370 2221.020 783.380 ;
        RECT 2398.020 783.370 2401.020 783.380 ;
        RECT 2578.020 783.370 2581.020 783.380 ;
        RECT 2758.020 783.370 2761.020 783.380 ;
        RECT 2954.200 783.370 2957.200 783.380 ;
        RECT -37.580 606.380 -34.580 606.390 ;
        RECT 58.020 606.380 61.020 606.390 ;
        RECT 238.020 606.380 241.020 606.390 ;
        RECT 418.020 606.380 421.020 606.390 ;
        RECT 598.020 606.380 601.020 606.390 ;
        RECT 778.020 606.380 781.020 606.390 ;
        RECT 958.020 606.380 961.020 606.390 ;
        RECT 1138.020 606.380 1141.020 606.390 ;
        RECT 1318.020 606.380 1321.020 606.390 ;
        RECT 1498.020 606.380 1501.020 606.390 ;
        RECT 1678.020 606.380 1681.020 606.390 ;
        RECT 1858.020 606.380 1861.020 606.390 ;
        RECT 2038.020 606.380 2041.020 606.390 ;
        RECT 2218.020 606.380 2221.020 606.390 ;
        RECT 2398.020 606.380 2401.020 606.390 ;
        RECT 2578.020 606.380 2581.020 606.390 ;
        RECT 2758.020 606.380 2761.020 606.390 ;
        RECT 2954.200 606.380 2957.200 606.390 ;
        RECT -42.180 603.380 2961.800 606.380 ;
        RECT -37.580 603.370 -34.580 603.380 ;
        RECT 58.020 603.370 61.020 603.380 ;
        RECT 238.020 603.370 241.020 603.380 ;
        RECT 418.020 603.370 421.020 603.380 ;
        RECT 598.020 603.370 601.020 603.380 ;
        RECT 778.020 603.370 781.020 603.380 ;
        RECT 958.020 603.370 961.020 603.380 ;
        RECT 1138.020 603.370 1141.020 603.380 ;
        RECT 1318.020 603.370 1321.020 603.380 ;
        RECT 1498.020 603.370 1501.020 603.380 ;
        RECT 1678.020 603.370 1681.020 603.380 ;
        RECT 1858.020 603.370 1861.020 603.380 ;
        RECT 2038.020 603.370 2041.020 603.380 ;
        RECT 2218.020 603.370 2221.020 603.380 ;
        RECT 2398.020 603.370 2401.020 603.380 ;
        RECT 2578.020 603.370 2581.020 603.380 ;
        RECT 2758.020 603.370 2761.020 603.380 ;
        RECT 2954.200 603.370 2957.200 603.380 ;
        RECT -37.580 426.380 -34.580 426.390 ;
        RECT 58.020 426.380 61.020 426.390 ;
        RECT 238.020 426.380 241.020 426.390 ;
        RECT 418.020 426.380 421.020 426.390 ;
        RECT 598.020 426.380 601.020 426.390 ;
        RECT 778.020 426.380 781.020 426.390 ;
        RECT 958.020 426.380 961.020 426.390 ;
        RECT 1138.020 426.380 1141.020 426.390 ;
        RECT 1318.020 426.380 1321.020 426.390 ;
        RECT 1498.020 426.380 1501.020 426.390 ;
        RECT 1678.020 426.380 1681.020 426.390 ;
        RECT 1858.020 426.380 1861.020 426.390 ;
        RECT 2038.020 426.380 2041.020 426.390 ;
        RECT 2218.020 426.380 2221.020 426.390 ;
        RECT 2398.020 426.380 2401.020 426.390 ;
        RECT 2578.020 426.380 2581.020 426.390 ;
        RECT 2758.020 426.380 2761.020 426.390 ;
        RECT 2954.200 426.380 2957.200 426.390 ;
        RECT -42.180 423.380 2961.800 426.380 ;
        RECT -37.580 423.370 -34.580 423.380 ;
        RECT 58.020 423.370 61.020 423.380 ;
        RECT 238.020 423.370 241.020 423.380 ;
        RECT 418.020 423.370 421.020 423.380 ;
        RECT 598.020 423.370 601.020 423.380 ;
        RECT 778.020 423.370 781.020 423.380 ;
        RECT 958.020 423.370 961.020 423.380 ;
        RECT 1138.020 423.370 1141.020 423.380 ;
        RECT 1318.020 423.370 1321.020 423.380 ;
        RECT 1498.020 423.370 1501.020 423.380 ;
        RECT 1678.020 423.370 1681.020 423.380 ;
        RECT 1858.020 423.370 1861.020 423.380 ;
        RECT 2038.020 423.370 2041.020 423.380 ;
        RECT 2218.020 423.370 2221.020 423.380 ;
        RECT 2398.020 423.370 2401.020 423.380 ;
        RECT 2578.020 423.370 2581.020 423.380 ;
        RECT 2758.020 423.370 2761.020 423.380 ;
        RECT 2954.200 423.370 2957.200 423.380 ;
        RECT -37.580 246.380 -34.580 246.390 ;
        RECT 58.020 246.380 61.020 246.390 ;
        RECT 238.020 246.380 241.020 246.390 ;
        RECT 418.020 246.380 421.020 246.390 ;
        RECT 598.020 246.380 601.020 246.390 ;
        RECT 778.020 246.380 781.020 246.390 ;
        RECT 958.020 246.380 961.020 246.390 ;
        RECT 1138.020 246.380 1141.020 246.390 ;
        RECT 1318.020 246.380 1321.020 246.390 ;
        RECT 1498.020 246.380 1501.020 246.390 ;
        RECT 1678.020 246.380 1681.020 246.390 ;
        RECT 1858.020 246.380 1861.020 246.390 ;
        RECT 2038.020 246.380 2041.020 246.390 ;
        RECT 2218.020 246.380 2221.020 246.390 ;
        RECT 2398.020 246.380 2401.020 246.390 ;
        RECT 2578.020 246.380 2581.020 246.390 ;
        RECT 2758.020 246.380 2761.020 246.390 ;
        RECT 2954.200 246.380 2957.200 246.390 ;
        RECT -42.180 243.380 2961.800 246.380 ;
        RECT -37.580 243.370 -34.580 243.380 ;
        RECT 58.020 243.370 61.020 243.380 ;
        RECT 238.020 243.370 241.020 243.380 ;
        RECT 418.020 243.370 421.020 243.380 ;
        RECT 598.020 243.370 601.020 243.380 ;
        RECT 778.020 243.370 781.020 243.380 ;
        RECT 958.020 243.370 961.020 243.380 ;
        RECT 1138.020 243.370 1141.020 243.380 ;
        RECT 1318.020 243.370 1321.020 243.380 ;
        RECT 1498.020 243.370 1501.020 243.380 ;
        RECT 1678.020 243.370 1681.020 243.380 ;
        RECT 1858.020 243.370 1861.020 243.380 ;
        RECT 2038.020 243.370 2041.020 243.380 ;
        RECT 2218.020 243.370 2221.020 243.380 ;
        RECT 2398.020 243.370 2401.020 243.380 ;
        RECT 2578.020 243.370 2581.020 243.380 ;
        RECT 2758.020 243.370 2761.020 243.380 ;
        RECT 2954.200 243.370 2957.200 243.380 ;
        RECT -37.580 66.380 -34.580 66.390 ;
        RECT 58.020 66.380 61.020 66.390 ;
        RECT 238.020 66.380 241.020 66.390 ;
        RECT 418.020 66.380 421.020 66.390 ;
        RECT 598.020 66.380 601.020 66.390 ;
        RECT 778.020 66.380 781.020 66.390 ;
        RECT 958.020 66.380 961.020 66.390 ;
        RECT 1138.020 66.380 1141.020 66.390 ;
        RECT 1318.020 66.380 1321.020 66.390 ;
        RECT 1498.020 66.380 1501.020 66.390 ;
        RECT 1678.020 66.380 1681.020 66.390 ;
        RECT 1858.020 66.380 1861.020 66.390 ;
        RECT 2038.020 66.380 2041.020 66.390 ;
        RECT 2218.020 66.380 2221.020 66.390 ;
        RECT 2398.020 66.380 2401.020 66.390 ;
        RECT 2578.020 66.380 2581.020 66.390 ;
        RECT 2758.020 66.380 2761.020 66.390 ;
        RECT 2954.200 66.380 2957.200 66.390 ;
        RECT -42.180 63.380 2961.800 66.380 ;
        RECT -37.580 63.370 -34.580 63.380 ;
        RECT 58.020 63.370 61.020 63.380 ;
        RECT 238.020 63.370 241.020 63.380 ;
        RECT 418.020 63.370 421.020 63.380 ;
        RECT 598.020 63.370 601.020 63.380 ;
        RECT 778.020 63.370 781.020 63.380 ;
        RECT 958.020 63.370 961.020 63.380 ;
        RECT 1138.020 63.370 1141.020 63.380 ;
        RECT 1318.020 63.370 1321.020 63.380 ;
        RECT 1498.020 63.370 1501.020 63.380 ;
        RECT 1678.020 63.370 1681.020 63.380 ;
        RECT 1858.020 63.370 1861.020 63.380 ;
        RECT 2038.020 63.370 2041.020 63.380 ;
        RECT 2218.020 63.370 2221.020 63.380 ;
        RECT 2398.020 63.370 2401.020 63.380 ;
        RECT 2578.020 63.370 2581.020 63.380 ;
        RECT 2758.020 63.370 2761.020 63.380 ;
        RECT 2954.200 63.370 2957.200 63.380 ;
        RECT -37.580 -29.220 -34.580 -29.210 ;
        RECT 58.020 -29.220 61.020 -29.210 ;
        RECT 238.020 -29.220 241.020 -29.210 ;
        RECT 418.020 -29.220 421.020 -29.210 ;
        RECT 598.020 -29.220 601.020 -29.210 ;
        RECT 778.020 -29.220 781.020 -29.210 ;
        RECT 958.020 -29.220 961.020 -29.210 ;
        RECT 1138.020 -29.220 1141.020 -29.210 ;
        RECT 1318.020 -29.220 1321.020 -29.210 ;
        RECT 1498.020 -29.220 1501.020 -29.210 ;
        RECT 1678.020 -29.220 1681.020 -29.210 ;
        RECT 1858.020 -29.220 1861.020 -29.210 ;
        RECT 2038.020 -29.220 2041.020 -29.210 ;
        RECT 2218.020 -29.220 2221.020 -29.210 ;
        RECT 2398.020 -29.220 2401.020 -29.210 ;
        RECT 2578.020 -29.220 2581.020 -29.210 ;
        RECT 2758.020 -29.220 2761.020 -29.210 ;
        RECT 2954.200 -29.220 2957.200 -29.210 ;
        RECT -37.580 -32.220 2957.200 -29.220 ;
        RECT -37.580 -32.230 -34.580 -32.220 ;
        RECT 58.020 -32.230 61.020 -32.220 ;
        RECT 238.020 -32.230 241.020 -32.220 ;
        RECT 418.020 -32.230 421.020 -32.220 ;
        RECT 598.020 -32.230 601.020 -32.220 ;
        RECT 778.020 -32.230 781.020 -32.220 ;
        RECT 958.020 -32.230 961.020 -32.220 ;
        RECT 1138.020 -32.230 1141.020 -32.220 ;
        RECT 1318.020 -32.230 1321.020 -32.220 ;
        RECT 1498.020 -32.230 1501.020 -32.220 ;
        RECT 1678.020 -32.230 1681.020 -32.220 ;
        RECT 1858.020 -32.230 1861.020 -32.220 ;
        RECT 2038.020 -32.230 2041.020 -32.220 ;
        RECT 2218.020 -32.230 2221.020 -32.220 ;
        RECT 2398.020 -32.230 2401.020 -32.220 ;
        RECT 2578.020 -32.230 2581.020 -32.220 ;
        RECT 2758.020 -32.230 2761.020 -32.220 ;
        RECT 2954.200 -32.230 2957.200 -32.220 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -42.180 -36.820 -39.180 3556.500 ;
        RECT 148.020 -36.820 151.020 3556.500 ;
        RECT 328.020 -36.820 331.020 3556.500 ;
        RECT 508.020 -36.820 511.020 3556.500 ;
        RECT 688.020 -36.820 691.020 3556.500 ;
        RECT 868.020 -36.820 871.020 3556.500 ;
        RECT 1048.020 -36.820 1051.020 3556.500 ;
        RECT 1228.020 -36.820 1231.020 3556.500 ;
        RECT 1408.020 -36.820 1411.020 3556.500 ;
        RECT 1588.020 -36.820 1591.020 3556.500 ;
        RECT 1768.020 -36.820 1771.020 3556.500 ;
        RECT 1948.020 -36.820 1951.020 3556.500 ;
        RECT 2128.020 -36.820 2131.020 3556.500 ;
        RECT 2308.020 -36.820 2311.020 3556.500 ;
        RECT 2488.020 -36.820 2491.020 3556.500 ;
        RECT 2668.020 -36.820 2671.020 3556.500 ;
        RECT 2848.020 -36.820 2851.020 3556.500 ;
        RECT 2958.800 -36.820 2961.800 3556.500 ;
      LAYER via4 ;
        RECT -41.270 3555.210 -40.090 3556.390 ;
        RECT -41.270 3553.610 -40.090 3554.790 ;
        RECT -41.270 3395.090 -40.090 3396.270 ;
        RECT -41.270 3393.490 -40.090 3394.670 ;
        RECT -41.270 3215.090 -40.090 3216.270 ;
        RECT -41.270 3213.490 -40.090 3214.670 ;
        RECT -41.270 3035.090 -40.090 3036.270 ;
        RECT -41.270 3033.490 -40.090 3034.670 ;
        RECT -41.270 2855.090 -40.090 2856.270 ;
        RECT -41.270 2853.490 -40.090 2854.670 ;
        RECT -41.270 2675.090 -40.090 2676.270 ;
        RECT -41.270 2673.490 -40.090 2674.670 ;
        RECT -41.270 2495.090 -40.090 2496.270 ;
        RECT -41.270 2493.490 -40.090 2494.670 ;
        RECT -41.270 2315.090 -40.090 2316.270 ;
        RECT -41.270 2313.490 -40.090 2314.670 ;
        RECT -41.270 2135.090 -40.090 2136.270 ;
        RECT -41.270 2133.490 -40.090 2134.670 ;
        RECT -41.270 1955.090 -40.090 1956.270 ;
        RECT -41.270 1953.490 -40.090 1954.670 ;
        RECT -41.270 1775.090 -40.090 1776.270 ;
        RECT -41.270 1773.490 -40.090 1774.670 ;
        RECT -41.270 1595.090 -40.090 1596.270 ;
        RECT -41.270 1593.490 -40.090 1594.670 ;
        RECT -41.270 1415.090 -40.090 1416.270 ;
        RECT -41.270 1413.490 -40.090 1414.670 ;
        RECT -41.270 1235.090 -40.090 1236.270 ;
        RECT -41.270 1233.490 -40.090 1234.670 ;
        RECT -41.270 1055.090 -40.090 1056.270 ;
        RECT -41.270 1053.490 -40.090 1054.670 ;
        RECT -41.270 875.090 -40.090 876.270 ;
        RECT -41.270 873.490 -40.090 874.670 ;
        RECT -41.270 695.090 -40.090 696.270 ;
        RECT -41.270 693.490 -40.090 694.670 ;
        RECT -41.270 515.090 -40.090 516.270 ;
        RECT -41.270 513.490 -40.090 514.670 ;
        RECT -41.270 335.090 -40.090 336.270 ;
        RECT -41.270 333.490 -40.090 334.670 ;
        RECT -41.270 155.090 -40.090 156.270 ;
        RECT -41.270 153.490 -40.090 154.670 ;
        RECT -41.270 -35.110 -40.090 -33.930 ;
        RECT -41.270 -36.710 -40.090 -35.530 ;
        RECT 148.930 3555.210 150.110 3556.390 ;
        RECT 148.930 3553.610 150.110 3554.790 ;
        RECT 148.930 3395.090 150.110 3396.270 ;
        RECT 148.930 3393.490 150.110 3394.670 ;
        RECT 148.930 3215.090 150.110 3216.270 ;
        RECT 148.930 3213.490 150.110 3214.670 ;
        RECT 148.930 3035.090 150.110 3036.270 ;
        RECT 148.930 3033.490 150.110 3034.670 ;
        RECT 148.930 2855.090 150.110 2856.270 ;
        RECT 148.930 2853.490 150.110 2854.670 ;
        RECT 148.930 2675.090 150.110 2676.270 ;
        RECT 148.930 2673.490 150.110 2674.670 ;
        RECT 148.930 2495.090 150.110 2496.270 ;
        RECT 148.930 2493.490 150.110 2494.670 ;
        RECT 148.930 2315.090 150.110 2316.270 ;
        RECT 148.930 2313.490 150.110 2314.670 ;
        RECT 148.930 2135.090 150.110 2136.270 ;
        RECT 148.930 2133.490 150.110 2134.670 ;
        RECT 148.930 1955.090 150.110 1956.270 ;
        RECT 148.930 1953.490 150.110 1954.670 ;
        RECT 148.930 1775.090 150.110 1776.270 ;
        RECT 148.930 1773.490 150.110 1774.670 ;
        RECT 148.930 1595.090 150.110 1596.270 ;
        RECT 148.930 1593.490 150.110 1594.670 ;
        RECT 148.930 1415.090 150.110 1416.270 ;
        RECT 148.930 1413.490 150.110 1414.670 ;
        RECT 148.930 1235.090 150.110 1236.270 ;
        RECT 148.930 1233.490 150.110 1234.670 ;
        RECT 148.930 1055.090 150.110 1056.270 ;
        RECT 148.930 1053.490 150.110 1054.670 ;
        RECT 148.930 875.090 150.110 876.270 ;
        RECT 148.930 873.490 150.110 874.670 ;
        RECT 148.930 695.090 150.110 696.270 ;
        RECT 148.930 693.490 150.110 694.670 ;
        RECT 148.930 515.090 150.110 516.270 ;
        RECT 148.930 513.490 150.110 514.670 ;
        RECT 148.930 335.090 150.110 336.270 ;
        RECT 148.930 333.490 150.110 334.670 ;
        RECT 148.930 155.090 150.110 156.270 ;
        RECT 148.930 153.490 150.110 154.670 ;
        RECT 148.930 -35.110 150.110 -33.930 ;
        RECT 148.930 -36.710 150.110 -35.530 ;
        RECT 328.930 3555.210 330.110 3556.390 ;
        RECT 328.930 3553.610 330.110 3554.790 ;
        RECT 328.930 3395.090 330.110 3396.270 ;
        RECT 328.930 3393.490 330.110 3394.670 ;
        RECT 328.930 3215.090 330.110 3216.270 ;
        RECT 328.930 3213.490 330.110 3214.670 ;
        RECT 328.930 3035.090 330.110 3036.270 ;
        RECT 328.930 3033.490 330.110 3034.670 ;
        RECT 328.930 2855.090 330.110 2856.270 ;
        RECT 328.930 2853.490 330.110 2854.670 ;
        RECT 328.930 2675.090 330.110 2676.270 ;
        RECT 328.930 2673.490 330.110 2674.670 ;
        RECT 328.930 2495.090 330.110 2496.270 ;
        RECT 328.930 2493.490 330.110 2494.670 ;
        RECT 328.930 2315.090 330.110 2316.270 ;
        RECT 328.930 2313.490 330.110 2314.670 ;
        RECT 328.930 2135.090 330.110 2136.270 ;
        RECT 328.930 2133.490 330.110 2134.670 ;
        RECT 328.930 1955.090 330.110 1956.270 ;
        RECT 328.930 1953.490 330.110 1954.670 ;
        RECT 328.930 1775.090 330.110 1776.270 ;
        RECT 328.930 1773.490 330.110 1774.670 ;
        RECT 328.930 1595.090 330.110 1596.270 ;
        RECT 328.930 1593.490 330.110 1594.670 ;
        RECT 328.930 1415.090 330.110 1416.270 ;
        RECT 328.930 1413.490 330.110 1414.670 ;
        RECT 328.930 1235.090 330.110 1236.270 ;
        RECT 328.930 1233.490 330.110 1234.670 ;
        RECT 328.930 1055.090 330.110 1056.270 ;
        RECT 328.930 1053.490 330.110 1054.670 ;
        RECT 328.930 875.090 330.110 876.270 ;
        RECT 328.930 873.490 330.110 874.670 ;
        RECT 328.930 695.090 330.110 696.270 ;
        RECT 328.930 693.490 330.110 694.670 ;
        RECT 328.930 515.090 330.110 516.270 ;
        RECT 328.930 513.490 330.110 514.670 ;
        RECT 328.930 335.090 330.110 336.270 ;
        RECT 328.930 333.490 330.110 334.670 ;
        RECT 328.930 155.090 330.110 156.270 ;
        RECT 328.930 153.490 330.110 154.670 ;
        RECT 328.930 -35.110 330.110 -33.930 ;
        RECT 328.930 -36.710 330.110 -35.530 ;
        RECT 508.930 3555.210 510.110 3556.390 ;
        RECT 508.930 3553.610 510.110 3554.790 ;
        RECT 508.930 3395.090 510.110 3396.270 ;
        RECT 508.930 3393.490 510.110 3394.670 ;
        RECT 508.930 3215.090 510.110 3216.270 ;
        RECT 508.930 3213.490 510.110 3214.670 ;
        RECT 508.930 3035.090 510.110 3036.270 ;
        RECT 508.930 3033.490 510.110 3034.670 ;
        RECT 508.930 2855.090 510.110 2856.270 ;
        RECT 508.930 2853.490 510.110 2854.670 ;
        RECT 508.930 2675.090 510.110 2676.270 ;
        RECT 508.930 2673.490 510.110 2674.670 ;
        RECT 508.930 2495.090 510.110 2496.270 ;
        RECT 508.930 2493.490 510.110 2494.670 ;
        RECT 508.930 2315.090 510.110 2316.270 ;
        RECT 508.930 2313.490 510.110 2314.670 ;
        RECT 508.930 2135.090 510.110 2136.270 ;
        RECT 508.930 2133.490 510.110 2134.670 ;
        RECT 508.930 1955.090 510.110 1956.270 ;
        RECT 508.930 1953.490 510.110 1954.670 ;
        RECT 508.930 1775.090 510.110 1776.270 ;
        RECT 508.930 1773.490 510.110 1774.670 ;
        RECT 508.930 1595.090 510.110 1596.270 ;
        RECT 508.930 1593.490 510.110 1594.670 ;
        RECT 508.930 1415.090 510.110 1416.270 ;
        RECT 508.930 1413.490 510.110 1414.670 ;
        RECT 508.930 1235.090 510.110 1236.270 ;
        RECT 508.930 1233.490 510.110 1234.670 ;
        RECT 508.930 1055.090 510.110 1056.270 ;
        RECT 508.930 1053.490 510.110 1054.670 ;
        RECT 508.930 875.090 510.110 876.270 ;
        RECT 508.930 873.490 510.110 874.670 ;
        RECT 508.930 695.090 510.110 696.270 ;
        RECT 508.930 693.490 510.110 694.670 ;
        RECT 508.930 515.090 510.110 516.270 ;
        RECT 508.930 513.490 510.110 514.670 ;
        RECT 508.930 335.090 510.110 336.270 ;
        RECT 508.930 333.490 510.110 334.670 ;
        RECT 508.930 155.090 510.110 156.270 ;
        RECT 508.930 153.490 510.110 154.670 ;
        RECT 508.930 -35.110 510.110 -33.930 ;
        RECT 508.930 -36.710 510.110 -35.530 ;
        RECT 688.930 3555.210 690.110 3556.390 ;
        RECT 688.930 3553.610 690.110 3554.790 ;
        RECT 688.930 3395.090 690.110 3396.270 ;
        RECT 688.930 3393.490 690.110 3394.670 ;
        RECT 688.930 3215.090 690.110 3216.270 ;
        RECT 688.930 3213.490 690.110 3214.670 ;
        RECT 688.930 3035.090 690.110 3036.270 ;
        RECT 688.930 3033.490 690.110 3034.670 ;
        RECT 688.930 2855.090 690.110 2856.270 ;
        RECT 688.930 2853.490 690.110 2854.670 ;
        RECT 688.930 2675.090 690.110 2676.270 ;
        RECT 688.930 2673.490 690.110 2674.670 ;
        RECT 688.930 2495.090 690.110 2496.270 ;
        RECT 688.930 2493.490 690.110 2494.670 ;
        RECT 688.930 2315.090 690.110 2316.270 ;
        RECT 688.930 2313.490 690.110 2314.670 ;
        RECT 688.930 2135.090 690.110 2136.270 ;
        RECT 688.930 2133.490 690.110 2134.670 ;
        RECT 688.930 1955.090 690.110 1956.270 ;
        RECT 688.930 1953.490 690.110 1954.670 ;
        RECT 688.930 1775.090 690.110 1776.270 ;
        RECT 688.930 1773.490 690.110 1774.670 ;
        RECT 688.930 1595.090 690.110 1596.270 ;
        RECT 688.930 1593.490 690.110 1594.670 ;
        RECT 688.930 1415.090 690.110 1416.270 ;
        RECT 688.930 1413.490 690.110 1414.670 ;
        RECT 688.930 1235.090 690.110 1236.270 ;
        RECT 688.930 1233.490 690.110 1234.670 ;
        RECT 688.930 1055.090 690.110 1056.270 ;
        RECT 688.930 1053.490 690.110 1054.670 ;
        RECT 688.930 875.090 690.110 876.270 ;
        RECT 688.930 873.490 690.110 874.670 ;
        RECT 688.930 695.090 690.110 696.270 ;
        RECT 688.930 693.490 690.110 694.670 ;
        RECT 688.930 515.090 690.110 516.270 ;
        RECT 688.930 513.490 690.110 514.670 ;
        RECT 688.930 335.090 690.110 336.270 ;
        RECT 688.930 333.490 690.110 334.670 ;
        RECT 688.930 155.090 690.110 156.270 ;
        RECT 688.930 153.490 690.110 154.670 ;
        RECT 688.930 -35.110 690.110 -33.930 ;
        RECT 688.930 -36.710 690.110 -35.530 ;
        RECT 868.930 3555.210 870.110 3556.390 ;
        RECT 868.930 3553.610 870.110 3554.790 ;
        RECT 868.930 3395.090 870.110 3396.270 ;
        RECT 868.930 3393.490 870.110 3394.670 ;
        RECT 868.930 3215.090 870.110 3216.270 ;
        RECT 868.930 3213.490 870.110 3214.670 ;
        RECT 868.930 3035.090 870.110 3036.270 ;
        RECT 868.930 3033.490 870.110 3034.670 ;
        RECT 868.930 2855.090 870.110 2856.270 ;
        RECT 868.930 2853.490 870.110 2854.670 ;
        RECT 868.930 2675.090 870.110 2676.270 ;
        RECT 868.930 2673.490 870.110 2674.670 ;
        RECT 868.930 2495.090 870.110 2496.270 ;
        RECT 868.930 2493.490 870.110 2494.670 ;
        RECT 868.930 2315.090 870.110 2316.270 ;
        RECT 868.930 2313.490 870.110 2314.670 ;
        RECT 868.930 2135.090 870.110 2136.270 ;
        RECT 868.930 2133.490 870.110 2134.670 ;
        RECT 868.930 1955.090 870.110 1956.270 ;
        RECT 868.930 1953.490 870.110 1954.670 ;
        RECT 868.930 1775.090 870.110 1776.270 ;
        RECT 868.930 1773.490 870.110 1774.670 ;
        RECT 868.930 1595.090 870.110 1596.270 ;
        RECT 868.930 1593.490 870.110 1594.670 ;
        RECT 868.930 1415.090 870.110 1416.270 ;
        RECT 868.930 1413.490 870.110 1414.670 ;
        RECT 868.930 1235.090 870.110 1236.270 ;
        RECT 868.930 1233.490 870.110 1234.670 ;
        RECT 868.930 1055.090 870.110 1056.270 ;
        RECT 868.930 1053.490 870.110 1054.670 ;
        RECT 868.930 875.090 870.110 876.270 ;
        RECT 868.930 873.490 870.110 874.670 ;
        RECT 868.930 695.090 870.110 696.270 ;
        RECT 868.930 693.490 870.110 694.670 ;
        RECT 868.930 515.090 870.110 516.270 ;
        RECT 868.930 513.490 870.110 514.670 ;
        RECT 868.930 335.090 870.110 336.270 ;
        RECT 868.930 333.490 870.110 334.670 ;
        RECT 868.930 155.090 870.110 156.270 ;
        RECT 868.930 153.490 870.110 154.670 ;
        RECT 868.930 -35.110 870.110 -33.930 ;
        RECT 868.930 -36.710 870.110 -35.530 ;
        RECT 1048.930 3555.210 1050.110 3556.390 ;
        RECT 1048.930 3553.610 1050.110 3554.790 ;
        RECT 1048.930 3395.090 1050.110 3396.270 ;
        RECT 1048.930 3393.490 1050.110 3394.670 ;
        RECT 1048.930 3215.090 1050.110 3216.270 ;
        RECT 1048.930 3213.490 1050.110 3214.670 ;
        RECT 1048.930 3035.090 1050.110 3036.270 ;
        RECT 1048.930 3033.490 1050.110 3034.670 ;
        RECT 1048.930 2855.090 1050.110 2856.270 ;
        RECT 1048.930 2853.490 1050.110 2854.670 ;
        RECT 1048.930 2675.090 1050.110 2676.270 ;
        RECT 1048.930 2673.490 1050.110 2674.670 ;
        RECT 1048.930 2495.090 1050.110 2496.270 ;
        RECT 1048.930 2493.490 1050.110 2494.670 ;
        RECT 1048.930 2315.090 1050.110 2316.270 ;
        RECT 1048.930 2313.490 1050.110 2314.670 ;
        RECT 1048.930 2135.090 1050.110 2136.270 ;
        RECT 1048.930 2133.490 1050.110 2134.670 ;
        RECT 1048.930 1955.090 1050.110 1956.270 ;
        RECT 1048.930 1953.490 1050.110 1954.670 ;
        RECT 1048.930 1775.090 1050.110 1776.270 ;
        RECT 1048.930 1773.490 1050.110 1774.670 ;
        RECT 1048.930 1595.090 1050.110 1596.270 ;
        RECT 1048.930 1593.490 1050.110 1594.670 ;
        RECT 1048.930 1415.090 1050.110 1416.270 ;
        RECT 1048.930 1413.490 1050.110 1414.670 ;
        RECT 1048.930 1235.090 1050.110 1236.270 ;
        RECT 1048.930 1233.490 1050.110 1234.670 ;
        RECT 1048.930 1055.090 1050.110 1056.270 ;
        RECT 1048.930 1053.490 1050.110 1054.670 ;
        RECT 1048.930 875.090 1050.110 876.270 ;
        RECT 1048.930 873.490 1050.110 874.670 ;
        RECT 1048.930 695.090 1050.110 696.270 ;
        RECT 1048.930 693.490 1050.110 694.670 ;
        RECT 1048.930 515.090 1050.110 516.270 ;
        RECT 1048.930 513.490 1050.110 514.670 ;
        RECT 1048.930 335.090 1050.110 336.270 ;
        RECT 1048.930 333.490 1050.110 334.670 ;
        RECT 1048.930 155.090 1050.110 156.270 ;
        RECT 1048.930 153.490 1050.110 154.670 ;
        RECT 1048.930 -35.110 1050.110 -33.930 ;
        RECT 1048.930 -36.710 1050.110 -35.530 ;
        RECT 1228.930 3555.210 1230.110 3556.390 ;
        RECT 1228.930 3553.610 1230.110 3554.790 ;
        RECT 1228.930 3395.090 1230.110 3396.270 ;
        RECT 1228.930 3393.490 1230.110 3394.670 ;
        RECT 1228.930 3215.090 1230.110 3216.270 ;
        RECT 1228.930 3213.490 1230.110 3214.670 ;
        RECT 1228.930 3035.090 1230.110 3036.270 ;
        RECT 1228.930 3033.490 1230.110 3034.670 ;
        RECT 1228.930 2855.090 1230.110 2856.270 ;
        RECT 1228.930 2853.490 1230.110 2854.670 ;
        RECT 1228.930 2675.090 1230.110 2676.270 ;
        RECT 1228.930 2673.490 1230.110 2674.670 ;
        RECT 1228.930 2495.090 1230.110 2496.270 ;
        RECT 1228.930 2493.490 1230.110 2494.670 ;
        RECT 1228.930 2315.090 1230.110 2316.270 ;
        RECT 1228.930 2313.490 1230.110 2314.670 ;
        RECT 1228.930 2135.090 1230.110 2136.270 ;
        RECT 1228.930 2133.490 1230.110 2134.670 ;
        RECT 1228.930 1955.090 1230.110 1956.270 ;
        RECT 1228.930 1953.490 1230.110 1954.670 ;
        RECT 1228.930 1775.090 1230.110 1776.270 ;
        RECT 1228.930 1773.490 1230.110 1774.670 ;
        RECT 1228.930 1595.090 1230.110 1596.270 ;
        RECT 1228.930 1593.490 1230.110 1594.670 ;
        RECT 1228.930 1415.090 1230.110 1416.270 ;
        RECT 1228.930 1413.490 1230.110 1414.670 ;
        RECT 1228.930 1235.090 1230.110 1236.270 ;
        RECT 1228.930 1233.490 1230.110 1234.670 ;
        RECT 1228.930 1055.090 1230.110 1056.270 ;
        RECT 1228.930 1053.490 1230.110 1054.670 ;
        RECT 1228.930 875.090 1230.110 876.270 ;
        RECT 1228.930 873.490 1230.110 874.670 ;
        RECT 1228.930 695.090 1230.110 696.270 ;
        RECT 1228.930 693.490 1230.110 694.670 ;
        RECT 1228.930 515.090 1230.110 516.270 ;
        RECT 1228.930 513.490 1230.110 514.670 ;
        RECT 1228.930 335.090 1230.110 336.270 ;
        RECT 1228.930 333.490 1230.110 334.670 ;
        RECT 1228.930 155.090 1230.110 156.270 ;
        RECT 1228.930 153.490 1230.110 154.670 ;
        RECT 1228.930 -35.110 1230.110 -33.930 ;
        RECT 1228.930 -36.710 1230.110 -35.530 ;
        RECT 1408.930 3555.210 1410.110 3556.390 ;
        RECT 1408.930 3553.610 1410.110 3554.790 ;
        RECT 1408.930 3395.090 1410.110 3396.270 ;
        RECT 1408.930 3393.490 1410.110 3394.670 ;
        RECT 1408.930 3215.090 1410.110 3216.270 ;
        RECT 1408.930 3213.490 1410.110 3214.670 ;
        RECT 1408.930 3035.090 1410.110 3036.270 ;
        RECT 1408.930 3033.490 1410.110 3034.670 ;
        RECT 1408.930 2855.090 1410.110 2856.270 ;
        RECT 1408.930 2853.490 1410.110 2854.670 ;
        RECT 1408.930 2675.090 1410.110 2676.270 ;
        RECT 1408.930 2673.490 1410.110 2674.670 ;
        RECT 1408.930 2495.090 1410.110 2496.270 ;
        RECT 1408.930 2493.490 1410.110 2494.670 ;
        RECT 1408.930 2315.090 1410.110 2316.270 ;
        RECT 1408.930 2313.490 1410.110 2314.670 ;
        RECT 1408.930 2135.090 1410.110 2136.270 ;
        RECT 1408.930 2133.490 1410.110 2134.670 ;
        RECT 1408.930 1955.090 1410.110 1956.270 ;
        RECT 1408.930 1953.490 1410.110 1954.670 ;
        RECT 1408.930 1775.090 1410.110 1776.270 ;
        RECT 1408.930 1773.490 1410.110 1774.670 ;
        RECT 1408.930 1595.090 1410.110 1596.270 ;
        RECT 1408.930 1593.490 1410.110 1594.670 ;
        RECT 1408.930 1415.090 1410.110 1416.270 ;
        RECT 1408.930 1413.490 1410.110 1414.670 ;
        RECT 1408.930 1235.090 1410.110 1236.270 ;
        RECT 1408.930 1233.490 1410.110 1234.670 ;
        RECT 1408.930 1055.090 1410.110 1056.270 ;
        RECT 1408.930 1053.490 1410.110 1054.670 ;
        RECT 1408.930 875.090 1410.110 876.270 ;
        RECT 1408.930 873.490 1410.110 874.670 ;
        RECT 1408.930 695.090 1410.110 696.270 ;
        RECT 1408.930 693.490 1410.110 694.670 ;
        RECT 1408.930 515.090 1410.110 516.270 ;
        RECT 1408.930 513.490 1410.110 514.670 ;
        RECT 1408.930 335.090 1410.110 336.270 ;
        RECT 1408.930 333.490 1410.110 334.670 ;
        RECT 1408.930 155.090 1410.110 156.270 ;
        RECT 1408.930 153.490 1410.110 154.670 ;
        RECT 1408.930 -35.110 1410.110 -33.930 ;
        RECT 1408.930 -36.710 1410.110 -35.530 ;
        RECT 1588.930 3555.210 1590.110 3556.390 ;
        RECT 1588.930 3553.610 1590.110 3554.790 ;
        RECT 1588.930 3395.090 1590.110 3396.270 ;
        RECT 1588.930 3393.490 1590.110 3394.670 ;
        RECT 1588.930 3215.090 1590.110 3216.270 ;
        RECT 1588.930 3213.490 1590.110 3214.670 ;
        RECT 1588.930 3035.090 1590.110 3036.270 ;
        RECT 1588.930 3033.490 1590.110 3034.670 ;
        RECT 1588.930 2855.090 1590.110 2856.270 ;
        RECT 1588.930 2853.490 1590.110 2854.670 ;
        RECT 1588.930 2675.090 1590.110 2676.270 ;
        RECT 1588.930 2673.490 1590.110 2674.670 ;
        RECT 1588.930 2495.090 1590.110 2496.270 ;
        RECT 1588.930 2493.490 1590.110 2494.670 ;
        RECT 1588.930 2315.090 1590.110 2316.270 ;
        RECT 1588.930 2313.490 1590.110 2314.670 ;
        RECT 1588.930 2135.090 1590.110 2136.270 ;
        RECT 1588.930 2133.490 1590.110 2134.670 ;
        RECT 1588.930 1955.090 1590.110 1956.270 ;
        RECT 1588.930 1953.490 1590.110 1954.670 ;
        RECT 1588.930 1775.090 1590.110 1776.270 ;
        RECT 1588.930 1773.490 1590.110 1774.670 ;
        RECT 1588.930 1595.090 1590.110 1596.270 ;
        RECT 1588.930 1593.490 1590.110 1594.670 ;
        RECT 1588.930 1415.090 1590.110 1416.270 ;
        RECT 1588.930 1413.490 1590.110 1414.670 ;
        RECT 1588.930 1235.090 1590.110 1236.270 ;
        RECT 1588.930 1233.490 1590.110 1234.670 ;
        RECT 1588.930 1055.090 1590.110 1056.270 ;
        RECT 1588.930 1053.490 1590.110 1054.670 ;
        RECT 1588.930 875.090 1590.110 876.270 ;
        RECT 1588.930 873.490 1590.110 874.670 ;
        RECT 1588.930 695.090 1590.110 696.270 ;
        RECT 1588.930 693.490 1590.110 694.670 ;
        RECT 1588.930 515.090 1590.110 516.270 ;
        RECT 1588.930 513.490 1590.110 514.670 ;
        RECT 1588.930 335.090 1590.110 336.270 ;
        RECT 1588.930 333.490 1590.110 334.670 ;
        RECT 1588.930 155.090 1590.110 156.270 ;
        RECT 1588.930 153.490 1590.110 154.670 ;
        RECT 1588.930 -35.110 1590.110 -33.930 ;
        RECT 1588.930 -36.710 1590.110 -35.530 ;
        RECT 1768.930 3555.210 1770.110 3556.390 ;
        RECT 1768.930 3553.610 1770.110 3554.790 ;
        RECT 1768.930 3395.090 1770.110 3396.270 ;
        RECT 1768.930 3393.490 1770.110 3394.670 ;
        RECT 1768.930 3215.090 1770.110 3216.270 ;
        RECT 1768.930 3213.490 1770.110 3214.670 ;
        RECT 1768.930 3035.090 1770.110 3036.270 ;
        RECT 1768.930 3033.490 1770.110 3034.670 ;
        RECT 1768.930 2855.090 1770.110 2856.270 ;
        RECT 1768.930 2853.490 1770.110 2854.670 ;
        RECT 1768.930 2675.090 1770.110 2676.270 ;
        RECT 1768.930 2673.490 1770.110 2674.670 ;
        RECT 1768.930 2495.090 1770.110 2496.270 ;
        RECT 1768.930 2493.490 1770.110 2494.670 ;
        RECT 1768.930 2315.090 1770.110 2316.270 ;
        RECT 1768.930 2313.490 1770.110 2314.670 ;
        RECT 1768.930 2135.090 1770.110 2136.270 ;
        RECT 1768.930 2133.490 1770.110 2134.670 ;
        RECT 1768.930 1955.090 1770.110 1956.270 ;
        RECT 1768.930 1953.490 1770.110 1954.670 ;
        RECT 1768.930 1775.090 1770.110 1776.270 ;
        RECT 1768.930 1773.490 1770.110 1774.670 ;
        RECT 1768.930 1595.090 1770.110 1596.270 ;
        RECT 1768.930 1593.490 1770.110 1594.670 ;
        RECT 1768.930 1415.090 1770.110 1416.270 ;
        RECT 1768.930 1413.490 1770.110 1414.670 ;
        RECT 1768.930 1235.090 1770.110 1236.270 ;
        RECT 1768.930 1233.490 1770.110 1234.670 ;
        RECT 1768.930 1055.090 1770.110 1056.270 ;
        RECT 1768.930 1053.490 1770.110 1054.670 ;
        RECT 1768.930 875.090 1770.110 876.270 ;
        RECT 1768.930 873.490 1770.110 874.670 ;
        RECT 1768.930 695.090 1770.110 696.270 ;
        RECT 1768.930 693.490 1770.110 694.670 ;
        RECT 1768.930 515.090 1770.110 516.270 ;
        RECT 1768.930 513.490 1770.110 514.670 ;
        RECT 1768.930 335.090 1770.110 336.270 ;
        RECT 1768.930 333.490 1770.110 334.670 ;
        RECT 1768.930 155.090 1770.110 156.270 ;
        RECT 1768.930 153.490 1770.110 154.670 ;
        RECT 1768.930 -35.110 1770.110 -33.930 ;
        RECT 1768.930 -36.710 1770.110 -35.530 ;
        RECT 1948.930 3555.210 1950.110 3556.390 ;
        RECT 1948.930 3553.610 1950.110 3554.790 ;
        RECT 1948.930 3395.090 1950.110 3396.270 ;
        RECT 1948.930 3393.490 1950.110 3394.670 ;
        RECT 1948.930 3215.090 1950.110 3216.270 ;
        RECT 1948.930 3213.490 1950.110 3214.670 ;
        RECT 1948.930 3035.090 1950.110 3036.270 ;
        RECT 1948.930 3033.490 1950.110 3034.670 ;
        RECT 1948.930 2855.090 1950.110 2856.270 ;
        RECT 1948.930 2853.490 1950.110 2854.670 ;
        RECT 1948.930 2675.090 1950.110 2676.270 ;
        RECT 1948.930 2673.490 1950.110 2674.670 ;
        RECT 1948.930 2495.090 1950.110 2496.270 ;
        RECT 1948.930 2493.490 1950.110 2494.670 ;
        RECT 1948.930 2315.090 1950.110 2316.270 ;
        RECT 1948.930 2313.490 1950.110 2314.670 ;
        RECT 1948.930 2135.090 1950.110 2136.270 ;
        RECT 1948.930 2133.490 1950.110 2134.670 ;
        RECT 1948.930 1955.090 1950.110 1956.270 ;
        RECT 1948.930 1953.490 1950.110 1954.670 ;
        RECT 1948.930 1775.090 1950.110 1776.270 ;
        RECT 1948.930 1773.490 1950.110 1774.670 ;
        RECT 1948.930 1595.090 1950.110 1596.270 ;
        RECT 1948.930 1593.490 1950.110 1594.670 ;
        RECT 1948.930 1415.090 1950.110 1416.270 ;
        RECT 1948.930 1413.490 1950.110 1414.670 ;
        RECT 1948.930 1235.090 1950.110 1236.270 ;
        RECT 1948.930 1233.490 1950.110 1234.670 ;
        RECT 1948.930 1055.090 1950.110 1056.270 ;
        RECT 1948.930 1053.490 1950.110 1054.670 ;
        RECT 1948.930 875.090 1950.110 876.270 ;
        RECT 1948.930 873.490 1950.110 874.670 ;
        RECT 1948.930 695.090 1950.110 696.270 ;
        RECT 1948.930 693.490 1950.110 694.670 ;
        RECT 1948.930 515.090 1950.110 516.270 ;
        RECT 1948.930 513.490 1950.110 514.670 ;
        RECT 1948.930 335.090 1950.110 336.270 ;
        RECT 1948.930 333.490 1950.110 334.670 ;
        RECT 1948.930 155.090 1950.110 156.270 ;
        RECT 1948.930 153.490 1950.110 154.670 ;
        RECT 1948.930 -35.110 1950.110 -33.930 ;
        RECT 1948.930 -36.710 1950.110 -35.530 ;
        RECT 2128.930 3555.210 2130.110 3556.390 ;
        RECT 2128.930 3553.610 2130.110 3554.790 ;
        RECT 2128.930 3395.090 2130.110 3396.270 ;
        RECT 2128.930 3393.490 2130.110 3394.670 ;
        RECT 2128.930 3215.090 2130.110 3216.270 ;
        RECT 2128.930 3213.490 2130.110 3214.670 ;
        RECT 2128.930 3035.090 2130.110 3036.270 ;
        RECT 2128.930 3033.490 2130.110 3034.670 ;
        RECT 2128.930 2855.090 2130.110 2856.270 ;
        RECT 2128.930 2853.490 2130.110 2854.670 ;
        RECT 2128.930 2675.090 2130.110 2676.270 ;
        RECT 2128.930 2673.490 2130.110 2674.670 ;
        RECT 2128.930 2495.090 2130.110 2496.270 ;
        RECT 2128.930 2493.490 2130.110 2494.670 ;
        RECT 2128.930 2315.090 2130.110 2316.270 ;
        RECT 2128.930 2313.490 2130.110 2314.670 ;
        RECT 2128.930 2135.090 2130.110 2136.270 ;
        RECT 2128.930 2133.490 2130.110 2134.670 ;
        RECT 2128.930 1955.090 2130.110 1956.270 ;
        RECT 2128.930 1953.490 2130.110 1954.670 ;
        RECT 2128.930 1775.090 2130.110 1776.270 ;
        RECT 2128.930 1773.490 2130.110 1774.670 ;
        RECT 2128.930 1595.090 2130.110 1596.270 ;
        RECT 2128.930 1593.490 2130.110 1594.670 ;
        RECT 2128.930 1415.090 2130.110 1416.270 ;
        RECT 2128.930 1413.490 2130.110 1414.670 ;
        RECT 2128.930 1235.090 2130.110 1236.270 ;
        RECT 2128.930 1233.490 2130.110 1234.670 ;
        RECT 2128.930 1055.090 2130.110 1056.270 ;
        RECT 2128.930 1053.490 2130.110 1054.670 ;
        RECT 2128.930 875.090 2130.110 876.270 ;
        RECT 2128.930 873.490 2130.110 874.670 ;
        RECT 2128.930 695.090 2130.110 696.270 ;
        RECT 2128.930 693.490 2130.110 694.670 ;
        RECT 2128.930 515.090 2130.110 516.270 ;
        RECT 2128.930 513.490 2130.110 514.670 ;
        RECT 2128.930 335.090 2130.110 336.270 ;
        RECT 2128.930 333.490 2130.110 334.670 ;
        RECT 2128.930 155.090 2130.110 156.270 ;
        RECT 2128.930 153.490 2130.110 154.670 ;
        RECT 2128.930 -35.110 2130.110 -33.930 ;
        RECT 2128.930 -36.710 2130.110 -35.530 ;
        RECT 2308.930 3555.210 2310.110 3556.390 ;
        RECT 2308.930 3553.610 2310.110 3554.790 ;
        RECT 2308.930 3395.090 2310.110 3396.270 ;
        RECT 2308.930 3393.490 2310.110 3394.670 ;
        RECT 2308.930 3215.090 2310.110 3216.270 ;
        RECT 2308.930 3213.490 2310.110 3214.670 ;
        RECT 2308.930 3035.090 2310.110 3036.270 ;
        RECT 2308.930 3033.490 2310.110 3034.670 ;
        RECT 2308.930 2855.090 2310.110 2856.270 ;
        RECT 2308.930 2853.490 2310.110 2854.670 ;
        RECT 2308.930 2675.090 2310.110 2676.270 ;
        RECT 2308.930 2673.490 2310.110 2674.670 ;
        RECT 2308.930 2495.090 2310.110 2496.270 ;
        RECT 2308.930 2493.490 2310.110 2494.670 ;
        RECT 2308.930 2315.090 2310.110 2316.270 ;
        RECT 2308.930 2313.490 2310.110 2314.670 ;
        RECT 2308.930 2135.090 2310.110 2136.270 ;
        RECT 2308.930 2133.490 2310.110 2134.670 ;
        RECT 2308.930 1955.090 2310.110 1956.270 ;
        RECT 2308.930 1953.490 2310.110 1954.670 ;
        RECT 2308.930 1775.090 2310.110 1776.270 ;
        RECT 2308.930 1773.490 2310.110 1774.670 ;
        RECT 2308.930 1595.090 2310.110 1596.270 ;
        RECT 2308.930 1593.490 2310.110 1594.670 ;
        RECT 2308.930 1415.090 2310.110 1416.270 ;
        RECT 2308.930 1413.490 2310.110 1414.670 ;
        RECT 2308.930 1235.090 2310.110 1236.270 ;
        RECT 2308.930 1233.490 2310.110 1234.670 ;
        RECT 2308.930 1055.090 2310.110 1056.270 ;
        RECT 2308.930 1053.490 2310.110 1054.670 ;
        RECT 2308.930 875.090 2310.110 876.270 ;
        RECT 2308.930 873.490 2310.110 874.670 ;
        RECT 2308.930 695.090 2310.110 696.270 ;
        RECT 2308.930 693.490 2310.110 694.670 ;
        RECT 2308.930 515.090 2310.110 516.270 ;
        RECT 2308.930 513.490 2310.110 514.670 ;
        RECT 2308.930 335.090 2310.110 336.270 ;
        RECT 2308.930 333.490 2310.110 334.670 ;
        RECT 2308.930 155.090 2310.110 156.270 ;
        RECT 2308.930 153.490 2310.110 154.670 ;
        RECT 2308.930 -35.110 2310.110 -33.930 ;
        RECT 2308.930 -36.710 2310.110 -35.530 ;
        RECT 2488.930 3555.210 2490.110 3556.390 ;
        RECT 2488.930 3553.610 2490.110 3554.790 ;
        RECT 2488.930 3395.090 2490.110 3396.270 ;
        RECT 2488.930 3393.490 2490.110 3394.670 ;
        RECT 2488.930 3215.090 2490.110 3216.270 ;
        RECT 2488.930 3213.490 2490.110 3214.670 ;
        RECT 2488.930 3035.090 2490.110 3036.270 ;
        RECT 2488.930 3033.490 2490.110 3034.670 ;
        RECT 2488.930 2855.090 2490.110 2856.270 ;
        RECT 2488.930 2853.490 2490.110 2854.670 ;
        RECT 2488.930 2675.090 2490.110 2676.270 ;
        RECT 2488.930 2673.490 2490.110 2674.670 ;
        RECT 2488.930 2495.090 2490.110 2496.270 ;
        RECT 2488.930 2493.490 2490.110 2494.670 ;
        RECT 2488.930 2315.090 2490.110 2316.270 ;
        RECT 2488.930 2313.490 2490.110 2314.670 ;
        RECT 2488.930 2135.090 2490.110 2136.270 ;
        RECT 2488.930 2133.490 2490.110 2134.670 ;
        RECT 2488.930 1955.090 2490.110 1956.270 ;
        RECT 2488.930 1953.490 2490.110 1954.670 ;
        RECT 2488.930 1775.090 2490.110 1776.270 ;
        RECT 2488.930 1773.490 2490.110 1774.670 ;
        RECT 2488.930 1595.090 2490.110 1596.270 ;
        RECT 2488.930 1593.490 2490.110 1594.670 ;
        RECT 2488.930 1415.090 2490.110 1416.270 ;
        RECT 2488.930 1413.490 2490.110 1414.670 ;
        RECT 2488.930 1235.090 2490.110 1236.270 ;
        RECT 2488.930 1233.490 2490.110 1234.670 ;
        RECT 2488.930 1055.090 2490.110 1056.270 ;
        RECT 2488.930 1053.490 2490.110 1054.670 ;
        RECT 2488.930 875.090 2490.110 876.270 ;
        RECT 2488.930 873.490 2490.110 874.670 ;
        RECT 2488.930 695.090 2490.110 696.270 ;
        RECT 2488.930 693.490 2490.110 694.670 ;
        RECT 2488.930 515.090 2490.110 516.270 ;
        RECT 2488.930 513.490 2490.110 514.670 ;
        RECT 2488.930 335.090 2490.110 336.270 ;
        RECT 2488.930 333.490 2490.110 334.670 ;
        RECT 2488.930 155.090 2490.110 156.270 ;
        RECT 2488.930 153.490 2490.110 154.670 ;
        RECT 2488.930 -35.110 2490.110 -33.930 ;
        RECT 2488.930 -36.710 2490.110 -35.530 ;
        RECT 2668.930 3555.210 2670.110 3556.390 ;
        RECT 2668.930 3553.610 2670.110 3554.790 ;
        RECT 2668.930 3395.090 2670.110 3396.270 ;
        RECT 2668.930 3393.490 2670.110 3394.670 ;
        RECT 2668.930 3215.090 2670.110 3216.270 ;
        RECT 2668.930 3213.490 2670.110 3214.670 ;
        RECT 2668.930 3035.090 2670.110 3036.270 ;
        RECT 2668.930 3033.490 2670.110 3034.670 ;
        RECT 2668.930 2855.090 2670.110 2856.270 ;
        RECT 2668.930 2853.490 2670.110 2854.670 ;
        RECT 2668.930 2675.090 2670.110 2676.270 ;
        RECT 2668.930 2673.490 2670.110 2674.670 ;
        RECT 2668.930 2495.090 2670.110 2496.270 ;
        RECT 2668.930 2493.490 2670.110 2494.670 ;
        RECT 2668.930 2315.090 2670.110 2316.270 ;
        RECT 2668.930 2313.490 2670.110 2314.670 ;
        RECT 2668.930 2135.090 2670.110 2136.270 ;
        RECT 2668.930 2133.490 2670.110 2134.670 ;
        RECT 2668.930 1955.090 2670.110 1956.270 ;
        RECT 2668.930 1953.490 2670.110 1954.670 ;
        RECT 2668.930 1775.090 2670.110 1776.270 ;
        RECT 2668.930 1773.490 2670.110 1774.670 ;
        RECT 2668.930 1595.090 2670.110 1596.270 ;
        RECT 2668.930 1593.490 2670.110 1594.670 ;
        RECT 2668.930 1415.090 2670.110 1416.270 ;
        RECT 2668.930 1413.490 2670.110 1414.670 ;
        RECT 2668.930 1235.090 2670.110 1236.270 ;
        RECT 2668.930 1233.490 2670.110 1234.670 ;
        RECT 2668.930 1055.090 2670.110 1056.270 ;
        RECT 2668.930 1053.490 2670.110 1054.670 ;
        RECT 2668.930 875.090 2670.110 876.270 ;
        RECT 2668.930 873.490 2670.110 874.670 ;
        RECT 2668.930 695.090 2670.110 696.270 ;
        RECT 2668.930 693.490 2670.110 694.670 ;
        RECT 2668.930 515.090 2670.110 516.270 ;
        RECT 2668.930 513.490 2670.110 514.670 ;
        RECT 2668.930 335.090 2670.110 336.270 ;
        RECT 2668.930 333.490 2670.110 334.670 ;
        RECT 2668.930 155.090 2670.110 156.270 ;
        RECT 2668.930 153.490 2670.110 154.670 ;
        RECT 2668.930 -35.110 2670.110 -33.930 ;
        RECT 2668.930 -36.710 2670.110 -35.530 ;
        RECT 2848.930 3555.210 2850.110 3556.390 ;
        RECT 2848.930 3553.610 2850.110 3554.790 ;
        RECT 2848.930 3395.090 2850.110 3396.270 ;
        RECT 2848.930 3393.490 2850.110 3394.670 ;
        RECT 2848.930 3215.090 2850.110 3216.270 ;
        RECT 2848.930 3213.490 2850.110 3214.670 ;
        RECT 2848.930 3035.090 2850.110 3036.270 ;
        RECT 2848.930 3033.490 2850.110 3034.670 ;
        RECT 2848.930 2855.090 2850.110 2856.270 ;
        RECT 2848.930 2853.490 2850.110 2854.670 ;
        RECT 2848.930 2675.090 2850.110 2676.270 ;
        RECT 2848.930 2673.490 2850.110 2674.670 ;
        RECT 2848.930 2495.090 2850.110 2496.270 ;
        RECT 2848.930 2493.490 2850.110 2494.670 ;
        RECT 2848.930 2315.090 2850.110 2316.270 ;
        RECT 2848.930 2313.490 2850.110 2314.670 ;
        RECT 2848.930 2135.090 2850.110 2136.270 ;
        RECT 2848.930 2133.490 2850.110 2134.670 ;
        RECT 2848.930 1955.090 2850.110 1956.270 ;
        RECT 2848.930 1953.490 2850.110 1954.670 ;
        RECT 2848.930 1775.090 2850.110 1776.270 ;
        RECT 2848.930 1773.490 2850.110 1774.670 ;
        RECT 2848.930 1595.090 2850.110 1596.270 ;
        RECT 2848.930 1593.490 2850.110 1594.670 ;
        RECT 2848.930 1415.090 2850.110 1416.270 ;
        RECT 2848.930 1413.490 2850.110 1414.670 ;
        RECT 2848.930 1235.090 2850.110 1236.270 ;
        RECT 2848.930 1233.490 2850.110 1234.670 ;
        RECT 2848.930 1055.090 2850.110 1056.270 ;
        RECT 2848.930 1053.490 2850.110 1054.670 ;
        RECT 2848.930 875.090 2850.110 876.270 ;
        RECT 2848.930 873.490 2850.110 874.670 ;
        RECT 2848.930 695.090 2850.110 696.270 ;
        RECT 2848.930 693.490 2850.110 694.670 ;
        RECT 2848.930 515.090 2850.110 516.270 ;
        RECT 2848.930 513.490 2850.110 514.670 ;
        RECT 2848.930 335.090 2850.110 336.270 ;
        RECT 2848.930 333.490 2850.110 334.670 ;
        RECT 2848.930 155.090 2850.110 156.270 ;
        RECT 2848.930 153.490 2850.110 154.670 ;
        RECT 2848.930 -35.110 2850.110 -33.930 ;
        RECT 2848.930 -36.710 2850.110 -35.530 ;
        RECT 2959.710 3555.210 2960.890 3556.390 ;
        RECT 2959.710 3553.610 2960.890 3554.790 ;
        RECT 2959.710 3395.090 2960.890 3396.270 ;
        RECT 2959.710 3393.490 2960.890 3394.670 ;
        RECT 2959.710 3215.090 2960.890 3216.270 ;
        RECT 2959.710 3213.490 2960.890 3214.670 ;
        RECT 2959.710 3035.090 2960.890 3036.270 ;
        RECT 2959.710 3033.490 2960.890 3034.670 ;
        RECT 2959.710 2855.090 2960.890 2856.270 ;
        RECT 2959.710 2853.490 2960.890 2854.670 ;
        RECT 2959.710 2675.090 2960.890 2676.270 ;
        RECT 2959.710 2673.490 2960.890 2674.670 ;
        RECT 2959.710 2495.090 2960.890 2496.270 ;
        RECT 2959.710 2493.490 2960.890 2494.670 ;
        RECT 2959.710 2315.090 2960.890 2316.270 ;
        RECT 2959.710 2313.490 2960.890 2314.670 ;
        RECT 2959.710 2135.090 2960.890 2136.270 ;
        RECT 2959.710 2133.490 2960.890 2134.670 ;
        RECT 2959.710 1955.090 2960.890 1956.270 ;
        RECT 2959.710 1953.490 2960.890 1954.670 ;
        RECT 2959.710 1775.090 2960.890 1776.270 ;
        RECT 2959.710 1773.490 2960.890 1774.670 ;
        RECT 2959.710 1595.090 2960.890 1596.270 ;
        RECT 2959.710 1593.490 2960.890 1594.670 ;
        RECT 2959.710 1415.090 2960.890 1416.270 ;
        RECT 2959.710 1413.490 2960.890 1414.670 ;
        RECT 2959.710 1235.090 2960.890 1236.270 ;
        RECT 2959.710 1233.490 2960.890 1234.670 ;
        RECT 2959.710 1055.090 2960.890 1056.270 ;
        RECT 2959.710 1053.490 2960.890 1054.670 ;
        RECT 2959.710 875.090 2960.890 876.270 ;
        RECT 2959.710 873.490 2960.890 874.670 ;
        RECT 2959.710 695.090 2960.890 696.270 ;
        RECT 2959.710 693.490 2960.890 694.670 ;
        RECT 2959.710 515.090 2960.890 516.270 ;
        RECT 2959.710 513.490 2960.890 514.670 ;
        RECT 2959.710 335.090 2960.890 336.270 ;
        RECT 2959.710 333.490 2960.890 334.670 ;
        RECT 2959.710 155.090 2960.890 156.270 ;
        RECT 2959.710 153.490 2960.890 154.670 ;
        RECT 2959.710 -35.110 2960.890 -33.930 ;
        RECT 2959.710 -36.710 2960.890 -35.530 ;
      LAYER met5 ;
        RECT -42.180 3556.500 -39.180 3556.510 ;
        RECT 148.020 3556.500 151.020 3556.510 ;
        RECT 328.020 3556.500 331.020 3556.510 ;
        RECT 508.020 3556.500 511.020 3556.510 ;
        RECT 688.020 3556.500 691.020 3556.510 ;
        RECT 868.020 3556.500 871.020 3556.510 ;
        RECT 1048.020 3556.500 1051.020 3556.510 ;
        RECT 1228.020 3556.500 1231.020 3556.510 ;
        RECT 1408.020 3556.500 1411.020 3556.510 ;
        RECT 1588.020 3556.500 1591.020 3556.510 ;
        RECT 1768.020 3556.500 1771.020 3556.510 ;
        RECT 1948.020 3556.500 1951.020 3556.510 ;
        RECT 2128.020 3556.500 2131.020 3556.510 ;
        RECT 2308.020 3556.500 2311.020 3556.510 ;
        RECT 2488.020 3556.500 2491.020 3556.510 ;
        RECT 2668.020 3556.500 2671.020 3556.510 ;
        RECT 2848.020 3556.500 2851.020 3556.510 ;
        RECT 2958.800 3556.500 2961.800 3556.510 ;
        RECT -42.180 3553.500 2961.800 3556.500 ;
        RECT -42.180 3553.490 -39.180 3553.500 ;
        RECT 148.020 3553.490 151.020 3553.500 ;
        RECT 328.020 3553.490 331.020 3553.500 ;
        RECT 508.020 3553.490 511.020 3553.500 ;
        RECT 688.020 3553.490 691.020 3553.500 ;
        RECT 868.020 3553.490 871.020 3553.500 ;
        RECT 1048.020 3553.490 1051.020 3553.500 ;
        RECT 1228.020 3553.490 1231.020 3553.500 ;
        RECT 1408.020 3553.490 1411.020 3553.500 ;
        RECT 1588.020 3553.490 1591.020 3553.500 ;
        RECT 1768.020 3553.490 1771.020 3553.500 ;
        RECT 1948.020 3553.490 1951.020 3553.500 ;
        RECT 2128.020 3553.490 2131.020 3553.500 ;
        RECT 2308.020 3553.490 2311.020 3553.500 ;
        RECT 2488.020 3553.490 2491.020 3553.500 ;
        RECT 2668.020 3553.490 2671.020 3553.500 ;
        RECT 2848.020 3553.490 2851.020 3553.500 ;
        RECT 2958.800 3553.490 2961.800 3553.500 ;
        RECT -42.180 3396.380 -39.180 3396.390 ;
        RECT 148.020 3396.380 151.020 3396.390 ;
        RECT 328.020 3396.380 331.020 3396.390 ;
        RECT 508.020 3396.380 511.020 3396.390 ;
        RECT 688.020 3396.380 691.020 3396.390 ;
        RECT 868.020 3396.380 871.020 3396.390 ;
        RECT 1048.020 3396.380 1051.020 3396.390 ;
        RECT 1228.020 3396.380 1231.020 3396.390 ;
        RECT 1408.020 3396.380 1411.020 3396.390 ;
        RECT 1588.020 3396.380 1591.020 3396.390 ;
        RECT 1768.020 3396.380 1771.020 3396.390 ;
        RECT 1948.020 3396.380 1951.020 3396.390 ;
        RECT 2128.020 3396.380 2131.020 3396.390 ;
        RECT 2308.020 3396.380 2311.020 3396.390 ;
        RECT 2488.020 3396.380 2491.020 3396.390 ;
        RECT 2668.020 3396.380 2671.020 3396.390 ;
        RECT 2848.020 3396.380 2851.020 3396.390 ;
        RECT 2958.800 3396.380 2961.800 3396.390 ;
        RECT -42.180 3393.380 2961.800 3396.380 ;
        RECT -42.180 3393.370 -39.180 3393.380 ;
        RECT 148.020 3393.370 151.020 3393.380 ;
        RECT 328.020 3393.370 331.020 3393.380 ;
        RECT 508.020 3393.370 511.020 3393.380 ;
        RECT 688.020 3393.370 691.020 3393.380 ;
        RECT 868.020 3393.370 871.020 3393.380 ;
        RECT 1048.020 3393.370 1051.020 3393.380 ;
        RECT 1228.020 3393.370 1231.020 3393.380 ;
        RECT 1408.020 3393.370 1411.020 3393.380 ;
        RECT 1588.020 3393.370 1591.020 3393.380 ;
        RECT 1768.020 3393.370 1771.020 3393.380 ;
        RECT 1948.020 3393.370 1951.020 3393.380 ;
        RECT 2128.020 3393.370 2131.020 3393.380 ;
        RECT 2308.020 3393.370 2311.020 3393.380 ;
        RECT 2488.020 3393.370 2491.020 3393.380 ;
        RECT 2668.020 3393.370 2671.020 3393.380 ;
        RECT 2848.020 3393.370 2851.020 3393.380 ;
        RECT 2958.800 3393.370 2961.800 3393.380 ;
        RECT -42.180 3216.380 -39.180 3216.390 ;
        RECT 148.020 3216.380 151.020 3216.390 ;
        RECT 328.020 3216.380 331.020 3216.390 ;
        RECT 508.020 3216.380 511.020 3216.390 ;
        RECT 688.020 3216.380 691.020 3216.390 ;
        RECT 868.020 3216.380 871.020 3216.390 ;
        RECT 1048.020 3216.380 1051.020 3216.390 ;
        RECT 1228.020 3216.380 1231.020 3216.390 ;
        RECT 1408.020 3216.380 1411.020 3216.390 ;
        RECT 1588.020 3216.380 1591.020 3216.390 ;
        RECT 1768.020 3216.380 1771.020 3216.390 ;
        RECT 1948.020 3216.380 1951.020 3216.390 ;
        RECT 2128.020 3216.380 2131.020 3216.390 ;
        RECT 2308.020 3216.380 2311.020 3216.390 ;
        RECT 2488.020 3216.380 2491.020 3216.390 ;
        RECT 2668.020 3216.380 2671.020 3216.390 ;
        RECT 2848.020 3216.380 2851.020 3216.390 ;
        RECT 2958.800 3216.380 2961.800 3216.390 ;
        RECT -42.180 3213.380 2961.800 3216.380 ;
        RECT -42.180 3213.370 -39.180 3213.380 ;
        RECT 148.020 3213.370 151.020 3213.380 ;
        RECT 328.020 3213.370 331.020 3213.380 ;
        RECT 508.020 3213.370 511.020 3213.380 ;
        RECT 688.020 3213.370 691.020 3213.380 ;
        RECT 868.020 3213.370 871.020 3213.380 ;
        RECT 1048.020 3213.370 1051.020 3213.380 ;
        RECT 1228.020 3213.370 1231.020 3213.380 ;
        RECT 1408.020 3213.370 1411.020 3213.380 ;
        RECT 1588.020 3213.370 1591.020 3213.380 ;
        RECT 1768.020 3213.370 1771.020 3213.380 ;
        RECT 1948.020 3213.370 1951.020 3213.380 ;
        RECT 2128.020 3213.370 2131.020 3213.380 ;
        RECT 2308.020 3213.370 2311.020 3213.380 ;
        RECT 2488.020 3213.370 2491.020 3213.380 ;
        RECT 2668.020 3213.370 2671.020 3213.380 ;
        RECT 2848.020 3213.370 2851.020 3213.380 ;
        RECT 2958.800 3213.370 2961.800 3213.380 ;
        RECT -42.180 3036.380 -39.180 3036.390 ;
        RECT 148.020 3036.380 151.020 3036.390 ;
        RECT 328.020 3036.380 331.020 3036.390 ;
        RECT 508.020 3036.380 511.020 3036.390 ;
        RECT 688.020 3036.380 691.020 3036.390 ;
        RECT 868.020 3036.380 871.020 3036.390 ;
        RECT 1048.020 3036.380 1051.020 3036.390 ;
        RECT 1228.020 3036.380 1231.020 3036.390 ;
        RECT 1408.020 3036.380 1411.020 3036.390 ;
        RECT 1588.020 3036.380 1591.020 3036.390 ;
        RECT 1768.020 3036.380 1771.020 3036.390 ;
        RECT 1948.020 3036.380 1951.020 3036.390 ;
        RECT 2128.020 3036.380 2131.020 3036.390 ;
        RECT 2308.020 3036.380 2311.020 3036.390 ;
        RECT 2488.020 3036.380 2491.020 3036.390 ;
        RECT 2668.020 3036.380 2671.020 3036.390 ;
        RECT 2848.020 3036.380 2851.020 3036.390 ;
        RECT 2958.800 3036.380 2961.800 3036.390 ;
        RECT -42.180 3033.380 2961.800 3036.380 ;
        RECT -42.180 3033.370 -39.180 3033.380 ;
        RECT 148.020 3033.370 151.020 3033.380 ;
        RECT 328.020 3033.370 331.020 3033.380 ;
        RECT 508.020 3033.370 511.020 3033.380 ;
        RECT 688.020 3033.370 691.020 3033.380 ;
        RECT 868.020 3033.370 871.020 3033.380 ;
        RECT 1048.020 3033.370 1051.020 3033.380 ;
        RECT 1228.020 3033.370 1231.020 3033.380 ;
        RECT 1408.020 3033.370 1411.020 3033.380 ;
        RECT 1588.020 3033.370 1591.020 3033.380 ;
        RECT 1768.020 3033.370 1771.020 3033.380 ;
        RECT 1948.020 3033.370 1951.020 3033.380 ;
        RECT 2128.020 3033.370 2131.020 3033.380 ;
        RECT 2308.020 3033.370 2311.020 3033.380 ;
        RECT 2488.020 3033.370 2491.020 3033.380 ;
        RECT 2668.020 3033.370 2671.020 3033.380 ;
        RECT 2848.020 3033.370 2851.020 3033.380 ;
        RECT 2958.800 3033.370 2961.800 3033.380 ;
        RECT -42.180 2856.380 -39.180 2856.390 ;
        RECT 148.020 2856.380 151.020 2856.390 ;
        RECT 328.020 2856.380 331.020 2856.390 ;
        RECT 508.020 2856.380 511.020 2856.390 ;
        RECT 688.020 2856.380 691.020 2856.390 ;
        RECT 868.020 2856.380 871.020 2856.390 ;
        RECT 1048.020 2856.380 1051.020 2856.390 ;
        RECT 1228.020 2856.380 1231.020 2856.390 ;
        RECT 1408.020 2856.380 1411.020 2856.390 ;
        RECT 1588.020 2856.380 1591.020 2856.390 ;
        RECT 1768.020 2856.380 1771.020 2856.390 ;
        RECT 1948.020 2856.380 1951.020 2856.390 ;
        RECT 2128.020 2856.380 2131.020 2856.390 ;
        RECT 2308.020 2856.380 2311.020 2856.390 ;
        RECT 2488.020 2856.380 2491.020 2856.390 ;
        RECT 2668.020 2856.380 2671.020 2856.390 ;
        RECT 2848.020 2856.380 2851.020 2856.390 ;
        RECT 2958.800 2856.380 2961.800 2856.390 ;
        RECT -42.180 2853.380 2961.800 2856.380 ;
        RECT -42.180 2853.370 -39.180 2853.380 ;
        RECT 148.020 2853.370 151.020 2853.380 ;
        RECT 328.020 2853.370 331.020 2853.380 ;
        RECT 508.020 2853.370 511.020 2853.380 ;
        RECT 688.020 2853.370 691.020 2853.380 ;
        RECT 868.020 2853.370 871.020 2853.380 ;
        RECT 1048.020 2853.370 1051.020 2853.380 ;
        RECT 1228.020 2853.370 1231.020 2853.380 ;
        RECT 1408.020 2853.370 1411.020 2853.380 ;
        RECT 1588.020 2853.370 1591.020 2853.380 ;
        RECT 1768.020 2853.370 1771.020 2853.380 ;
        RECT 1948.020 2853.370 1951.020 2853.380 ;
        RECT 2128.020 2853.370 2131.020 2853.380 ;
        RECT 2308.020 2853.370 2311.020 2853.380 ;
        RECT 2488.020 2853.370 2491.020 2853.380 ;
        RECT 2668.020 2853.370 2671.020 2853.380 ;
        RECT 2848.020 2853.370 2851.020 2853.380 ;
        RECT 2958.800 2853.370 2961.800 2853.380 ;
        RECT -42.180 2676.380 -39.180 2676.390 ;
        RECT 148.020 2676.380 151.020 2676.390 ;
        RECT 328.020 2676.380 331.020 2676.390 ;
        RECT 508.020 2676.380 511.020 2676.390 ;
        RECT 688.020 2676.380 691.020 2676.390 ;
        RECT 868.020 2676.380 871.020 2676.390 ;
        RECT 1048.020 2676.380 1051.020 2676.390 ;
        RECT 1228.020 2676.380 1231.020 2676.390 ;
        RECT 1408.020 2676.380 1411.020 2676.390 ;
        RECT 1588.020 2676.380 1591.020 2676.390 ;
        RECT 1768.020 2676.380 1771.020 2676.390 ;
        RECT 1948.020 2676.380 1951.020 2676.390 ;
        RECT 2128.020 2676.380 2131.020 2676.390 ;
        RECT 2308.020 2676.380 2311.020 2676.390 ;
        RECT 2488.020 2676.380 2491.020 2676.390 ;
        RECT 2668.020 2676.380 2671.020 2676.390 ;
        RECT 2848.020 2676.380 2851.020 2676.390 ;
        RECT 2958.800 2676.380 2961.800 2676.390 ;
        RECT -42.180 2673.380 2961.800 2676.380 ;
        RECT -42.180 2673.370 -39.180 2673.380 ;
        RECT 148.020 2673.370 151.020 2673.380 ;
        RECT 328.020 2673.370 331.020 2673.380 ;
        RECT 508.020 2673.370 511.020 2673.380 ;
        RECT 688.020 2673.370 691.020 2673.380 ;
        RECT 868.020 2673.370 871.020 2673.380 ;
        RECT 1048.020 2673.370 1051.020 2673.380 ;
        RECT 1228.020 2673.370 1231.020 2673.380 ;
        RECT 1408.020 2673.370 1411.020 2673.380 ;
        RECT 1588.020 2673.370 1591.020 2673.380 ;
        RECT 1768.020 2673.370 1771.020 2673.380 ;
        RECT 1948.020 2673.370 1951.020 2673.380 ;
        RECT 2128.020 2673.370 2131.020 2673.380 ;
        RECT 2308.020 2673.370 2311.020 2673.380 ;
        RECT 2488.020 2673.370 2491.020 2673.380 ;
        RECT 2668.020 2673.370 2671.020 2673.380 ;
        RECT 2848.020 2673.370 2851.020 2673.380 ;
        RECT 2958.800 2673.370 2961.800 2673.380 ;
        RECT -42.180 2496.380 -39.180 2496.390 ;
        RECT 148.020 2496.380 151.020 2496.390 ;
        RECT 328.020 2496.380 331.020 2496.390 ;
        RECT 508.020 2496.380 511.020 2496.390 ;
        RECT 688.020 2496.380 691.020 2496.390 ;
        RECT 868.020 2496.380 871.020 2496.390 ;
        RECT 1048.020 2496.380 1051.020 2496.390 ;
        RECT 1228.020 2496.380 1231.020 2496.390 ;
        RECT 1408.020 2496.380 1411.020 2496.390 ;
        RECT 1588.020 2496.380 1591.020 2496.390 ;
        RECT 1768.020 2496.380 1771.020 2496.390 ;
        RECT 1948.020 2496.380 1951.020 2496.390 ;
        RECT 2128.020 2496.380 2131.020 2496.390 ;
        RECT 2308.020 2496.380 2311.020 2496.390 ;
        RECT 2488.020 2496.380 2491.020 2496.390 ;
        RECT 2668.020 2496.380 2671.020 2496.390 ;
        RECT 2848.020 2496.380 2851.020 2496.390 ;
        RECT 2958.800 2496.380 2961.800 2496.390 ;
        RECT -42.180 2493.380 2961.800 2496.380 ;
        RECT -42.180 2493.370 -39.180 2493.380 ;
        RECT 148.020 2493.370 151.020 2493.380 ;
        RECT 328.020 2493.370 331.020 2493.380 ;
        RECT 508.020 2493.370 511.020 2493.380 ;
        RECT 688.020 2493.370 691.020 2493.380 ;
        RECT 868.020 2493.370 871.020 2493.380 ;
        RECT 1048.020 2493.370 1051.020 2493.380 ;
        RECT 1228.020 2493.370 1231.020 2493.380 ;
        RECT 1408.020 2493.370 1411.020 2493.380 ;
        RECT 1588.020 2493.370 1591.020 2493.380 ;
        RECT 1768.020 2493.370 1771.020 2493.380 ;
        RECT 1948.020 2493.370 1951.020 2493.380 ;
        RECT 2128.020 2493.370 2131.020 2493.380 ;
        RECT 2308.020 2493.370 2311.020 2493.380 ;
        RECT 2488.020 2493.370 2491.020 2493.380 ;
        RECT 2668.020 2493.370 2671.020 2493.380 ;
        RECT 2848.020 2493.370 2851.020 2493.380 ;
        RECT 2958.800 2493.370 2961.800 2493.380 ;
        RECT -42.180 2316.380 -39.180 2316.390 ;
        RECT 148.020 2316.380 151.020 2316.390 ;
        RECT 328.020 2316.380 331.020 2316.390 ;
        RECT 508.020 2316.380 511.020 2316.390 ;
        RECT 688.020 2316.380 691.020 2316.390 ;
        RECT 868.020 2316.380 871.020 2316.390 ;
        RECT 1048.020 2316.380 1051.020 2316.390 ;
        RECT 1228.020 2316.380 1231.020 2316.390 ;
        RECT 1408.020 2316.380 1411.020 2316.390 ;
        RECT 1588.020 2316.380 1591.020 2316.390 ;
        RECT 1768.020 2316.380 1771.020 2316.390 ;
        RECT 1948.020 2316.380 1951.020 2316.390 ;
        RECT 2128.020 2316.380 2131.020 2316.390 ;
        RECT 2308.020 2316.380 2311.020 2316.390 ;
        RECT 2488.020 2316.380 2491.020 2316.390 ;
        RECT 2668.020 2316.380 2671.020 2316.390 ;
        RECT 2848.020 2316.380 2851.020 2316.390 ;
        RECT 2958.800 2316.380 2961.800 2316.390 ;
        RECT -42.180 2313.380 2961.800 2316.380 ;
        RECT -42.180 2313.370 -39.180 2313.380 ;
        RECT 148.020 2313.370 151.020 2313.380 ;
        RECT 328.020 2313.370 331.020 2313.380 ;
        RECT 508.020 2313.370 511.020 2313.380 ;
        RECT 688.020 2313.370 691.020 2313.380 ;
        RECT 868.020 2313.370 871.020 2313.380 ;
        RECT 1048.020 2313.370 1051.020 2313.380 ;
        RECT 1228.020 2313.370 1231.020 2313.380 ;
        RECT 1408.020 2313.370 1411.020 2313.380 ;
        RECT 1588.020 2313.370 1591.020 2313.380 ;
        RECT 1768.020 2313.370 1771.020 2313.380 ;
        RECT 1948.020 2313.370 1951.020 2313.380 ;
        RECT 2128.020 2313.370 2131.020 2313.380 ;
        RECT 2308.020 2313.370 2311.020 2313.380 ;
        RECT 2488.020 2313.370 2491.020 2313.380 ;
        RECT 2668.020 2313.370 2671.020 2313.380 ;
        RECT 2848.020 2313.370 2851.020 2313.380 ;
        RECT 2958.800 2313.370 2961.800 2313.380 ;
        RECT -42.180 2136.380 -39.180 2136.390 ;
        RECT 148.020 2136.380 151.020 2136.390 ;
        RECT 328.020 2136.380 331.020 2136.390 ;
        RECT 508.020 2136.380 511.020 2136.390 ;
        RECT 688.020 2136.380 691.020 2136.390 ;
        RECT 868.020 2136.380 871.020 2136.390 ;
        RECT 1048.020 2136.380 1051.020 2136.390 ;
        RECT 1228.020 2136.380 1231.020 2136.390 ;
        RECT 1408.020 2136.380 1411.020 2136.390 ;
        RECT 1588.020 2136.380 1591.020 2136.390 ;
        RECT 1768.020 2136.380 1771.020 2136.390 ;
        RECT 1948.020 2136.380 1951.020 2136.390 ;
        RECT 2128.020 2136.380 2131.020 2136.390 ;
        RECT 2308.020 2136.380 2311.020 2136.390 ;
        RECT 2488.020 2136.380 2491.020 2136.390 ;
        RECT 2668.020 2136.380 2671.020 2136.390 ;
        RECT 2848.020 2136.380 2851.020 2136.390 ;
        RECT 2958.800 2136.380 2961.800 2136.390 ;
        RECT -42.180 2133.380 2961.800 2136.380 ;
        RECT -42.180 2133.370 -39.180 2133.380 ;
        RECT 148.020 2133.370 151.020 2133.380 ;
        RECT 328.020 2133.370 331.020 2133.380 ;
        RECT 508.020 2133.370 511.020 2133.380 ;
        RECT 688.020 2133.370 691.020 2133.380 ;
        RECT 868.020 2133.370 871.020 2133.380 ;
        RECT 1048.020 2133.370 1051.020 2133.380 ;
        RECT 1228.020 2133.370 1231.020 2133.380 ;
        RECT 1408.020 2133.370 1411.020 2133.380 ;
        RECT 1588.020 2133.370 1591.020 2133.380 ;
        RECT 1768.020 2133.370 1771.020 2133.380 ;
        RECT 1948.020 2133.370 1951.020 2133.380 ;
        RECT 2128.020 2133.370 2131.020 2133.380 ;
        RECT 2308.020 2133.370 2311.020 2133.380 ;
        RECT 2488.020 2133.370 2491.020 2133.380 ;
        RECT 2668.020 2133.370 2671.020 2133.380 ;
        RECT 2848.020 2133.370 2851.020 2133.380 ;
        RECT 2958.800 2133.370 2961.800 2133.380 ;
        RECT -42.180 1956.380 -39.180 1956.390 ;
        RECT 148.020 1956.380 151.020 1956.390 ;
        RECT 328.020 1956.380 331.020 1956.390 ;
        RECT 508.020 1956.380 511.020 1956.390 ;
        RECT 688.020 1956.380 691.020 1956.390 ;
        RECT 868.020 1956.380 871.020 1956.390 ;
        RECT 1048.020 1956.380 1051.020 1956.390 ;
        RECT 1228.020 1956.380 1231.020 1956.390 ;
        RECT 1408.020 1956.380 1411.020 1956.390 ;
        RECT 1588.020 1956.380 1591.020 1956.390 ;
        RECT 1768.020 1956.380 1771.020 1956.390 ;
        RECT 1948.020 1956.380 1951.020 1956.390 ;
        RECT 2128.020 1956.380 2131.020 1956.390 ;
        RECT 2308.020 1956.380 2311.020 1956.390 ;
        RECT 2488.020 1956.380 2491.020 1956.390 ;
        RECT 2668.020 1956.380 2671.020 1956.390 ;
        RECT 2848.020 1956.380 2851.020 1956.390 ;
        RECT 2958.800 1956.380 2961.800 1956.390 ;
        RECT -42.180 1953.380 2961.800 1956.380 ;
        RECT -42.180 1953.370 -39.180 1953.380 ;
        RECT 148.020 1953.370 151.020 1953.380 ;
        RECT 328.020 1953.370 331.020 1953.380 ;
        RECT 508.020 1953.370 511.020 1953.380 ;
        RECT 688.020 1953.370 691.020 1953.380 ;
        RECT 868.020 1953.370 871.020 1953.380 ;
        RECT 1048.020 1953.370 1051.020 1953.380 ;
        RECT 1228.020 1953.370 1231.020 1953.380 ;
        RECT 1408.020 1953.370 1411.020 1953.380 ;
        RECT 1588.020 1953.370 1591.020 1953.380 ;
        RECT 1768.020 1953.370 1771.020 1953.380 ;
        RECT 1948.020 1953.370 1951.020 1953.380 ;
        RECT 2128.020 1953.370 2131.020 1953.380 ;
        RECT 2308.020 1953.370 2311.020 1953.380 ;
        RECT 2488.020 1953.370 2491.020 1953.380 ;
        RECT 2668.020 1953.370 2671.020 1953.380 ;
        RECT 2848.020 1953.370 2851.020 1953.380 ;
        RECT 2958.800 1953.370 2961.800 1953.380 ;
        RECT -42.180 1776.380 -39.180 1776.390 ;
        RECT 148.020 1776.380 151.020 1776.390 ;
        RECT 328.020 1776.380 331.020 1776.390 ;
        RECT 508.020 1776.380 511.020 1776.390 ;
        RECT 688.020 1776.380 691.020 1776.390 ;
        RECT 868.020 1776.380 871.020 1776.390 ;
        RECT 1048.020 1776.380 1051.020 1776.390 ;
        RECT 1228.020 1776.380 1231.020 1776.390 ;
        RECT 1408.020 1776.380 1411.020 1776.390 ;
        RECT 1588.020 1776.380 1591.020 1776.390 ;
        RECT 1768.020 1776.380 1771.020 1776.390 ;
        RECT 1948.020 1776.380 1951.020 1776.390 ;
        RECT 2128.020 1776.380 2131.020 1776.390 ;
        RECT 2308.020 1776.380 2311.020 1776.390 ;
        RECT 2488.020 1776.380 2491.020 1776.390 ;
        RECT 2668.020 1776.380 2671.020 1776.390 ;
        RECT 2848.020 1776.380 2851.020 1776.390 ;
        RECT 2958.800 1776.380 2961.800 1776.390 ;
        RECT -42.180 1773.380 2961.800 1776.380 ;
        RECT -42.180 1773.370 -39.180 1773.380 ;
        RECT 148.020 1773.370 151.020 1773.380 ;
        RECT 328.020 1773.370 331.020 1773.380 ;
        RECT 508.020 1773.370 511.020 1773.380 ;
        RECT 688.020 1773.370 691.020 1773.380 ;
        RECT 868.020 1773.370 871.020 1773.380 ;
        RECT 1048.020 1773.370 1051.020 1773.380 ;
        RECT 1228.020 1773.370 1231.020 1773.380 ;
        RECT 1408.020 1773.370 1411.020 1773.380 ;
        RECT 1588.020 1773.370 1591.020 1773.380 ;
        RECT 1768.020 1773.370 1771.020 1773.380 ;
        RECT 1948.020 1773.370 1951.020 1773.380 ;
        RECT 2128.020 1773.370 2131.020 1773.380 ;
        RECT 2308.020 1773.370 2311.020 1773.380 ;
        RECT 2488.020 1773.370 2491.020 1773.380 ;
        RECT 2668.020 1773.370 2671.020 1773.380 ;
        RECT 2848.020 1773.370 2851.020 1773.380 ;
        RECT 2958.800 1773.370 2961.800 1773.380 ;
        RECT -42.180 1596.380 -39.180 1596.390 ;
        RECT 148.020 1596.380 151.020 1596.390 ;
        RECT 328.020 1596.380 331.020 1596.390 ;
        RECT 508.020 1596.380 511.020 1596.390 ;
        RECT 688.020 1596.380 691.020 1596.390 ;
        RECT 868.020 1596.380 871.020 1596.390 ;
        RECT 1048.020 1596.380 1051.020 1596.390 ;
        RECT 1228.020 1596.380 1231.020 1596.390 ;
        RECT 1408.020 1596.380 1411.020 1596.390 ;
        RECT 1588.020 1596.380 1591.020 1596.390 ;
        RECT 1768.020 1596.380 1771.020 1596.390 ;
        RECT 1948.020 1596.380 1951.020 1596.390 ;
        RECT 2128.020 1596.380 2131.020 1596.390 ;
        RECT 2308.020 1596.380 2311.020 1596.390 ;
        RECT 2488.020 1596.380 2491.020 1596.390 ;
        RECT 2668.020 1596.380 2671.020 1596.390 ;
        RECT 2848.020 1596.380 2851.020 1596.390 ;
        RECT 2958.800 1596.380 2961.800 1596.390 ;
        RECT -42.180 1593.380 2961.800 1596.380 ;
        RECT -42.180 1593.370 -39.180 1593.380 ;
        RECT 148.020 1593.370 151.020 1593.380 ;
        RECT 328.020 1593.370 331.020 1593.380 ;
        RECT 508.020 1593.370 511.020 1593.380 ;
        RECT 688.020 1593.370 691.020 1593.380 ;
        RECT 868.020 1593.370 871.020 1593.380 ;
        RECT 1048.020 1593.370 1051.020 1593.380 ;
        RECT 1228.020 1593.370 1231.020 1593.380 ;
        RECT 1408.020 1593.370 1411.020 1593.380 ;
        RECT 1588.020 1593.370 1591.020 1593.380 ;
        RECT 1768.020 1593.370 1771.020 1593.380 ;
        RECT 1948.020 1593.370 1951.020 1593.380 ;
        RECT 2128.020 1593.370 2131.020 1593.380 ;
        RECT 2308.020 1593.370 2311.020 1593.380 ;
        RECT 2488.020 1593.370 2491.020 1593.380 ;
        RECT 2668.020 1593.370 2671.020 1593.380 ;
        RECT 2848.020 1593.370 2851.020 1593.380 ;
        RECT 2958.800 1593.370 2961.800 1593.380 ;
        RECT -42.180 1416.380 -39.180 1416.390 ;
        RECT 148.020 1416.380 151.020 1416.390 ;
        RECT 328.020 1416.380 331.020 1416.390 ;
        RECT 508.020 1416.380 511.020 1416.390 ;
        RECT 688.020 1416.380 691.020 1416.390 ;
        RECT 868.020 1416.380 871.020 1416.390 ;
        RECT 1048.020 1416.380 1051.020 1416.390 ;
        RECT 1228.020 1416.380 1231.020 1416.390 ;
        RECT 1408.020 1416.380 1411.020 1416.390 ;
        RECT 1588.020 1416.380 1591.020 1416.390 ;
        RECT 1768.020 1416.380 1771.020 1416.390 ;
        RECT 1948.020 1416.380 1951.020 1416.390 ;
        RECT 2128.020 1416.380 2131.020 1416.390 ;
        RECT 2308.020 1416.380 2311.020 1416.390 ;
        RECT 2488.020 1416.380 2491.020 1416.390 ;
        RECT 2668.020 1416.380 2671.020 1416.390 ;
        RECT 2848.020 1416.380 2851.020 1416.390 ;
        RECT 2958.800 1416.380 2961.800 1416.390 ;
        RECT -42.180 1413.380 2961.800 1416.380 ;
        RECT -42.180 1413.370 -39.180 1413.380 ;
        RECT 148.020 1413.370 151.020 1413.380 ;
        RECT 328.020 1413.370 331.020 1413.380 ;
        RECT 508.020 1413.370 511.020 1413.380 ;
        RECT 688.020 1413.370 691.020 1413.380 ;
        RECT 868.020 1413.370 871.020 1413.380 ;
        RECT 1048.020 1413.370 1051.020 1413.380 ;
        RECT 1228.020 1413.370 1231.020 1413.380 ;
        RECT 1408.020 1413.370 1411.020 1413.380 ;
        RECT 1588.020 1413.370 1591.020 1413.380 ;
        RECT 1768.020 1413.370 1771.020 1413.380 ;
        RECT 1948.020 1413.370 1951.020 1413.380 ;
        RECT 2128.020 1413.370 2131.020 1413.380 ;
        RECT 2308.020 1413.370 2311.020 1413.380 ;
        RECT 2488.020 1413.370 2491.020 1413.380 ;
        RECT 2668.020 1413.370 2671.020 1413.380 ;
        RECT 2848.020 1413.370 2851.020 1413.380 ;
        RECT 2958.800 1413.370 2961.800 1413.380 ;
        RECT -42.180 1236.380 -39.180 1236.390 ;
        RECT 148.020 1236.380 151.020 1236.390 ;
        RECT 328.020 1236.380 331.020 1236.390 ;
        RECT 508.020 1236.380 511.020 1236.390 ;
        RECT 688.020 1236.380 691.020 1236.390 ;
        RECT 868.020 1236.380 871.020 1236.390 ;
        RECT 1048.020 1236.380 1051.020 1236.390 ;
        RECT 1228.020 1236.380 1231.020 1236.390 ;
        RECT 1408.020 1236.380 1411.020 1236.390 ;
        RECT 1588.020 1236.380 1591.020 1236.390 ;
        RECT 1768.020 1236.380 1771.020 1236.390 ;
        RECT 1948.020 1236.380 1951.020 1236.390 ;
        RECT 2128.020 1236.380 2131.020 1236.390 ;
        RECT 2308.020 1236.380 2311.020 1236.390 ;
        RECT 2488.020 1236.380 2491.020 1236.390 ;
        RECT 2668.020 1236.380 2671.020 1236.390 ;
        RECT 2848.020 1236.380 2851.020 1236.390 ;
        RECT 2958.800 1236.380 2961.800 1236.390 ;
        RECT -42.180 1233.380 2961.800 1236.380 ;
        RECT -42.180 1233.370 -39.180 1233.380 ;
        RECT 148.020 1233.370 151.020 1233.380 ;
        RECT 328.020 1233.370 331.020 1233.380 ;
        RECT 508.020 1233.370 511.020 1233.380 ;
        RECT 688.020 1233.370 691.020 1233.380 ;
        RECT 868.020 1233.370 871.020 1233.380 ;
        RECT 1048.020 1233.370 1051.020 1233.380 ;
        RECT 1228.020 1233.370 1231.020 1233.380 ;
        RECT 1408.020 1233.370 1411.020 1233.380 ;
        RECT 1588.020 1233.370 1591.020 1233.380 ;
        RECT 1768.020 1233.370 1771.020 1233.380 ;
        RECT 1948.020 1233.370 1951.020 1233.380 ;
        RECT 2128.020 1233.370 2131.020 1233.380 ;
        RECT 2308.020 1233.370 2311.020 1233.380 ;
        RECT 2488.020 1233.370 2491.020 1233.380 ;
        RECT 2668.020 1233.370 2671.020 1233.380 ;
        RECT 2848.020 1233.370 2851.020 1233.380 ;
        RECT 2958.800 1233.370 2961.800 1233.380 ;
        RECT -42.180 1056.380 -39.180 1056.390 ;
        RECT 148.020 1056.380 151.020 1056.390 ;
        RECT 328.020 1056.380 331.020 1056.390 ;
        RECT 508.020 1056.380 511.020 1056.390 ;
        RECT 688.020 1056.380 691.020 1056.390 ;
        RECT 868.020 1056.380 871.020 1056.390 ;
        RECT 1048.020 1056.380 1051.020 1056.390 ;
        RECT 1228.020 1056.380 1231.020 1056.390 ;
        RECT 1408.020 1056.380 1411.020 1056.390 ;
        RECT 1588.020 1056.380 1591.020 1056.390 ;
        RECT 1768.020 1056.380 1771.020 1056.390 ;
        RECT 1948.020 1056.380 1951.020 1056.390 ;
        RECT 2128.020 1056.380 2131.020 1056.390 ;
        RECT 2308.020 1056.380 2311.020 1056.390 ;
        RECT 2488.020 1056.380 2491.020 1056.390 ;
        RECT 2668.020 1056.380 2671.020 1056.390 ;
        RECT 2848.020 1056.380 2851.020 1056.390 ;
        RECT 2958.800 1056.380 2961.800 1056.390 ;
        RECT -42.180 1053.380 2961.800 1056.380 ;
        RECT -42.180 1053.370 -39.180 1053.380 ;
        RECT 148.020 1053.370 151.020 1053.380 ;
        RECT 328.020 1053.370 331.020 1053.380 ;
        RECT 508.020 1053.370 511.020 1053.380 ;
        RECT 688.020 1053.370 691.020 1053.380 ;
        RECT 868.020 1053.370 871.020 1053.380 ;
        RECT 1048.020 1053.370 1051.020 1053.380 ;
        RECT 1228.020 1053.370 1231.020 1053.380 ;
        RECT 1408.020 1053.370 1411.020 1053.380 ;
        RECT 1588.020 1053.370 1591.020 1053.380 ;
        RECT 1768.020 1053.370 1771.020 1053.380 ;
        RECT 1948.020 1053.370 1951.020 1053.380 ;
        RECT 2128.020 1053.370 2131.020 1053.380 ;
        RECT 2308.020 1053.370 2311.020 1053.380 ;
        RECT 2488.020 1053.370 2491.020 1053.380 ;
        RECT 2668.020 1053.370 2671.020 1053.380 ;
        RECT 2848.020 1053.370 2851.020 1053.380 ;
        RECT 2958.800 1053.370 2961.800 1053.380 ;
        RECT -42.180 876.380 -39.180 876.390 ;
        RECT 148.020 876.380 151.020 876.390 ;
        RECT 328.020 876.380 331.020 876.390 ;
        RECT 508.020 876.380 511.020 876.390 ;
        RECT 688.020 876.380 691.020 876.390 ;
        RECT 868.020 876.380 871.020 876.390 ;
        RECT 1048.020 876.380 1051.020 876.390 ;
        RECT 1228.020 876.380 1231.020 876.390 ;
        RECT 1408.020 876.380 1411.020 876.390 ;
        RECT 1588.020 876.380 1591.020 876.390 ;
        RECT 1768.020 876.380 1771.020 876.390 ;
        RECT 1948.020 876.380 1951.020 876.390 ;
        RECT 2128.020 876.380 2131.020 876.390 ;
        RECT 2308.020 876.380 2311.020 876.390 ;
        RECT 2488.020 876.380 2491.020 876.390 ;
        RECT 2668.020 876.380 2671.020 876.390 ;
        RECT 2848.020 876.380 2851.020 876.390 ;
        RECT 2958.800 876.380 2961.800 876.390 ;
        RECT -42.180 873.380 2961.800 876.380 ;
        RECT -42.180 873.370 -39.180 873.380 ;
        RECT 148.020 873.370 151.020 873.380 ;
        RECT 328.020 873.370 331.020 873.380 ;
        RECT 508.020 873.370 511.020 873.380 ;
        RECT 688.020 873.370 691.020 873.380 ;
        RECT 868.020 873.370 871.020 873.380 ;
        RECT 1048.020 873.370 1051.020 873.380 ;
        RECT 1228.020 873.370 1231.020 873.380 ;
        RECT 1408.020 873.370 1411.020 873.380 ;
        RECT 1588.020 873.370 1591.020 873.380 ;
        RECT 1768.020 873.370 1771.020 873.380 ;
        RECT 1948.020 873.370 1951.020 873.380 ;
        RECT 2128.020 873.370 2131.020 873.380 ;
        RECT 2308.020 873.370 2311.020 873.380 ;
        RECT 2488.020 873.370 2491.020 873.380 ;
        RECT 2668.020 873.370 2671.020 873.380 ;
        RECT 2848.020 873.370 2851.020 873.380 ;
        RECT 2958.800 873.370 2961.800 873.380 ;
        RECT -42.180 696.380 -39.180 696.390 ;
        RECT 148.020 696.380 151.020 696.390 ;
        RECT 328.020 696.380 331.020 696.390 ;
        RECT 508.020 696.380 511.020 696.390 ;
        RECT 688.020 696.380 691.020 696.390 ;
        RECT 868.020 696.380 871.020 696.390 ;
        RECT 1048.020 696.380 1051.020 696.390 ;
        RECT 1228.020 696.380 1231.020 696.390 ;
        RECT 1408.020 696.380 1411.020 696.390 ;
        RECT 1588.020 696.380 1591.020 696.390 ;
        RECT 1768.020 696.380 1771.020 696.390 ;
        RECT 1948.020 696.380 1951.020 696.390 ;
        RECT 2128.020 696.380 2131.020 696.390 ;
        RECT 2308.020 696.380 2311.020 696.390 ;
        RECT 2488.020 696.380 2491.020 696.390 ;
        RECT 2668.020 696.380 2671.020 696.390 ;
        RECT 2848.020 696.380 2851.020 696.390 ;
        RECT 2958.800 696.380 2961.800 696.390 ;
        RECT -42.180 693.380 2961.800 696.380 ;
        RECT -42.180 693.370 -39.180 693.380 ;
        RECT 148.020 693.370 151.020 693.380 ;
        RECT 328.020 693.370 331.020 693.380 ;
        RECT 508.020 693.370 511.020 693.380 ;
        RECT 688.020 693.370 691.020 693.380 ;
        RECT 868.020 693.370 871.020 693.380 ;
        RECT 1048.020 693.370 1051.020 693.380 ;
        RECT 1228.020 693.370 1231.020 693.380 ;
        RECT 1408.020 693.370 1411.020 693.380 ;
        RECT 1588.020 693.370 1591.020 693.380 ;
        RECT 1768.020 693.370 1771.020 693.380 ;
        RECT 1948.020 693.370 1951.020 693.380 ;
        RECT 2128.020 693.370 2131.020 693.380 ;
        RECT 2308.020 693.370 2311.020 693.380 ;
        RECT 2488.020 693.370 2491.020 693.380 ;
        RECT 2668.020 693.370 2671.020 693.380 ;
        RECT 2848.020 693.370 2851.020 693.380 ;
        RECT 2958.800 693.370 2961.800 693.380 ;
        RECT -42.180 516.380 -39.180 516.390 ;
        RECT 148.020 516.380 151.020 516.390 ;
        RECT 328.020 516.380 331.020 516.390 ;
        RECT 508.020 516.380 511.020 516.390 ;
        RECT 688.020 516.380 691.020 516.390 ;
        RECT 868.020 516.380 871.020 516.390 ;
        RECT 1048.020 516.380 1051.020 516.390 ;
        RECT 1228.020 516.380 1231.020 516.390 ;
        RECT 1408.020 516.380 1411.020 516.390 ;
        RECT 1588.020 516.380 1591.020 516.390 ;
        RECT 1768.020 516.380 1771.020 516.390 ;
        RECT 1948.020 516.380 1951.020 516.390 ;
        RECT 2128.020 516.380 2131.020 516.390 ;
        RECT 2308.020 516.380 2311.020 516.390 ;
        RECT 2488.020 516.380 2491.020 516.390 ;
        RECT 2668.020 516.380 2671.020 516.390 ;
        RECT 2848.020 516.380 2851.020 516.390 ;
        RECT 2958.800 516.380 2961.800 516.390 ;
        RECT -42.180 513.380 2961.800 516.380 ;
        RECT -42.180 513.370 -39.180 513.380 ;
        RECT 148.020 513.370 151.020 513.380 ;
        RECT 328.020 513.370 331.020 513.380 ;
        RECT 508.020 513.370 511.020 513.380 ;
        RECT 688.020 513.370 691.020 513.380 ;
        RECT 868.020 513.370 871.020 513.380 ;
        RECT 1048.020 513.370 1051.020 513.380 ;
        RECT 1228.020 513.370 1231.020 513.380 ;
        RECT 1408.020 513.370 1411.020 513.380 ;
        RECT 1588.020 513.370 1591.020 513.380 ;
        RECT 1768.020 513.370 1771.020 513.380 ;
        RECT 1948.020 513.370 1951.020 513.380 ;
        RECT 2128.020 513.370 2131.020 513.380 ;
        RECT 2308.020 513.370 2311.020 513.380 ;
        RECT 2488.020 513.370 2491.020 513.380 ;
        RECT 2668.020 513.370 2671.020 513.380 ;
        RECT 2848.020 513.370 2851.020 513.380 ;
        RECT 2958.800 513.370 2961.800 513.380 ;
        RECT -42.180 336.380 -39.180 336.390 ;
        RECT 148.020 336.380 151.020 336.390 ;
        RECT 328.020 336.380 331.020 336.390 ;
        RECT 508.020 336.380 511.020 336.390 ;
        RECT 688.020 336.380 691.020 336.390 ;
        RECT 868.020 336.380 871.020 336.390 ;
        RECT 1048.020 336.380 1051.020 336.390 ;
        RECT 1228.020 336.380 1231.020 336.390 ;
        RECT 1408.020 336.380 1411.020 336.390 ;
        RECT 1588.020 336.380 1591.020 336.390 ;
        RECT 1768.020 336.380 1771.020 336.390 ;
        RECT 1948.020 336.380 1951.020 336.390 ;
        RECT 2128.020 336.380 2131.020 336.390 ;
        RECT 2308.020 336.380 2311.020 336.390 ;
        RECT 2488.020 336.380 2491.020 336.390 ;
        RECT 2668.020 336.380 2671.020 336.390 ;
        RECT 2848.020 336.380 2851.020 336.390 ;
        RECT 2958.800 336.380 2961.800 336.390 ;
        RECT -42.180 333.380 2961.800 336.380 ;
        RECT -42.180 333.370 -39.180 333.380 ;
        RECT 148.020 333.370 151.020 333.380 ;
        RECT 328.020 333.370 331.020 333.380 ;
        RECT 508.020 333.370 511.020 333.380 ;
        RECT 688.020 333.370 691.020 333.380 ;
        RECT 868.020 333.370 871.020 333.380 ;
        RECT 1048.020 333.370 1051.020 333.380 ;
        RECT 1228.020 333.370 1231.020 333.380 ;
        RECT 1408.020 333.370 1411.020 333.380 ;
        RECT 1588.020 333.370 1591.020 333.380 ;
        RECT 1768.020 333.370 1771.020 333.380 ;
        RECT 1948.020 333.370 1951.020 333.380 ;
        RECT 2128.020 333.370 2131.020 333.380 ;
        RECT 2308.020 333.370 2311.020 333.380 ;
        RECT 2488.020 333.370 2491.020 333.380 ;
        RECT 2668.020 333.370 2671.020 333.380 ;
        RECT 2848.020 333.370 2851.020 333.380 ;
        RECT 2958.800 333.370 2961.800 333.380 ;
        RECT -42.180 156.380 -39.180 156.390 ;
        RECT 148.020 156.380 151.020 156.390 ;
        RECT 328.020 156.380 331.020 156.390 ;
        RECT 508.020 156.380 511.020 156.390 ;
        RECT 688.020 156.380 691.020 156.390 ;
        RECT 868.020 156.380 871.020 156.390 ;
        RECT 1048.020 156.380 1051.020 156.390 ;
        RECT 1228.020 156.380 1231.020 156.390 ;
        RECT 1408.020 156.380 1411.020 156.390 ;
        RECT 1588.020 156.380 1591.020 156.390 ;
        RECT 1768.020 156.380 1771.020 156.390 ;
        RECT 1948.020 156.380 1951.020 156.390 ;
        RECT 2128.020 156.380 2131.020 156.390 ;
        RECT 2308.020 156.380 2311.020 156.390 ;
        RECT 2488.020 156.380 2491.020 156.390 ;
        RECT 2668.020 156.380 2671.020 156.390 ;
        RECT 2848.020 156.380 2851.020 156.390 ;
        RECT 2958.800 156.380 2961.800 156.390 ;
        RECT -42.180 153.380 2961.800 156.380 ;
        RECT -42.180 153.370 -39.180 153.380 ;
        RECT 148.020 153.370 151.020 153.380 ;
        RECT 328.020 153.370 331.020 153.380 ;
        RECT 508.020 153.370 511.020 153.380 ;
        RECT 688.020 153.370 691.020 153.380 ;
        RECT 868.020 153.370 871.020 153.380 ;
        RECT 1048.020 153.370 1051.020 153.380 ;
        RECT 1228.020 153.370 1231.020 153.380 ;
        RECT 1408.020 153.370 1411.020 153.380 ;
        RECT 1588.020 153.370 1591.020 153.380 ;
        RECT 1768.020 153.370 1771.020 153.380 ;
        RECT 1948.020 153.370 1951.020 153.380 ;
        RECT 2128.020 153.370 2131.020 153.380 ;
        RECT 2308.020 153.370 2311.020 153.380 ;
        RECT 2488.020 153.370 2491.020 153.380 ;
        RECT 2668.020 153.370 2671.020 153.380 ;
        RECT 2848.020 153.370 2851.020 153.380 ;
        RECT 2958.800 153.370 2961.800 153.380 ;
        RECT -42.180 -33.820 -39.180 -33.810 ;
        RECT 148.020 -33.820 151.020 -33.810 ;
        RECT 328.020 -33.820 331.020 -33.810 ;
        RECT 508.020 -33.820 511.020 -33.810 ;
        RECT 688.020 -33.820 691.020 -33.810 ;
        RECT 868.020 -33.820 871.020 -33.810 ;
        RECT 1048.020 -33.820 1051.020 -33.810 ;
        RECT 1228.020 -33.820 1231.020 -33.810 ;
        RECT 1408.020 -33.820 1411.020 -33.810 ;
        RECT 1588.020 -33.820 1591.020 -33.810 ;
        RECT 1768.020 -33.820 1771.020 -33.810 ;
        RECT 1948.020 -33.820 1951.020 -33.810 ;
        RECT 2128.020 -33.820 2131.020 -33.810 ;
        RECT 2308.020 -33.820 2311.020 -33.810 ;
        RECT 2488.020 -33.820 2491.020 -33.810 ;
        RECT 2668.020 -33.820 2671.020 -33.810 ;
        RECT 2848.020 -33.820 2851.020 -33.810 ;
        RECT 2958.800 -33.820 2961.800 -33.810 ;
        RECT -42.180 -36.820 2961.800 -33.820 ;
        RECT -42.180 -36.830 -39.180 -36.820 ;
        RECT 148.020 -36.830 151.020 -36.820 ;
        RECT 328.020 -36.830 331.020 -36.820 ;
        RECT 508.020 -36.830 511.020 -36.820 ;
        RECT 688.020 -36.830 691.020 -36.820 ;
        RECT 868.020 -36.830 871.020 -36.820 ;
        RECT 1048.020 -36.830 1051.020 -36.820 ;
        RECT 1228.020 -36.830 1231.020 -36.820 ;
        RECT 1408.020 -36.830 1411.020 -36.820 ;
        RECT 1588.020 -36.830 1591.020 -36.820 ;
        RECT 1768.020 -36.830 1771.020 -36.820 ;
        RECT 1948.020 -36.830 1951.020 -36.820 ;
        RECT 2128.020 -36.830 2131.020 -36.820 ;
        RECT 2308.020 -36.830 2311.020 -36.820 ;
        RECT 2488.020 -36.830 2491.020 -36.820 ;
        RECT 2668.020 -36.830 2671.020 -36.820 ;
        RECT 2848.020 -36.830 2851.020 -36.820 ;
        RECT 2958.800 -36.830 2961.800 -36.820 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 1154.070 1710.795 2642.630 3187.925 ;
      LAYER met1 ;
        RECT 1150.000 1704.460 2647.160 3188.080 ;
      LAYER met2 ;
        RECT 1150.030 3195.720 1154.800 3196.000 ;
        RECT 1155.640 3195.720 1167.680 3196.000 ;
        RECT 1168.520 3195.720 1181.020 3196.000 ;
        RECT 1181.860 3195.720 1193.900 3196.000 ;
        RECT 1194.740 3195.720 1207.240 3196.000 ;
        RECT 1208.080 3195.720 1220.580 3196.000 ;
        RECT 1221.420 3195.720 1233.460 3196.000 ;
        RECT 1234.300 3195.720 1246.800 3196.000 ;
        RECT 1247.640 3195.720 1259.680 3196.000 ;
        RECT 1260.520 3195.720 1273.020 3196.000 ;
        RECT 1273.860 3195.720 1286.360 3196.000 ;
        RECT 1287.200 3195.720 1299.240 3196.000 ;
        RECT 1300.080 3195.720 1312.580 3196.000 ;
        RECT 1313.420 3195.720 1325.460 3196.000 ;
        RECT 1326.300 3195.720 1338.800 3196.000 ;
        RECT 1339.640 3195.720 1352.140 3196.000 ;
        RECT 1352.980 3195.720 1365.020 3196.000 ;
        RECT 1365.860 3195.720 1378.360 3196.000 ;
        RECT 1379.200 3195.720 1391.240 3196.000 ;
        RECT 1392.080 3195.720 1404.580 3196.000 ;
        RECT 1405.420 3195.720 1417.920 3196.000 ;
        RECT 1418.760 3195.720 1430.800 3196.000 ;
        RECT 1431.640 3195.720 1444.140 3196.000 ;
        RECT 1444.980 3195.720 1457.020 3196.000 ;
        RECT 1457.860 3195.720 1470.360 3196.000 ;
        RECT 1471.200 3195.720 1483.700 3196.000 ;
        RECT 1484.540 3195.720 1496.580 3196.000 ;
        RECT 1497.420 3195.720 1509.920 3196.000 ;
        RECT 1510.760 3195.720 1522.800 3196.000 ;
        RECT 1523.640 3195.720 1536.140 3196.000 ;
        RECT 1536.980 3195.720 1549.480 3196.000 ;
        RECT 1550.320 3195.720 1562.360 3196.000 ;
        RECT 1563.200 3195.720 1575.700 3196.000 ;
        RECT 1576.540 3195.720 1588.580 3196.000 ;
        RECT 1589.420 3195.720 1601.920 3196.000 ;
        RECT 1602.760 3195.720 1615.260 3196.000 ;
        RECT 1616.100 3195.720 1628.140 3196.000 ;
        RECT 1628.980 3195.720 1641.480 3196.000 ;
        RECT 1642.320 3195.720 1654.820 3196.000 ;
        RECT 1655.660 3195.720 1667.700 3196.000 ;
        RECT 1668.540 3195.720 1681.040 3196.000 ;
        RECT 1681.880 3195.720 1693.920 3196.000 ;
        RECT 1694.760 3195.720 1707.260 3196.000 ;
        RECT 1708.100 3195.720 1720.600 3196.000 ;
        RECT 1721.440 3195.720 1733.480 3196.000 ;
        RECT 1734.320 3195.720 1746.820 3196.000 ;
        RECT 1747.660 3195.720 1759.700 3196.000 ;
        RECT 1760.540 3195.720 1773.040 3196.000 ;
        RECT 1773.880 3195.720 1786.380 3196.000 ;
        RECT 1787.220 3195.720 1799.260 3196.000 ;
        RECT 1800.100 3195.720 1812.600 3196.000 ;
        RECT 1813.440 3195.720 1825.480 3196.000 ;
        RECT 1826.320 3195.720 1838.820 3196.000 ;
        RECT 1839.660 3195.720 1852.160 3196.000 ;
        RECT 1853.000 3195.720 1865.040 3196.000 ;
        RECT 1865.880 3195.720 1878.380 3196.000 ;
        RECT 1879.220 3195.720 1891.260 3196.000 ;
        RECT 1892.100 3195.720 1904.600 3196.000 ;
        RECT 1905.440 3195.720 1917.940 3196.000 ;
        RECT 1918.780 3195.720 1930.820 3196.000 ;
        RECT 1931.660 3195.720 1944.160 3196.000 ;
        RECT 1945.000 3195.720 1957.040 3196.000 ;
        RECT 1957.880 3195.720 1970.380 3196.000 ;
        RECT 1971.220 3195.720 1983.720 3196.000 ;
        RECT 1984.560 3195.720 1996.600 3196.000 ;
        RECT 1997.440 3195.720 2009.940 3196.000 ;
        RECT 2010.780 3195.720 2022.820 3196.000 ;
        RECT 2023.660 3195.720 2036.160 3196.000 ;
        RECT 2037.000 3195.720 2049.500 3196.000 ;
        RECT 2050.340 3195.720 2062.380 3196.000 ;
        RECT 2063.220 3195.720 2075.720 3196.000 ;
        RECT 2076.560 3195.720 2088.600 3196.000 ;
        RECT 2089.440 3195.720 2101.940 3196.000 ;
        RECT 2102.780 3195.720 2115.280 3196.000 ;
        RECT 2116.120 3195.720 2128.160 3196.000 ;
        RECT 2129.000 3195.720 2141.500 3196.000 ;
        RECT 2142.340 3195.720 2154.840 3196.000 ;
        RECT 2155.680 3195.720 2167.720 3196.000 ;
        RECT 2168.560 3195.720 2181.060 3196.000 ;
        RECT 2181.900 3195.720 2193.940 3196.000 ;
        RECT 2194.780 3195.720 2207.280 3196.000 ;
        RECT 2208.120 3195.720 2220.620 3196.000 ;
        RECT 2221.460 3195.720 2233.500 3196.000 ;
        RECT 2234.340 3195.720 2246.840 3196.000 ;
        RECT 2247.680 3195.720 2259.720 3196.000 ;
        RECT 2260.560 3195.720 2273.060 3196.000 ;
        RECT 2273.900 3195.720 2286.400 3196.000 ;
        RECT 2287.240 3195.720 2299.280 3196.000 ;
        RECT 2300.120 3195.720 2312.620 3196.000 ;
        RECT 2313.460 3195.720 2325.500 3196.000 ;
        RECT 2326.340 3195.720 2338.840 3196.000 ;
        RECT 2339.680 3195.720 2352.180 3196.000 ;
        RECT 2353.020 3195.720 2365.060 3196.000 ;
        RECT 2365.900 3195.720 2378.400 3196.000 ;
        RECT 2379.240 3195.720 2391.280 3196.000 ;
        RECT 2392.120 3195.720 2404.620 3196.000 ;
        RECT 2405.460 3195.720 2417.960 3196.000 ;
        RECT 2418.800 3195.720 2430.840 3196.000 ;
        RECT 2431.680 3195.720 2444.180 3196.000 ;
        RECT 2445.020 3195.720 2457.060 3196.000 ;
        RECT 2457.900 3195.720 2470.400 3196.000 ;
        RECT 2471.240 3195.720 2483.740 3196.000 ;
        RECT 2484.580 3195.720 2496.620 3196.000 ;
        RECT 2497.460 3195.720 2509.960 3196.000 ;
        RECT 2510.800 3195.720 2522.840 3196.000 ;
        RECT 2523.680 3195.720 2536.180 3196.000 ;
        RECT 2537.020 3195.720 2549.520 3196.000 ;
        RECT 2550.360 3195.720 2562.400 3196.000 ;
        RECT 2563.240 3195.720 2575.740 3196.000 ;
        RECT 2576.580 3195.720 2588.620 3196.000 ;
        RECT 2589.460 3195.720 2601.960 3196.000 ;
        RECT 2602.800 3195.720 2615.300 3196.000 ;
        RECT 2616.140 3195.720 2628.180 3196.000 ;
        RECT 2629.020 3195.720 2641.520 3196.000 ;
        RECT 2642.360 3195.720 2647.130 3196.000 ;
        RECT 1150.030 1704.280 2647.130 3195.720 ;
        RECT 1150.580 1704.000 1152.500 1704.280 ;
        RECT 1153.340 1704.000 1155.720 1704.280 ;
        RECT 1156.560 1704.000 1158.480 1704.280 ;
        RECT 1159.320 1704.000 1161.700 1704.280 ;
        RECT 1162.540 1704.000 1164.920 1704.280 ;
        RECT 1165.760 1704.000 1167.680 1704.280 ;
        RECT 1168.520 1704.000 1170.900 1704.280 ;
        RECT 1171.740 1704.000 1174.120 1704.280 ;
        RECT 1174.960 1704.000 1176.880 1704.280 ;
        RECT 1177.720 1704.000 1180.100 1704.280 ;
        RECT 1180.940 1704.000 1183.320 1704.280 ;
        RECT 1184.160 1704.000 1186.080 1704.280 ;
        RECT 1186.920 1704.000 1189.300 1704.280 ;
        RECT 1190.140 1704.000 1192.520 1704.280 ;
        RECT 1193.360 1704.000 1195.280 1704.280 ;
        RECT 1196.120 1704.000 1198.500 1704.280 ;
        RECT 1199.340 1704.000 1201.720 1704.280 ;
        RECT 1202.560 1704.000 1204.480 1704.280 ;
        RECT 1205.320 1704.000 1207.700 1704.280 ;
        RECT 1208.540 1704.000 1210.920 1704.280 ;
        RECT 1211.760 1704.000 1213.680 1704.280 ;
        RECT 1214.520 1704.000 1216.900 1704.280 ;
        RECT 1217.740 1704.000 1220.120 1704.280 ;
        RECT 1220.960 1704.000 1222.880 1704.280 ;
        RECT 1223.720 1704.000 1226.100 1704.280 ;
        RECT 1226.940 1704.000 1229.320 1704.280 ;
        RECT 1230.160 1704.000 1232.080 1704.280 ;
        RECT 1232.920 1704.000 1235.300 1704.280 ;
        RECT 1236.140 1704.000 1238.060 1704.280 ;
        RECT 1238.900 1704.000 1241.280 1704.280 ;
        RECT 1242.120 1704.000 1244.500 1704.280 ;
        RECT 1245.340 1704.000 1247.260 1704.280 ;
        RECT 1248.100 1704.000 1250.480 1704.280 ;
        RECT 1251.320 1704.000 1253.700 1704.280 ;
        RECT 1254.540 1704.000 1256.460 1704.280 ;
        RECT 1257.300 1704.000 1259.680 1704.280 ;
        RECT 1260.520 1704.000 1262.900 1704.280 ;
        RECT 1263.740 1704.000 1265.660 1704.280 ;
        RECT 1266.500 1704.000 1268.880 1704.280 ;
        RECT 1269.720 1704.000 1272.100 1704.280 ;
        RECT 1272.940 1704.000 1274.860 1704.280 ;
        RECT 1275.700 1704.000 1278.080 1704.280 ;
        RECT 1278.920 1704.000 1281.300 1704.280 ;
        RECT 1282.140 1704.000 1284.060 1704.280 ;
        RECT 1284.900 1704.000 1287.280 1704.280 ;
        RECT 1288.120 1704.000 1290.500 1704.280 ;
        RECT 1291.340 1704.000 1293.260 1704.280 ;
        RECT 1294.100 1704.000 1296.480 1704.280 ;
        RECT 1297.320 1704.000 1299.700 1704.280 ;
        RECT 1300.540 1704.000 1302.460 1704.280 ;
        RECT 1303.300 1704.000 1305.680 1704.280 ;
        RECT 1306.520 1704.000 1308.900 1704.280 ;
        RECT 1309.740 1704.000 1311.660 1704.280 ;
        RECT 1312.500 1704.000 1314.880 1704.280 ;
        RECT 1315.720 1704.000 1318.100 1704.280 ;
        RECT 1318.940 1704.000 1320.860 1704.280 ;
        RECT 1321.700 1704.000 1324.080 1704.280 ;
        RECT 1324.920 1704.000 1326.840 1704.280 ;
        RECT 1327.680 1704.000 1330.060 1704.280 ;
        RECT 1330.900 1704.000 1333.280 1704.280 ;
        RECT 1334.120 1704.000 1336.040 1704.280 ;
        RECT 1336.880 1704.000 1339.260 1704.280 ;
        RECT 1340.100 1704.000 1342.480 1704.280 ;
        RECT 1343.320 1704.000 1345.240 1704.280 ;
        RECT 1346.080 1704.000 1348.460 1704.280 ;
        RECT 1349.300 1704.000 1351.680 1704.280 ;
        RECT 1352.520 1704.000 1354.440 1704.280 ;
        RECT 1355.280 1704.000 1357.660 1704.280 ;
        RECT 1358.500 1704.000 1360.880 1704.280 ;
        RECT 1361.720 1704.000 1363.640 1704.280 ;
        RECT 1364.480 1704.000 1366.860 1704.280 ;
        RECT 1367.700 1704.000 1370.080 1704.280 ;
        RECT 1370.920 1704.000 1372.840 1704.280 ;
        RECT 1373.680 1704.000 1376.060 1704.280 ;
        RECT 1376.900 1704.000 1379.280 1704.280 ;
        RECT 1380.120 1704.000 1382.040 1704.280 ;
        RECT 1382.880 1704.000 1385.260 1704.280 ;
        RECT 1386.100 1704.000 1388.480 1704.280 ;
        RECT 1389.320 1704.000 1391.240 1704.280 ;
        RECT 1392.080 1704.000 1394.460 1704.280 ;
        RECT 1395.300 1704.000 1397.680 1704.280 ;
        RECT 1398.520 1704.000 1400.440 1704.280 ;
        RECT 1401.280 1704.000 1403.660 1704.280 ;
        RECT 1404.500 1704.000 1406.880 1704.280 ;
        RECT 1407.720 1704.000 1409.640 1704.280 ;
        RECT 1410.480 1704.000 1412.860 1704.280 ;
        RECT 1413.700 1704.000 1415.620 1704.280 ;
        RECT 1416.460 1704.000 1418.840 1704.280 ;
        RECT 1419.680 1704.000 1422.060 1704.280 ;
        RECT 1422.900 1704.000 1424.820 1704.280 ;
        RECT 1425.660 1704.000 1428.040 1704.280 ;
        RECT 1428.880 1704.000 1431.260 1704.280 ;
        RECT 1432.100 1704.000 1434.020 1704.280 ;
        RECT 1434.860 1704.000 1437.240 1704.280 ;
        RECT 1438.080 1704.000 1440.460 1704.280 ;
        RECT 1441.300 1704.000 1443.220 1704.280 ;
        RECT 1444.060 1704.000 1446.440 1704.280 ;
        RECT 1447.280 1704.000 1449.660 1704.280 ;
        RECT 1450.500 1704.000 1452.420 1704.280 ;
        RECT 1453.260 1704.000 1455.640 1704.280 ;
        RECT 1456.480 1704.000 1458.860 1704.280 ;
        RECT 1459.700 1704.000 1461.620 1704.280 ;
        RECT 1462.460 1704.000 1464.840 1704.280 ;
        RECT 1465.680 1704.000 1468.060 1704.280 ;
        RECT 1468.900 1704.000 1470.820 1704.280 ;
        RECT 1471.660 1704.000 1474.040 1704.280 ;
        RECT 1474.880 1704.000 1477.260 1704.280 ;
        RECT 1478.100 1704.000 1480.020 1704.280 ;
        RECT 1480.860 1704.000 1483.240 1704.280 ;
        RECT 1484.080 1704.000 1486.460 1704.280 ;
        RECT 1487.300 1704.000 1489.220 1704.280 ;
        RECT 1490.060 1704.000 1492.440 1704.280 ;
        RECT 1493.280 1704.000 1495.660 1704.280 ;
        RECT 1496.500 1704.000 1498.420 1704.280 ;
        RECT 1499.260 1704.000 1501.640 1704.280 ;
        RECT 1502.480 1704.000 1504.400 1704.280 ;
        RECT 1505.240 1704.000 1507.620 1704.280 ;
        RECT 1508.460 1704.000 1510.840 1704.280 ;
        RECT 1511.680 1704.000 1513.600 1704.280 ;
        RECT 1514.440 1704.000 1516.820 1704.280 ;
        RECT 1517.660 1704.000 1520.040 1704.280 ;
        RECT 1520.880 1704.000 1522.800 1704.280 ;
        RECT 1523.640 1704.000 1526.020 1704.280 ;
        RECT 1526.860 1704.000 1529.240 1704.280 ;
        RECT 1530.080 1704.000 1532.000 1704.280 ;
        RECT 1532.840 1704.000 1535.220 1704.280 ;
        RECT 1536.060 1704.000 1538.440 1704.280 ;
        RECT 1539.280 1704.000 1541.200 1704.280 ;
        RECT 1542.040 1704.000 1544.420 1704.280 ;
        RECT 1545.260 1704.000 1547.640 1704.280 ;
        RECT 1548.480 1704.000 1550.400 1704.280 ;
        RECT 1551.240 1704.000 1553.620 1704.280 ;
        RECT 1554.460 1704.000 1556.840 1704.280 ;
        RECT 1557.680 1704.000 1559.600 1704.280 ;
        RECT 1560.440 1704.000 1562.820 1704.280 ;
        RECT 1563.660 1704.000 1566.040 1704.280 ;
        RECT 1566.880 1704.000 1568.800 1704.280 ;
        RECT 1569.640 1704.000 1572.020 1704.280 ;
        RECT 1572.860 1704.000 1575.240 1704.280 ;
        RECT 1576.080 1704.000 1578.000 1704.280 ;
        RECT 1578.840 1704.000 1581.220 1704.280 ;
        RECT 1582.060 1704.000 1584.440 1704.280 ;
        RECT 1585.280 1704.000 1587.200 1704.280 ;
        RECT 1588.040 1704.000 1590.420 1704.280 ;
        RECT 1591.260 1704.000 1593.180 1704.280 ;
        RECT 1594.020 1704.000 1596.400 1704.280 ;
        RECT 1597.240 1704.000 1599.620 1704.280 ;
        RECT 1600.460 1704.000 1602.380 1704.280 ;
        RECT 1603.220 1704.000 1605.600 1704.280 ;
        RECT 1606.440 1704.000 1608.820 1704.280 ;
        RECT 1609.660 1704.000 1611.580 1704.280 ;
        RECT 1612.420 1704.000 1614.800 1704.280 ;
        RECT 1615.640 1704.000 1618.020 1704.280 ;
        RECT 1618.860 1704.000 1620.780 1704.280 ;
        RECT 1621.620 1704.000 1624.000 1704.280 ;
        RECT 1624.840 1704.000 1627.220 1704.280 ;
        RECT 1628.060 1704.000 1629.980 1704.280 ;
        RECT 1630.820 1704.000 1633.200 1704.280 ;
        RECT 1634.040 1704.000 1636.420 1704.280 ;
        RECT 1637.260 1704.000 1639.180 1704.280 ;
        RECT 1640.020 1704.000 1642.400 1704.280 ;
        RECT 1643.240 1704.000 1645.620 1704.280 ;
        RECT 1646.460 1704.000 1648.380 1704.280 ;
        RECT 1649.220 1704.000 1651.600 1704.280 ;
        RECT 1652.440 1704.000 1654.820 1704.280 ;
        RECT 1655.660 1704.000 1657.580 1704.280 ;
        RECT 1658.420 1704.000 1660.800 1704.280 ;
        RECT 1661.640 1704.000 1664.020 1704.280 ;
        RECT 1664.860 1704.000 1666.780 1704.280 ;
        RECT 1667.620 1704.000 1670.000 1704.280 ;
        RECT 1670.840 1704.000 1673.220 1704.280 ;
        RECT 1674.060 1704.000 1675.980 1704.280 ;
        RECT 1676.820 1704.000 1679.200 1704.280 ;
        RECT 1680.040 1704.000 1681.960 1704.280 ;
        RECT 1682.800 1704.000 1685.180 1704.280 ;
        RECT 1686.020 1704.000 1688.400 1704.280 ;
        RECT 1689.240 1704.000 1691.160 1704.280 ;
        RECT 1692.000 1704.000 1694.380 1704.280 ;
        RECT 1695.220 1704.000 1697.600 1704.280 ;
        RECT 1698.440 1704.000 1700.360 1704.280 ;
        RECT 1701.200 1704.000 1703.580 1704.280 ;
        RECT 1704.420 1704.000 1706.800 1704.280 ;
        RECT 1707.640 1704.000 1709.560 1704.280 ;
        RECT 1710.400 1704.000 1712.780 1704.280 ;
        RECT 1713.620 1704.000 1716.000 1704.280 ;
        RECT 1716.840 1704.000 1718.760 1704.280 ;
        RECT 1719.600 1704.000 1721.980 1704.280 ;
        RECT 1722.820 1704.000 1725.200 1704.280 ;
        RECT 1726.040 1704.000 1727.960 1704.280 ;
        RECT 1728.800 1704.000 1731.180 1704.280 ;
        RECT 1732.020 1704.000 1734.400 1704.280 ;
        RECT 1735.240 1704.000 1737.160 1704.280 ;
        RECT 1738.000 1704.000 1740.380 1704.280 ;
        RECT 1741.220 1704.000 1743.600 1704.280 ;
        RECT 1744.440 1704.000 1746.360 1704.280 ;
        RECT 1747.200 1704.000 1749.580 1704.280 ;
        RECT 1750.420 1704.000 1752.800 1704.280 ;
        RECT 1753.640 1704.000 1755.560 1704.280 ;
        RECT 1756.400 1704.000 1758.780 1704.280 ;
        RECT 1759.620 1704.000 1762.000 1704.280 ;
        RECT 1762.840 1704.000 1764.760 1704.280 ;
        RECT 1765.600 1704.000 1767.980 1704.280 ;
        RECT 1768.820 1704.000 1770.740 1704.280 ;
        RECT 1771.580 1704.000 1773.960 1704.280 ;
        RECT 1774.800 1704.000 1777.180 1704.280 ;
        RECT 1778.020 1704.000 1779.940 1704.280 ;
        RECT 1780.780 1704.000 1783.160 1704.280 ;
        RECT 1784.000 1704.000 1786.380 1704.280 ;
        RECT 1787.220 1704.000 1789.140 1704.280 ;
        RECT 1789.980 1704.000 1792.360 1704.280 ;
        RECT 1793.200 1704.000 1795.580 1704.280 ;
        RECT 1796.420 1704.000 1798.340 1704.280 ;
        RECT 1799.180 1704.000 1801.560 1704.280 ;
        RECT 1802.400 1704.000 1804.780 1704.280 ;
        RECT 1805.620 1704.000 1807.540 1704.280 ;
        RECT 1808.380 1704.000 1810.760 1704.280 ;
        RECT 1811.600 1704.000 1813.980 1704.280 ;
        RECT 1814.820 1704.000 1816.740 1704.280 ;
        RECT 1817.580 1704.000 1819.960 1704.280 ;
        RECT 1820.800 1704.000 1823.180 1704.280 ;
        RECT 1824.020 1704.000 1825.940 1704.280 ;
        RECT 1826.780 1704.000 1829.160 1704.280 ;
        RECT 1830.000 1704.000 1832.380 1704.280 ;
        RECT 1833.220 1704.000 1835.140 1704.280 ;
        RECT 1835.980 1704.000 1838.360 1704.280 ;
        RECT 1839.200 1704.000 1841.580 1704.280 ;
        RECT 1842.420 1704.000 1844.340 1704.280 ;
        RECT 1845.180 1704.000 1847.560 1704.280 ;
        RECT 1848.400 1704.000 1850.780 1704.280 ;
        RECT 1851.620 1704.000 1853.540 1704.280 ;
        RECT 1854.380 1704.000 1856.760 1704.280 ;
        RECT 1857.600 1704.000 1859.520 1704.280 ;
        RECT 1860.360 1704.000 1862.740 1704.280 ;
        RECT 1863.580 1704.000 1865.960 1704.280 ;
        RECT 1866.800 1704.000 1868.720 1704.280 ;
        RECT 1869.560 1704.000 1871.940 1704.280 ;
        RECT 1872.780 1704.000 1875.160 1704.280 ;
        RECT 1876.000 1704.000 1877.920 1704.280 ;
        RECT 1878.760 1704.000 1881.140 1704.280 ;
        RECT 1881.980 1704.000 1884.360 1704.280 ;
        RECT 1885.200 1704.000 1887.120 1704.280 ;
        RECT 1887.960 1704.000 1890.340 1704.280 ;
        RECT 1891.180 1704.000 1893.560 1704.280 ;
        RECT 1894.400 1704.000 1896.320 1704.280 ;
        RECT 1897.160 1704.000 1899.540 1704.280 ;
        RECT 1900.380 1704.000 1902.760 1704.280 ;
        RECT 1903.600 1704.000 1905.520 1704.280 ;
        RECT 1906.360 1704.000 1908.740 1704.280 ;
        RECT 1909.580 1704.000 1911.960 1704.280 ;
        RECT 1912.800 1704.000 1914.720 1704.280 ;
        RECT 1915.560 1704.000 1917.940 1704.280 ;
        RECT 1918.780 1704.000 1921.160 1704.280 ;
        RECT 1922.000 1704.000 1923.920 1704.280 ;
        RECT 1924.760 1704.000 1927.140 1704.280 ;
        RECT 1927.980 1704.000 1930.360 1704.280 ;
        RECT 1931.200 1704.000 1933.120 1704.280 ;
        RECT 1933.960 1704.000 1936.340 1704.280 ;
        RECT 1937.180 1704.000 1939.560 1704.280 ;
        RECT 1940.400 1704.000 1942.320 1704.280 ;
        RECT 1943.160 1704.000 1945.540 1704.280 ;
        RECT 1946.380 1704.000 1948.300 1704.280 ;
        RECT 1949.140 1704.000 1951.520 1704.280 ;
        RECT 1952.360 1704.000 1954.740 1704.280 ;
        RECT 1955.580 1704.000 1957.500 1704.280 ;
        RECT 1958.340 1704.000 1960.720 1704.280 ;
        RECT 1961.560 1704.000 1963.940 1704.280 ;
        RECT 1964.780 1704.000 1966.700 1704.280 ;
        RECT 1967.540 1704.000 1969.920 1704.280 ;
        RECT 1970.760 1704.000 1973.140 1704.280 ;
        RECT 1973.980 1704.000 1975.900 1704.280 ;
        RECT 1976.740 1704.000 1979.120 1704.280 ;
        RECT 1979.960 1704.000 1982.340 1704.280 ;
        RECT 1983.180 1704.000 1985.100 1704.280 ;
        RECT 1985.940 1704.000 1988.320 1704.280 ;
        RECT 1989.160 1704.000 1991.540 1704.280 ;
        RECT 1992.380 1704.000 1994.300 1704.280 ;
        RECT 1995.140 1704.000 1997.520 1704.280 ;
        RECT 1998.360 1704.000 2000.740 1704.280 ;
        RECT 2001.580 1704.000 2003.500 1704.280 ;
        RECT 2004.340 1704.000 2006.720 1704.280 ;
        RECT 2007.560 1704.000 2009.940 1704.280 ;
        RECT 2010.780 1704.000 2012.700 1704.280 ;
        RECT 2013.540 1704.000 2015.920 1704.280 ;
        RECT 2016.760 1704.000 2019.140 1704.280 ;
        RECT 2019.980 1704.000 2021.900 1704.280 ;
        RECT 2022.740 1704.000 2025.120 1704.280 ;
        RECT 2025.960 1704.000 2028.340 1704.280 ;
        RECT 2029.180 1704.000 2031.100 1704.280 ;
        RECT 2031.940 1704.000 2034.320 1704.280 ;
        RECT 2035.160 1704.000 2037.080 1704.280 ;
        RECT 2037.920 1704.000 2040.300 1704.280 ;
        RECT 2041.140 1704.000 2043.520 1704.280 ;
        RECT 2044.360 1704.000 2046.280 1704.280 ;
        RECT 2047.120 1704.000 2049.500 1704.280 ;
        RECT 2050.340 1704.000 2052.720 1704.280 ;
        RECT 2053.560 1704.000 2055.480 1704.280 ;
        RECT 2056.320 1704.000 2058.700 1704.280 ;
        RECT 2059.540 1704.000 2061.920 1704.280 ;
        RECT 2062.760 1704.000 2064.680 1704.280 ;
        RECT 2065.520 1704.000 2067.900 1704.280 ;
        RECT 2068.740 1704.000 2071.120 1704.280 ;
        RECT 2071.960 1704.000 2073.880 1704.280 ;
        RECT 2074.720 1704.000 2077.100 1704.280 ;
        RECT 2077.940 1704.000 2080.320 1704.280 ;
        RECT 2081.160 1704.000 2083.080 1704.280 ;
        RECT 2083.920 1704.000 2086.300 1704.280 ;
        RECT 2087.140 1704.000 2089.520 1704.280 ;
        RECT 2090.360 1704.000 2092.280 1704.280 ;
        RECT 2093.120 1704.000 2095.500 1704.280 ;
        RECT 2096.340 1704.000 2098.720 1704.280 ;
        RECT 2099.560 1704.000 2101.480 1704.280 ;
        RECT 2102.320 1704.000 2104.700 1704.280 ;
        RECT 2105.540 1704.000 2107.920 1704.280 ;
        RECT 2108.760 1704.000 2110.680 1704.280 ;
        RECT 2111.520 1704.000 2113.900 1704.280 ;
        RECT 2114.740 1704.000 2117.120 1704.280 ;
        RECT 2117.960 1704.000 2119.880 1704.280 ;
        RECT 2120.720 1704.000 2123.100 1704.280 ;
        RECT 2123.940 1704.000 2125.860 1704.280 ;
        RECT 2126.700 1704.000 2129.080 1704.280 ;
        RECT 2129.920 1704.000 2132.300 1704.280 ;
        RECT 2133.140 1704.000 2135.060 1704.280 ;
        RECT 2135.900 1704.000 2138.280 1704.280 ;
        RECT 2139.120 1704.000 2141.500 1704.280 ;
        RECT 2142.340 1704.000 2144.260 1704.280 ;
        RECT 2145.100 1704.000 2147.480 1704.280 ;
        RECT 2148.320 1704.000 2150.700 1704.280 ;
        RECT 2151.540 1704.000 2153.460 1704.280 ;
        RECT 2154.300 1704.000 2156.680 1704.280 ;
        RECT 2157.520 1704.000 2159.900 1704.280 ;
        RECT 2160.740 1704.000 2162.660 1704.280 ;
        RECT 2163.500 1704.000 2165.880 1704.280 ;
        RECT 2166.720 1704.000 2169.100 1704.280 ;
        RECT 2169.940 1704.000 2171.860 1704.280 ;
        RECT 2172.700 1704.000 2175.080 1704.280 ;
        RECT 2175.920 1704.000 2178.300 1704.280 ;
        RECT 2179.140 1704.000 2181.060 1704.280 ;
        RECT 2181.900 1704.000 2184.280 1704.280 ;
        RECT 2185.120 1704.000 2187.500 1704.280 ;
        RECT 2188.340 1704.000 2190.260 1704.280 ;
        RECT 2191.100 1704.000 2193.480 1704.280 ;
        RECT 2194.320 1704.000 2196.700 1704.280 ;
        RECT 2197.540 1704.000 2199.460 1704.280 ;
        RECT 2200.300 1704.000 2202.680 1704.280 ;
        RECT 2203.520 1704.000 2205.900 1704.280 ;
        RECT 2206.740 1704.000 2208.660 1704.280 ;
        RECT 2209.500 1704.000 2211.880 1704.280 ;
        RECT 2212.720 1704.000 2214.640 1704.280 ;
        RECT 2215.480 1704.000 2217.860 1704.280 ;
        RECT 2218.700 1704.000 2221.080 1704.280 ;
        RECT 2221.920 1704.000 2223.840 1704.280 ;
        RECT 2224.680 1704.000 2227.060 1704.280 ;
        RECT 2227.900 1704.000 2230.280 1704.280 ;
        RECT 2231.120 1704.000 2233.040 1704.280 ;
        RECT 2233.880 1704.000 2236.260 1704.280 ;
        RECT 2237.100 1704.000 2239.480 1704.280 ;
        RECT 2240.320 1704.000 2242.240 1704.280 ;
        RECT 2243.080 1704.000 2245.460 1704.280 ;
        RECT 2246.300 1704.000 2248.680 1704.280 ;
        RECT 2249.520 1704.000 2251.440 1704.280 ;
        RECT 2252.280 1704.000 2254.660 1704.280 ;
        RECT 2255.500 1704.000 2257.880 1704.280 ;
        RECT 2258.720 1704.000 2260.640 1704.280 ;
        RECT 2261.480 1704.000 2263.860 1704.280 ;
        RECT 2264.700 1704.000 2267.080 1704.280 ;
        RECT 2267.920 1704.000 2269.840 1704.280 ;
        RECT 2270.680 1704.000 2273.060 1704.280 ;
        RECT 2273.900 1704.000 2276.280 1704.280 ;
        RECT 2277.120 1704.000 2279.040 1704.280 ;
        RECT 2279.880 1704.000 2282.260 1704.280 ;
        RECT 2283.100 1704.000 2285.480 1704.280 ;
        RECT 2286.320 1704.000 2288.240 1704.280 ;
        RECT 2289.080 1704.000 2291.460 1704.280 ;
        RECT 2292.300 1704.000 2294.680 1704.280 ;
        RECT 2295.520 1704.000 2297.440 1704.280 ;
        RECT 2298.280 1704.000 2300.660 1704.280 ;
        RECT 2301.500 1704.000 2303.420 1704.280 ;
        RECT 2304.260 1704.000 2306.640 1704.280 ;
        RECT 2307.480 1704.000 2309.860 1704.280 ;
        RECT 2310.700 1704.000 2312.620 1704.280 ;
        RECT 2313.460 1704.000 2315.840 1704.280 ;
        RECT 2316.680 1704.000 2319.060 1704.280 ;
        RECT 2319.900 1704.000 2321.820 1704.280 ;
        RECT 2322.660 1704.000 2325.040 1704.280 ;
        RECT 2325.880 1704.000 2328.260 1704.280 ;
        RECT 2329.100 1704.000 2331.020 1704.280 ;
        RECT 2331.860 1704.000 2334.240 1704.280 ;
        RECT 2335.080 1704.000 2337.460 1704.280 ;
        RECT 2338.300 1704.000 2340.220 1704.280 ;
        RECT 2341.060 1704.000 2343.440 1704.280 ;
        RECT 2344.280 1704.000 2346.660 1704.280 ;
        RECT 2347.500 1704.000 2349.420 1704.280 ;
        RECT 2350.260 1704.000 2352.640 1704.280 ;
        RECT 2353.480 1704.000 2355.860 1704.280 ;
        RECT 2356.700 1704.000 2358.620 1704.280 ;
        RECT 2359.460 1704.000 2361.840 1704.280 ;
        RECT 2362.680 1704.000 2365.060 1704.280 ;
        RECT 2365.900 1704.000 2367.820 1704.280 ;
        RECT 2368.660 1704.000 2371.040 1704.280 ;
        RECT 2371.880 1704.000 2374.260 1704.280 ;
        RECT 2375.100 1704.000 2377.020 1704.280 ;
        RECT 2377.860 1704.000 2380.240 1704.280 ;
        RECT 2381.080 1704.000 2383.460 1704.280 ;
        RECT 2384.300 1704.000 2386.220 1704.280 ;
        RECT 2387.060 1704.000 2389.440 1704.280 ;
        RECT 2390.280 1704.000 2392.200 1704.280 ;
        RECT 2393.040 1704.000 2395.420 1704.280 ;
        RECT 2396.260 1704.000 2398.640 1704.280 ;
        RECT 2399.480 1704.000 2401.400 1704.280 ;
        RECT 2402.240 1704.000 2404.620 1704.280 ;
        RECT 2405.460 1704.000 2407.840 1704.280 ;
        RECT 2408.680 1704.000 2410.600 1704.280 ;
        RECT 2411.440 1704.000 2413.820 1704.280 ;
        RECT 2414.660 1704.000 2417.040 1704.280 ;
        RECT 2417.880 1704.000 2419.800 1704.280 ;
        RECT 2420.640 1704.000 2423.020 1704.280 ;
        RECT 2423.860 1704.000 2426.240 1704.280 ;
        RECT 2427.080 1704.000 2429.000 1704.280 ;
        RECT 2429.840 1704.000 2432.220 1704.280 ;
        RECT 2433.060 1704.000 2435.440 1704.280 ;
        RECT 2436.280 1704.000 2438.200 1704.280 ;
        RECT 2439.040 1704.000 2441.420 1704.280 ;
        RECT 2442.260 1704.000 2444.640 1704.280 ;
        RECT 2445.480 1704.000 2447.400 1704.280 ;
        RECT 2448.240 1704.000 2450.620 1704.280 ;
        RECT 2451.460 1704.000 2453.840 1704.280 ;
        RECT 2454.680 1704.000 2456.600 1704.280 ;
        RECT 2457.440 1704.000 2459.820 1704.280 ;
        RECT 2460.660 1704.000 2463.040 1704.280 ;
        RECT 2463.880 1704.000 2465.800 1704.280 ;
        RECT 2466.640 1704.000 2469.020 1704.280 ;
        RECT 2469.860 1704.000 2472.240 1704.280 ;
        RECT 2473.080 1704.000 2475.000 1704.280 ;
        RECT 2475.840 1704.000 2478.220 1704.280 ;
        RECT 2479.060 1704.000 2480.980 1704.280 ;
        RECT 2481.820 1704.000 2484.200 1704.280 ;
        RECT 2485.040 1704.000 2487.420 1704.280 ;
        RECT 2488.260 1704.000 2490.180 1704.280 ;
        RECT 2491.020 1704.000 2493.400 1704.280 ;
        RECT 2494.240 1704.000 2496.620 1704.280 ;
        RECT 2497.460 1704.000 2499.380 1704.280 ;
        RECT 2500.220 1704.000 2502.600 1704.280 ;
        RECT 2503.440 1704.000 2505.820 1704.280 ;
        RECT 2506.660 1704.000 2508.580 1704.280 ;
        RECT 2509.420 1704.000 2511.800 1704.280 ;
        RECT 2512.640 1704.000 2515.020 1704.280 ;
        RECT 2515.860 1704.000 2517.780 1704.280 ;
        RECT 2518.620 1704.000 2521.000 1704.280 ;
        RECT 2521.840 1704.000 2524.220 1704.280 ;
        RECT 2525.060 1704.000 2526.980 1704.280 ;
        RECT 2527.820 1704.000 2530.200 1704.280 ;
        RECT 2531.040 1704.000 2533.420 1704.280 ;
        RECT 2534.260 1704.000 2536.180 1704.280 ;
        RECT 2537.020 1704.000 2539.400 1704.280 ;
        RECT 2540.240 1704.000 2542.620 1704.280 ;
        RECT 2543.460 1704.000 2545.380 1704.280 ;
        RECT 2546.220 1704.000 2548.600 1704.280 ;
        RECT 2549.440 1704.000 2551.820 1704.280 ;
        RECT 2552.660 1704.000 2554.580 1704.280 ;
        RECT 2555.420 1704.000 2557.800 1704.280 ;
        RECT 2558.640 1704.000 2561.020 1704.280 ;
        RECT 2561.860 1704.000 2563.780 1704.280 ;
        RECT 2564.620 1704.000 2567.000 1704.280 ;
        RECT 2567.840 1704.000 2569.760 1704.280 ;
        RECT 2570.600 1704.000 2572.980 1704.280 ;
        RECT 2573.820 1704.000 2576.200 1704.280 ;
        RECT 2577.040 1704.000 2578.960 1704.280 ;
        RECT 2579.800 1704.000 2582.180 1704.280 ;
        RECT 2583.020 1704.000 2585.400 1704.280 ;
        RECT 2586.240 1704.000 2588.160 1704.280 ;
        RECT 2589.000 1704.000 2591.380 1704.280 ;
        RECT 2592.220 1704.000 2594.600 1704.280 ;
        RECT 2595.440 1704.000 2597.360 1704.280 ;
        RECT 2598.200 1704.000 2600.580 1704.280 ;
        RECT 2601.420 1704.000 2603.800 1704.280 ;
        RECT 2604.640 1704.000 2606.560 1704.280 ;
        RECT 2607.400 1704.000 2609.780 1704.280 ;
        RECT 2610.620 1704.000 2613.000 1704.280 ;
        RECT 2613.840 1704.000 2615.760 1704.280 ;
        RECT 2616.600 1704.000 2618.980 1704.280 ;
        RECT 2619.820 1704.000 2622.200 1704.280 ;
        RECT 2623.040 1704.000 2624.960 1704.280 ;
        RECT 2625.800 1704.000 2628.180 1704.280 ;
        RECT 2629.020 1704.000 2631.400 1704.280 ;
        RECT 2632.240 1704.000 2634.160 1704.280 ;
        RECT 2635.000 1704.000 2637.380 1704.280 ;
        RECT 2638.220 1704.000 2640.600 1704.280 ;
        RECT 2641.440 1704.000 2643.360 1704.280 ;
        RECT 2644.200 1704.000 2646.580 1704.280 ;
      LAYER met3 ;
        RECT 1161.955 1704.255 2633.825 3188.005 ;
      LAYER met4 ;
        RECT 1169.590 1710.640 1171.190 3188.080 ;
        RECT 1246.390 1710.640 1247.990 3188.080 ;
      LAYER met4 ;
        RECT 1323.190 1710.640 1354.020 3188.080 ;
        RECT 1357.020 1710.640 1372.020 3188.080 ;
        RECT 1375.020 1710.640 1390.020 3188.080 ;
        RECT 1393.020 1710.640 1408.020 3188.080 ;
        RECT 1411.020 1710.640 1444.020 3188.080 ;
        RECT 1447.020 1710.640 1462.020 3188.080 ;
        RECT 1465.020 1710.640 1480.020 3188.080 ;
        RECT 1483.020 1710.640 1498.020 3188.080 ;
        RECT 1501.020 1710.640 1534.020 3188.080 ;
        RECT 1537.020 1710.640 1552.020 3188.080 ;
        RECT 1555.020 1710.640 1570.020 3188.080 ;
        RECT 1573.020 1710.640 1588.020 3188.080 ;
        RECT 1591.020 1710.640 1624.020 3188.080 ;
        RECT 1627.020 1710.640 1642.020 3188.080 ;
        RECT 1645.020 1710.640 1660.020 3188.080 ;
        RECT 1663.020 1710.640 1678.020 3188.080 ;
        RECT 1681.020 1710.640 1714.020 3188.080 ;
        RECT 1717.020 1710.640 1732.020 3188.080 ;
        RECT 1735.020 1710.640 1750.020 3188.080 ;
        RECT 1753.020 1710.640 1768.020 3188.080 ;
        RECT 1771.020 1710.640 1804.020 3188.080 ;
        RECT 1807.020 1710.640 1822.020 3188.080 ;
        RECT 1825.020 1710.640 1840.020 3188.080 ;
        RECT 1843.020 1710.640 1858.020 3188.080 ;
        RECT 1861.020 1710.640 1894.020 3188.080 ;
        RECT 1897.020 1710.640 1912.020 3188.080 ;
        RECT 1915.020 1710.640 1930.020 3188.080 ;
        RECT 1933.020 1710.640 1948.020 3188.080 ;
        RECT 1951.020 1710.640 1984.020 3188.080 ;
        RECT 1987.020 1710.640 2002.020 3188.080 ;
        RECT 2005.020 1710.640 2020.020 3188.080 ;
        RECT 2023.020 1710.640 2038.020 3188.080 ;
        RECT 2041.020 1710.640 2074.020 3188.080 ;
        RECT 2077.020 1710.640 2092.020 3188.080 ;
        RECT 2095.020 1710.640 2110.020 3188.080 ;
        RECT 2113.020 1710.640 2128.020 3188.080 ;
        RECT 2131.020 1710.640 2164.020 3188.080 ;
        RECT 2167.020 1710.640 2182.020 3188.080 ;
        RECT 2185.020 1710.640 2200.020 3188.080 ;
        RECT 2203.020 1710.640 2218.020 3188.080 ;
        RECT 2221.020 1710.640 2254.020 3188.080 ;
        RECT 2257.020 1710.640 2272.020 3188.080 ;
        RECT 2275.020 1710.640 2290.020 3188.080 ;
        RECT 2293.020 1710.640 2308.020 3188.080 ;
        RECT 2311.020 1710.640 2344.020 3188.080 ;
        RECT 2347.020 1710.640 2362.020 3188.080 ;
        RECT 2365.020 1710.640 2380.020 3188.080 ;
        RECT 2383.020 1710.640 2398.020 3188.080 ;
        RECT 2401.020 1710.640 2434.020 3188.080 ;
        RECT 2437.020 1710.640 2452.020 3188.080 ;
        RECT 2455.020 1710.640 2470.020 3188.080 ;
        RECT 2473.020 1710.640 2488.020 3188.080 ;
        RECT 2491.020 1710.640 2524.020 3188.080 ;
        RECT 2527.020 1710.640 2542.020 3188.080 ;
        RECT 2545.020 1710.640 2560.020 3188.080 ;
        RECT 2563.020 1710.640 2578.020 3188.080 ;
        RECT 2581.020 1710.640 2614.020 3188.080 ;
        RECT 2617.020 1710.640 2630.390 3188.080 ;
  END
END user_project_wrapper
END LIBRARY

