magic
tech sky130A
magscale 1 2
timestamp 1607890414
<< obsli1 >>
rect 908 2159 218672 217617
<< obsm1 >>
rect 830 1572 219578 219224
<< metal2 >>
rect 742 219200 798 220000
rect 2582 219200 2638 220000
rect 4514 219200 4570 220000
rect 6446 219200 6502 220000
rect 8378 219200 8434 220000
rect 10310 219200 10366 220000
rect 12242 219200 12298 220000
rect 14174 219200 14230 220000
rect 16106 219200 16162 220000
rect 18038 219200 18094 220000
rect 19970 219200 20026 220000
rect 21902 219200 21958 220000
rect 23834 219200 23890 220000
rect 25766 219200 25822 220000
rect 27698 219200 27754 220000
rect 29630 219200 29686 220000
rect 31562 219200 31618 220000
rect 33494 219200 33550 220000
rect 35426 219200 35482 220000
rect 37358 219200 37414 220000
rect 39290 219200 39346 220000
rect 41222 219200 41278 220000
rect 43154 219200 43210 220000
rect 45086 219200 45142 220000
rect 47018 219200 47074 220000
rect 48950 219200 49006 220000
rect 50882 219200 50938 220000
rect 52814 219200 52870 220000
rect 54746 219200 54802 220000
rect 56678 219200 56734 220000
rect 58610 219200 58666 220000
rect 60542 219200 60598 220000
rect 62474 219200 62530 220000
rect 64406 219200 64462 220000
rect 66338 219200 66394 220000
rect 68270 219200 68326 220000
rect 70202 219200 70258 220000
rect 72134 219200 72190 220000
rect 74066 219200 74122 220000
rect 75906 219200 75962 220000
rect 77838 219200 77894 220000
rect 79770 219200 79826 220000
rect 81702 219200 81758 220000
rect 83634 219200 83690 220000
rect 85566 219200 85622 220000
rect 87498 219200 87554 220000
rect 89430 219200 89486 220000
rect 91362 219200 91418 220000
rect 93294 219200 93350 220000
rect 95226 219200 95282 220000
rect 97158 219200 97214 220000
rect 99090 219200 99146 220000
rect 101022 219200 101078 220000
rect 102954 219200 103010 220000
rect 104886 219200 104942 220000
rect 106818 219200 106874 220000
rect 108750 219200 108806 220000
rect 110682 219200 110738 220000
rect 112614 219200 112670 220000
rect 114546 219200 114602 220000
rect 116478 219200 116534 220000
rect 118410 219200 118466 220000
rect 120342 219200 120398 220000
rect 122274 219200 122330 220000
rect 124206 219200 124262 220000
rect 126138 219200 126194 220000
rect 128070 219200 128126 220000
rect 130002 219200 130058 220000
rect 131934 219200 131990 220000
rect 133866 219200 133922 220000
rect 135798 219200 135854 220000
rect 137730 219200 137786 220000
rect 139662 219200 139718 220000
rect 141594 219200 141650 220000
rect 143526 219200 143582 220000
rect 145458 219200 145514 220000
rect 147390 219200 147446 220000
rect 149230 219200 149286 220000
rect 151162 219200 151218 220000
rect 153094 219200 153150 220000
rect 155026 219200 155082 220000
rect 156958 219200 157014 220000
rect 158890 219200 158946 220000
rect 160822 219200 160878 220000
rect 162754 219200 162810 220000
rect 164686 219200 164742 220000
rect 166618 219200 166674 220000
rect 168550 219200 168606 220000
rect 170482 219200 170538 220000
rect 172414 219200 172470 220000
rect 174346 219200 174402 220000
rect 176278 219200 176334 220000
rect 178210 219200 178266 220000
rect 180142 219200 180198 220000
rect 182074 219200 182130 220000
rect 184006 219200 184062 220000
rect 185938 219200 185994 220000
rect 187870 219200 187926 220000
rect 189802 219200 189858 220000
rect 191734 219200 191790 220000
rect 193666 219200 193722 220000
rect 195598 219200 195654 220000
rect 197530 219200 197586 220000
rect 199462 219200 199518 220000
rect 201394 219200 201450 220000
rect 203326 219200 203382 220000
rect 205258 219200 205314 220000
rect 207190 219200 207246 220000
rect 209122 219200 209178 220000
rect 211054 219200 211110 220000
rect 212986 219200 213042 220000
rect 214918 219200 214974 220000
rect 216850 219200 216906 220000
rect 218782 219200 218838 220000
rect 6 0 62 800
rect 374 0 430 800
rect 834 0 890 800
rect 1294 0 1350 800
rect 1754 0 1810 800
rect 2214 0 2270 800
rect 2674 0 2730 800
rect 3134 0 3190 800
rect 3594 0 3650 800
rect 3962 0 4018 800
rect 4422 0 4478 800
rect 4882 0 4938 800
rect 5342 0 5398 800
rect 5802 0 5858 800
rect 6262 0 6318 800
rect 6722 0 6778 800
rect 7182 0 7238 800
rect 7550 0 7606 800
rect 8010 0 8066 800
rect 8470 0 8526 800
rect 8930 0 8986 800
rect 9390 0 9446 800
rect 9850 0 9906 800
rect 10310 0 10366 800
rect 10770 0 10826 800
rect 11138 0 11194 800
rect 11598 0 11654 800
rect 12058 0 12114 800
rect 12518 0 12574 800
rect 12978 0 13034 800
rect 13438 0 13494 800
rect 13898 0 13954 800
rect 14358 0 14414 800
rect 14818 0 14874 800
rect 15186 0 15242 800
rect 15646 0 15702 800
rect 16106 0 16162 800
rect 16566 0 16622 800
rect 17026 0 17082 800
rect 17486 0 17542 800
rect 17946 0 18002 800
rect 18406 0 18462 800
rect 18774 0 18830 800
rect 19234 0 19290 800
rect 19694 0 19750 800
rect 20154 0 20210 800
rect 20614 0 20670 800
rect 21074 0 21130 800
rect 21534 0 21590 800
rect 21994 0 22050 800
rect 22362 0 22418 800
rect 22822 0 22878 800
rect 23282 0 23338 800
rect 23742 0 23798 800
rect 24202 0 24258 800
rect 24662 0 24718 800
rect 25122 0 25178 800
rect 25582 0 25638 800
rect 26042 0 26098 800
rect 26410 0 26466 800
rect 26870 0 26926 800
rect 27330 0 27386 800
rect 27790 0 27846 800
rect 28250 0 28306 800
rect 28710 0 28766 800
rect 29170 0 29226 800
rect 29630 0 29686 800
rect 29998 0 30054 800
rect 30458 0 30514 800
rect 30918 0 30974 800
rect 31378 0 31434 800
rect 31838 0 31894 800
rect 32298 0 32354 800
rect 32758 0 32814 800
rect 33218 0 33274 800
rect 33586 0 33642 800
rect 34046 0 34102 800
rect 34506 0 34562 800
rect 34966 0 35022 800
rect 35426 0 35482 800
rect 35886 0 35942 800
rect 36346 0 36402 800
rect 36806 0 36862 800
rect 37266 0 37322 800
rect 37634 0 37690 800
rect 38094 0 38150 800
rect 38554 0 38610 800
rect 39014 0 39070 800
rect 39474 0 39530 800
rect 39934 0 39990 800
rect 40394 0 40450 800
rect 40854 0 40910 800
rect 41222 0 41278 800
rect 41682 0 41738 800
rect 42142 0 42198 800
rect 42602 0 42658 800
rect 43062 0 43118 800
rect 43522 0 43578 800
rect 43982 0 44038 800
rect 44442 0 44498 800
rect 44810 0 44866 800
rect 45270 0 45326 800
rect 45730 0 45786 800
rect 46190 0 46246 800
rect 46650 0 46706 800
rect 47110 0 47166 800
rect 47570 0 47626 800
rect 48030 0 48086 800
rect 48398 0 48454 800
rect 48858 0 48914 800
rect 49318 0 49374 800
rect 49778 0 49834 800
rect 50238 0 50294 800
rect 50698 0 50754 800
rect 51158 0 51214 800
rect 51618 0 51674 800
rect 52078 0 52134 800
rect 52446 0 52502 800
rect 52906 0 52962 800
rect 53366 0 53422 800
rect 53826 0 53882 800
rect 54286 0 54342 800
rect 54746 0 54802 800
rect 55206 0 55262 800
rect 55666 0 55722 800
rect 56034 0 56090 800
rect 56494 0 56550 800
rect 56954 0 57010 800
rect 57414 0 57470 800
rect 57874 0 57930 800
rect 58334 0 58390 800
rect 58794 0 58850 800
rect 59254 0 59310 800
rect 59622 0 59678 800
rect 60082 0 60138 800
rect 60542 0 60598 800
rect 61002 0 61058 800
rect 61462 0 61518 800
rect 61922 0 61978 800
rect 62382 0 62438 800
rect 62842 0 62898 800
rect 63302 0 63358 800
rect 63670 0 63726 800
rect 64130 0 64186 800
rect 64590 0 64646 800
rect 65050 0 65106 800
rect 65510 0 65566 800
rect 65970 0 66026 800
rect 66430 0 66486 800
rect 66890 0 66946 800
rect 67258 0 67314 800
rect 67718 0 67774 800
rect 68178 0 68234 800
rect 68638 0 68694 800
rect 69098 0 69154 800
rect 69558 0 69614 800
rect 70018 0 70074 800
rect 70478 0 70534 800
rect 70846 0 70902 800
rect 71306 0 71362 800
rect 71766 0 71822 800
rect 72226 0 72282 800
rect 72686 0 72742 800
rect 73146 0 73202 800
rect 73606 0 73662 800
rect 74066 0 74122 800
rect 74526 0 74582 800
rect 74894 0 74950 800
rect 75354 0 75410 800
rect 75814 0 75870 800
rect 76274 0 76330 800
rect 76734 0 76790 800
rect 77194 0 77250 800
rect 77654 0 77710 800
rect 78114 0 78170 800
rect 78482 0 78538 800
rect 78942 0 78998 800
rect 79402 0 79458 800
rect 79862 0 79918 800
rect 80322 0 80378 800
rect 80782 0 80838 800
rect 81242 0 81298 800
rect 81702 0 81758 800
rect 82070 0 82126 800
rect 82530 0 82586 800
rect 82990 0 83046 800
rect 83450 0 83506 800
rect 83910 0 83966 800
rect 84370 0 84426 800
rect 84830 0 84886 800
rect 85290 0 85346 800
rect 85750 0 85806 800
rect 86118 0 86174 800
rect 86578 0 86634 800
rect 87038 0 87094 800
rect 87498 0 87554 800
rect 87958 0 88014 800
rect 88418 0 88474 800
rect 88878 0 88934 800
rect 89338 0 89394 800
rect 89706 0 89762 800
rect 90166 0 90222 800
rect 90626 0 90682 800
rect 91086 0 91142 800
rect 91546 0 91602 800
rect 92006 0 92062 800
rect 92466 0 92522 800
rect 92926 0 92982 800
rect 93294 0 93350 800
rect 93754 0 93810 800
rect 94214 0 94270 800
rect 94674 0 94730 800
rect 95134 0 95190 800
rect 95594 0 95650 800
rect 96054 0 96110 800
rect 96514 0 96570 800
rect 96882 0 96938 800
rect 97342 0 97398 800
rect 97802 0 97858 800
rect 98262 0 98318 800
rect 98722 0 98778 800
rect 99182 0 99238 800
rect 99642 0 99698 800
rect 100102 0 100158 800
rect 100562 0 100618 800
rect 100930 0 100986 800
rect 101390 0 101446 800
rect 101850 0 101906 800
rect 102310 0 102366 800
rect 102770 0 102826 800
rect 103230 0 103286 800
rect 103690 0 103746 800
rect 104150 0 104206 800
rect 104518 0 104574 800
rect 104978 0 105034 800
rect 105438 0 105494 800
rect 105898 0 105954 800
rect 106358 0 106414 800
rect 106818 0 106874 800
rect 107278 0 107334 800
rect 107738 0 107794 800
rect 108106 0 108162 800
rect 108566 0 108622 800
rect 109026 0 109082 800
rect 109486 0 109542 800
rect 109946 0 110002 800
rect 110406 0 110462 800
rect 110866 0 110922 800
rect 111326 0 111382 800
rect 111786 0 111842 800
rect 112154 0 112210 800
rect 112614 0 112670 800
rect 113074 0 113130 800
rect 113534 0 113590 800
rect 113994 0 114050 800
rect 114454 0 114510 800
rect 114914 0 114970 800
rect 115374 0 115430 800
rect 115742 0 115798 800
rect 116202 0 116258 800
rect 116662 0 116718 800
rect 117122 0 117178 800
rect 117582 0 117638 800
rect 118042 0 118098 800
rect 118502 0 118558 800
rect 118962 0 119018 800
rect 119330 0 119386 800
rect 119790 0 119846 800
rect 120250 0 120306 800
rect 120710 0 120766 800
rect 121170 0 121226 800
rect 121630 0 121686 800
rect 122090 0 122146 800
rect 122550 0 122606 800
rect 123010 0 123066 800
rect 123378 0 123434 800
rect 123838 0 123894 800
rect 124298 0 124354 800
rect 124758 0 124814 800
rect 125218 0 125274 800
rect 125678 0 125734 800
rect 126138 0 126194 800
rect 126598 0 126654 800
rect 126966 0 127022 800
rect 127426 0 127482 800
rect 127886 0 127942 800
rect 128346 0 128402 800
rect 128806 0 128862 800
rect 129266 0 129322 800
rect 129726 0 129782 800
rect 130186 0 130242 800
rect 130554 0 130610 800
rect 131014 0 131070 800
rect 131474 0 131530 800
rect 131934 0 131990 800
rect 132394 0 132450 800
rect 132854 0 132910 800
rect 133314 0 133370 800
rect 133774 0 133830 800
rect 134142 0 134198 800
rect 134602 0 134658 800
rect 135062 0 135118 800
rect 135522 0 135578 800
rect 135982 0 136038 800
rect 136442 0 136498 800
rect 136902 0 136958 800
rect 137362 0 137418 800
rect 137822 0 137878 800
rect 138190 0 138246 800
rect 138650 0 138706 800
rect 139110 0 139166 800
rect 139570 0 139626 800
rect 140030 0 140086 800
rect 140490 0 140546 800
rect 140950 0 141006 800
rect 141410 0 141466 800
rect 141778 0 141834 800
rect 142238 0 142294 800
rect 142698 0 142754 800
rect 143158 0 143214 800
rect 143618 0 143674 800
rect 144078 0 144134 800
rect 144538 0 144594 800
rect 144998 0 145054 800
rect 145366 0 145422 800
rect 145826 0 145882 800
rect 146286 0 146342 800
rect 146746 0 146802 800
rect 147206 0 147262 800
rect 147666 0 147722 800
rect 148126 0 148182 800
rect 148586 0 148642 800
rect 149046 0 149102 800
rect 149414 0 149470 800
rect 149874 0 149930 800
rect 150334 0 150390 800
rect 150794 0 150850 800
rect 151254 0 151310 800
rect 151714 0 151770 800
rect 152174 0 152230 800
rect 152634 0 152690 800
rect 153002 0 153058 800
rect 153462 0 153518 800
rect 153922 0 153978 800
rect 154382 0 154438 800
rect 154842 0 154898 800
rect 155302 0 155358 800
rect 155762 0 155818 800
rect 156222 0 156278 800
rect 156590 0 156646 800
rect 157050 0 157106 800
rect 157510 0 157566 800
rect 157970 0 158026 800
rect 158430 0 158486 800
rect 158890 0 158946 800
rect 159350 0 159406 800
rect 159810 0 159866 800
rect 160270 0 160326 800
rect 160638 0 160694 800
rect 161098 0 161154 800
rect 161558 0 161614 800
rect 162018 0 162074 800
rect 162478 0 162534 800
rect 162938 0 162994 800
rect 163398 0 163454 800
rect 163858 0 163914 800
rect 164226 0 164282 800
rect 164686 0 164742 800
rect 165146 0 165202 800
rect 165606 0 165662 800
rect 166066 0 166122 800
rect 166526 0 166582 800
rect 166986 0 167042 800
rect 167446 0 167502 800
rect 167814 0 167870 800
rect 168274 0 168330 800
rect 168734 0 168790 800
rect 169194 0 169250 800
rect 169654 0 169710 800
rect 170114 0 170170 800
rect 170574 0 170630 800
rect 171034 0 171090 800
rect 171494 0 171550 800
rect 171862 0 171918 800
rect 172322 0 172378 800
rect 172782 0 172838 800
rect 173242 0 173298 800
rect 173702 0 173758 800
rect 174162 0 174218 800
rect 174622 0 174678 800
rect 175082 0 175138 800
rect 175450 0 175506 800
rect 175910 0 175966 800
rect 176370 0 176426 800
rect 176830 0 176886 800
rect 177290 0 177346 800
rect 177750 0 177806 800
rect 178210 0 178266 800
rect 178670 0 178726 800
rect 179038 0 179094 800
rect 179498 0 179554 800
rect 179958 0 180014 800
rect 180418 0 180474 800
rect 180878 0 180934 800
rect 181338 0 181394 800
rect 181798 0 181854 800
rect 182258 0 182314 800
rect 182626 0 182682 800
rect 183086 0 183142 800
rect 183546 0 183602 800
rect 184006 0 184062 800
rect 184466 0 184522 800
rect 184926 0 184982 800
rect 185386 0 185442 800
rect 185846 0 185902 800
rect 186306 0 186362 800
rect 186674 0 186730 800
rect 187134 0 187190 800
rect 187594 0 187650 800
rect 188054 0 188110 800
rect 188514 0 188570 800
rect 188974 0 189030 800
rect 189434 0 189490 800
rect 189894 0 189950 800
rect 190262 0 190318 800
rect 190722 0 190778 800
rect 191182 0 191238 800
rect 191642 0 191698 800
rect 192102 0 192158 800
rect 192562 0 192618 800
rect 193022 0 193078 800
rect 193482 0 193538 800
rect 193850 0 193906 800
rect 194310 0 194366 800
rect 194770 0 194826 800
rect 195230 0 195286 800
rect 195690 0 195746 800
rect 196150 0 196206 800
rect 196610 0 196666 800
rect 197070 0 197126 800
rect 197530 0 197586 800
rect 197898 0 197954 800
rect 198358 0 198414 800
rect 198818 0 198874 800
rect 199278 0 199334 800
rect 199738 0 199794 800
rect 200198 0 200254 800
rect 200658 0 200714 800
rect 201118 0 201174 800
rect 201486 0 201542 800
rect 201946 0 202002 800
rect 202406 0 202462 800
rect 202866 0 202922 800
rect 203326 0 203382 800
rect 203786 0 203842 800
rect 204246 0 204302 800
rect 204706 0 204762 800
rect 205074 0 205130 800
rect 205534 0 205590 800
rect 205994 0 206050 800
rect 206454 0 206510 800
rect 206914 0 206970 800
rect 207374 0 207430 800
rect 207834 0 207890 800
rect 208294 0 208350 800
rect 208754 0 208810 800
rect 209122 0 209178 800
rect 209582 0 209638 800
rect 210042 0 210098 800
rect 210502 0 210558 800
rect 210962 0 211018 800
rect 211422 0 211478 800
rect 211882 0 211938 800
rect 212342 0 212398 800
rect 212710 0 212766 800
rect 213170 0 213226 800
rect 213630 0 213686 800
rect 214090 0 214146 800
rect 214550 0 214606 800
rect 215010 0 215066 800
rect 215470 0 215526 800
rect 215930 0 215986 800
rect 216298 0 216354 800
rect 216758 0 216814 800
rect 217218 0 217274 800
rect 217678 0 217734 800
rect 218138 0 218194 800
rect 218598 0 218654 800
rect 219058 0 219114 800
rect 219518 0 219574 800
<< obsm2 >>
rect 6 219144 686 219230
rect 854 219144 2526 219230
rect 2694 219144 4458 219230
rect 4626 219144 6390 219230
rect 6558 219144 8322 219230
rect 8490 219144 10254 219230
rect 10422 219144 12186 219230
rect 12354 219144 14118 219230
rect 14286 219144 16050 219230
rect 16218 219144 17982 219230
rect 18150 219144 19914 219230
rect 20082 219144 21846 219230
rect 22014 219144 23778 219230
rect 23946 219144 25710 219230
rect 25878 219144 27642 219230
rect 27810 219144 29574 219230
rect 29742 219144 31506 219230
rect 31674 219144 33438 219230
rect 33606 219144 35370 219230
rect 35538 219144 37302 219230
rect 37470 219144 39234 219230
rect 39402 219144 41166 219230
rect 41334 219144 43098 219230
rect 43266 219144 45030 219230
rect 45198 219144 46962 219230
rect 47130 219144 48894 219230
rect 49062 219144 50826 219230
rect 50994 219144 52758 219230
rect 52926 219144 54690 219230
rect 54858 219144 56622 219230
rect 56790 219144 58554 219230
rect 58722 219144 60486 219230
rect 60654 219144 62418 219230
rect 62586 219144 64350 219230
rect 64518 219144 66282 219230
rect 66450 219144 68214 219230
rect 68382 219144 70146 219230
rect 70314 219144 72078 219230
rect 72246 219144 74010 219230
rect 74178 219144 75850 219230
rect 76018 219144 77782 219230
rect 77950 219144 79714 219230
rect 79882 219144 81646 219230
rect 81814 219144 83578 219230
rect 83746 219144 85510 219230
rect 85678 219144 87442 219230
rect 87610 219144 89374 219230
rect 89542 219144 91306 219230
rect 91474 219144 93238 219230
rect 93406 219144 95170 219230
rect 95338 219144 97102 219230
rect 97270 219144 99034 219230
rect 99202 219144 100966 219230
rect 101134 219144 102898 219230
rect 103066 219144 104830 219230
rect 104998 219144 106762 219230
rect 106930 219144 108694 219230
rect 108862 219144 110626 219230
rect 110794 219144 112558 219230
rect 112726 219144 114490 219230
rect 114658 219144 116422 219230
rect 116590 219144 118354 219230
rect 118522 219144 120286 219230
rect 120454 219144 122218 219230
rect 122386 219144 124150 219230
rect 124318 219144 126082 219230
rect 126250 219144 128014 219230
rect 128182 219144 129946 219230
rect 130114 219144 131878 219230
rect 132046 219144 133810 219230
rect 133978 219144 135742 219230
rect 135910 219144 137674 219230
rect 137842 219144 139606 219230
rect 139774 219144 141538 219230
rect 141706 219144 143470 219230
rect 143638 219144 145402 219230
rect 145570 219144 147334 219230
rect 147502 219144 149174 219230
rect 149342 219144 151106 219230
rect 151274 219144 153038 219230
rect 153206 219144 154970 219230
rect 155138 219144 156902 219230
rect 157070 219144 158834 219230
rect 159002 219144 160766 219230
rect 160934 219144 162698 219230
rect 162866 219144 164630 219230
rect 164798 219144 166562 219230
rect 166730 219144 168494 219230
rect 168662 219144 170426 219230
rect 170594 219144 172358 219230
rect 172526 219144 174290 219230
rect 174458 219144 176222 219230
rect 176390 219144 178154 219230
rect 178322 219144 180086 219230
rect 180254 219144 182018 219230
rect 182186 219144 183950 219230
rect 184118 219144 185882 219230
rect 186050 219144 187814 219230
rect 187982 219144 189746 219230
rect 189914 219144 191678 219230
rect 191846 219144 193610 219230
rect 193778 219144 195542 219230
rect 195710 219144 197474 219230
rect 197642 219144 199406 219230
rect 199574 219144 201338 219230
rect 201506 219144 203270 219230
rect 203438 219144 205202 219230
rect 205370 219144 207134 219230
rect 207302 219144 209066 219230
rect 209234 219144 210998 219230
rect 211166 219144 212930 219230
rect 213098 219144 214862 219230
rect 215030 219144 216794 219230
rect 216962 219144 218726 219230
rect 218894 219144 219572 219230
rect 6 856 219572 219144
rect 118 800 318 856
rect 486 800 778 856
rect 946 800 1238 856
rect 1406 800 1698 856
rect 1866 800 2158 856
rect 2326 800 2618 856
rect 2786 800 3078 856
rect 3246 800 3538 856
rect 3706 800 3906 856
rect 4074 800 4366 856
rect 4534 800 4826 856
rect 4994 800 5286 856
rect 5454 800 5746 856
rect 5914 800 6206 856
rect 6374 800 6666 856
rect 6834 800 7126 856
rect 7294 800 7494 856
rect 7662 800 7954 856
rect 8122 800 8414 856
rect 8582 800 8874 856
rect 9042 800 9334 856
rect 9502 800 9794 856
rect 9962 800 10254 856
rect 10422 800 10714 856
rect 10882 800 11082 856
rect 11250 800 11542 856
rect 11710 800 12002 856
rect 12170 800 12462 856
rect 12630 800 12922 856
rect 13090 800 13382 856
rect 13550 800 13842 856
rect 14010 800 14302 856
rect 14470 800 14762 856
rect 14930 800 15130 856
rect 15298 800 15590 856
rect 15758 800 16050 856
rect 16218 800 16510 856
rect 16678 800 16970 856
rect 17138 800 17430 856
rect 17598 800 17890 856
rect 18058 800 18350 856
rect 18518 800 18718 856
rect 18886 800 19178 856
rect 19346 800 19638 856
rect 19806 800 20098 856
rect 20266 800 20558 856
rect 20726 800 21018 856
rect 21186 800 21478 856
rect 21646 800 21938 856
rect 22106 800 22306 856
rect 22474 800 22766 856
rect 22934 800 23226 856
rect 23394 800 23686 856
rect 23854 800 24146 856
rect 24314 800 24606 856
rect 24774 800 25066 856
rect 25234 800 25526 856
rect 25694 800 25986 856
rect 26154 800 26354 856
rect 26522 800 26814 856
rect 26982 800 27274 856
rect 27442 800 27734 856
rect 27902 800 28194 856
rect 28362 800 28654 856
rect 28822 800 29114 856
rect 29282 800 29574 856
rect 29742 800 29942 856
rect 30110 800 30402 856
rect 30570 800 30862 856
rect 31030 800 31322 856
rect 31490 800 31782 856
rect 31950 800 32242 856
rect 32410 800 32702 856
rect 32870 800 33162 856
rect 33330 800 33530 856
rect 33698 800 33990 856
rect 34158 800 34450 856
rect 34618 800 34910 856
rect 35078 800 35370 856
rect 35538 800 35830 856
rect 35998 800 36290 856
rect 36458 800 36750 856
rect 36918 800 37210 856
rect 37378 800 37578 856
rect 37746 800 38038 856
rect 38206 800 38498 856
rect 38666 800 38958 856
rect 39126 800 39418 856
rect 39586 800 39878 856
rect 40046 800 40338 856
rect 40506 800 40798 856
rect 40966 800 41166 856
rect 41334 800 41626 856
rect 41794 800 42086 856
rect 42254 800 42546 856
rect 42714 800 43006 856
rect 43174 800 43466 856
rect 43634 800 43926 856
rect 44094 800 44386 856
rect 44554 800 44754 856
rect 44922 800 45214 856
rect 45382 800 45674 856
rect 45842 800 46134 856
rect 46302 800 46594 856
rect 46762 800 47054 856
rect 47222 800 47514 856
rect 47682 800 47974 856
rect 48142 800 48342 856
rect 48510 800 48802 856
rect 48970 800 49262 856
rect 49430 800 49722 856
rect 49890 800 50182 856
rect 50350 800 50642 856
rect 50810 800 51102 856
rect 51270 800 51562 856
rect 51730 800 52022 856
rect 52190 800 52390 856
rect 52558 800 52850 856
rect 53018 800 53310 856
rect 53478 800 53770 856
rect 53938 800 54230 856
rect 54398 800 54690 856
rect 54858 800 55150 856
rect 55318 800 55610 856
rect 55778 800 55978 856
rect 56146 800 56438 856
rect 56606 800 56898 856
rect 57066 800 57358 856
rect 57526 800 57818 856
rect 57986 800 58278 856
rect 58446 800 58738 856
rect 58906 800 59198 856
rect 59366 800 59566 856
rect 59734 800 60026 856
rect 60194 800 60486 856
rect 60654 800 60946 856
rect 61114 800 61406 856
rect 61574 800 61866 856
rect 62034 800 62326 856
rect 62494 800 62786 856
rect 62954 800 63246 856
rect 63414 800 63614 856
rect 63782 800 64074 856
rect 64242 800 64534 856
rect 64702 800 64994 856
rect 65162 800 65454 856
rect 65622 800 65914 856
rect 66082 800 66374 856
rect 66542 800 66834 856
rect 67002 800 67202 856
rect 67370 800 67662 856
rect 67830 800 68122 856
rect 68290 800 68582 856
rect 68750 800 69042 856
rect 69210 800 69502 856
rect 69670 800 69962 856
rect 70130 800 70422 856
rect 70590 800 70790 856
rect 70958 800 71250 856
rect 71418 800 71710 856
rect 71878 800 72170 856
rect 72338 800 72630 856
rect 72798 800 73090 856
rect 73258 800 73550 856
rect 73718 800 74010 856
rect 74178 800 74470 856
rect 74638 800 74838 856
rect 75006 800 75298 856
rect 75466 800 75758 856
rect 75926 800 76218 856
rect 76386 800 76678 856
rect 76846 800 77138 856
rect 77306 800 77598 856
rect 77766 800 78058 856
rect 78226 800 78426 856
rect 78594 800 78886 856
rect 79054 800 79346 856
rect 79514 800 79806 856
rect 79974 800 80266 856
rect 80434 800 80726 856
rect 80894 800 81186 856
rect 81354 800 81646 856
rect 81814 800 82014 856
rect 82182 800 82474 856
rect 82642 800 82934 856
rect 83102 800 83394 856
rect 83562 800 83854 856
rect 84022 800 84314 856
rect 84482 800 84774 856
rect 84942 800 85234 856
rect 85402 800 85694 856
rect 85862 800 86062 856
rect 86230 800 86522 856
rect 86690 800 86982 856
rect 87150 800 87442 856
rect 87610 800 87902 856
rect 88070 800 88362 856
rect 88530 800 88822 856
rect 88990 800 89282 856
rect 89450 800 89650 856
rect 89818 800 90110 856
rect 90278 800 90570 856
rect 90738 800 91030 856
rect 91198 800 91490 856
rect 91658 800 91950 856
rect 92118 800 92410 856
rect 92578 800 92870 856
rect 93038 800 93238 856
rect 93406 800 93698 856
rect 93866 800 94158 856
rect 94326 800 94618 856
rect 94786 800 95078 856
rect 95246 800 95538 856
rect 95706 800 95998 856
rect 96166 800 96458 856
rect 96626 800 96826 856
rect 96994 800 97286 856
rect 97454 800 97746 856
rect 97914 800 98206 856
rect 98374 800 98666 856
rect 98834 800 99126 856
rect 99294 800 99586 856
rect 99754 800 100046 856
rect 100214 800 100506 856
rect 100674 800 100874 856
rect 101042 800 101334 856
rect 101502 800 101794 856
rect 101962 800 102254 856
rect 102422 800 102714 856
rect 102882 800 103174 856
rect 103342 800 103634 856
rect 103802 800 104094 856
rect 104262 800 104462 856
rect 104630 800 104922 856
rect 105090 800 105382 856
rect 105550 800 105842 856
rect 106010 800 106302 856
rect 106470 800 106762 856
rect 106930 800 107222 856
rect 107390 800 107682 856
rect 107850 800 108050 856
rect 108218 800 108510 856
rect 108678 800 108970 856
rect 109138 800 109430 856
rect 109598 800 109890 856
rect 110058 800 110350 856
rect 110518 800 110810 856
rect 110978 800 111270 856
rect 111438 800 111730 856
rect 111898 800 112098 856
rect 112266 800 112558 856
rect 112726 800 113018 856
rect 113186 800 113478 856
rect 113646 800 113938 856
rect 114106 800 114398 856
rect 114566 800 114858 856
rect 115026 800 115318 856
rect 115486 800 115686 856
rect 115854 800 116146 856
rect 116314 800 116606 856
rect 116774 800 117066 856
rect 117234 800 117526 856
rect 117694 800 117986 856
rect 118154 800 118446 856
rect 118614 800 118906 856
rect 119074 800 119274 856
rect 119442 800 119734 856
rect 119902 800 120194 856
rect 120362 800 120654 856
rect 120822 800 121114 856
rect 121282 800 121574 856
rect 121742 800 122034 856
rect 122202 800 122494 856
rect 122662 800 122954 856
rect 123122 800 123322 856
rect 123490 800 123782 856
rect 123950 800 124242 856
rect 124410 800 124702 856
rect 124870 800 125162 856
rect 125330 800 125622 856
rect 125790 800 126082 856
rect 126250 800 126542 856
rect 126710 800 126910 856
rect 127078 800 127370 856
rect 127538 800 127830 856
rect 127998 800 128290 856
rect 128458 800 128750 856
rect 128918 800 129210 856
rect 129378 800 129670 856
rect 129838 800 130130 856
rect 130298 800 130498 856
rect 130666 800 130958 856
rect 131126 800 131418 856
rect 131586 800 131878 856
rect 132046 800 132338 856
rect 132506 800 132798 856
rect 132966 800 133258 856
rect 133426 800 133718 856
rect 133886 800 134086 856
rect 134254 800 134546 856
rect 134714 800 135006 856
rect 135174 800 135466 856
rect 135634 800 135926 856
rect 136094 800 136386 856
rect 136554 800 136846 856
rect 137014 800 137306 856
rect 137474 800 137766 856
rect 137934 800 138134 856
rect 138302 800 138594 856
rect 138762 800 139054 856
rect 139222 800 139514 856
rect 139682 800 139974 856
rect 140142 800 140434 856
rect 140602 800 140894 856
rect 141062 800 141354 856
rect 141522 800 141722 856
rect 141890 800 142182 856
rect 142350 800 142642 856
rect 142810 800 143102 856
rect 143270 800 143562 856
rect 143730 800 144022 856
rect 144190 800 144482 856
rect 144650 800 144942 856
rect 145110 800 145310 856
rect 145478 800 145770 856
rect 145938 800 146230 856
rect 146398 800 146690 856
rect 146858 800 147150 856
rect 147318 800 147610 856
rect 147778 800 148070 856
rect 148238 800 148530 856
rect 148698 800 148990 856
rect 149158 800 149358 856
rect 149526 800 149818 856
rect 149986 800 150278 856
rect 150446 800 150738 856
rect 150906 800 151198 856
rect 151366 800 151658 856
rect 151826 800 152118 856
rect 152286 800 152578 856
rect 152746 800 152946 856
rect 153114 800 153406 856
rect 153574 800 153866 856
rect 154034 800 154326 856
rect 154494 800 154786 856
rect 154954 800 155246 856
rect 155414 800 155706 856
rect 155874 800 156166 856
rect 156334 800 156534 856
rect 156702 800 156994 856
rect 157162 800 157454 856
rect 157622 800 157914 856
rect 158082 800 158374 856
rect 158542 800 158834 856
rect 159002 800 159294 856
rect 159462 800 159754 856
rect 159922 800 160214 856
rect 160382 800 160582 856
rect 160750 800 161042 856
rect 161210 800 161502 856
rect 161670 800 161962 856
rect 162130 800 162422 856
rect 162590 800 162882 856
rect 163050 800 163342 856
rect 163510 800 163802 856
rect 163970 800 164170 856
rect 164338 800 164630 856
rect 164798 800 165090 856
rect 165258 800 165550 856
rect 165718 800 166010 856
rect 166178 800 166470 856
rect 166638 800 166930 856
rect 167098 800 167390 856
rect 167558 800 167758 856
rect 167926 800 168218 856
rect 168386 800 168678 856
rect 168846 800 169138 856
rect 169306 800 169598 856
rect 169766 800 170058 856
rect 170226 800 170518 856
rect 170686 800 170978 856
rect 171146 800 171438 856
rect 171606 800 171806 856
rect 171974 800 172266 856
rect 172434 800 172726 856
rect 172894 800 173186 856
rect 173354 800 173646 856
rect 173814 800 174106 856
rect 174274 800 174566 856
rect 174734 800 175026 856
rect 175194 800 175394 856
rect 175562 800 175854 856
rect 176022 800 176314 856
rect 176482 800 176774 856
rect 176942 800 177234 856
rect 177402 800 177694 856
rect 177862 800 178154 856
rect 178322 800 178614 856
rect 178782 800 178982 856
rect 179150 800 179442 856
rect 179610 800 179902 856
rect 180070 800 180362 856
rect 180530 800 180822 856
rect 180990 800 181282 856
rect 181450 800 181742 856
rect 181910 800 182202 856
rect 182370 800 182570 856
rect 182738 800 183030 856
rect 183198 800 183490 856
rect 183658 800 183950 856
rect 184118 800 184410 856
rect 184578 800 184870 856
rect 185038 800 185330 856
rect 185498 800 185790 856
rect 185958 800 186250 856
rect 186418 800 186618 856
rect 186786 800 187078 856
rect 187246 800 187538 856
rect 187706 800 187998 856
rect 188166 800 188458 856
rect 188626 800 188918 856
rect 189086 800 189378 856
rect 189546 800 189838 856
rect 190006 800 190206 856
rect 190374 800 190666 856
rect 190834 800 191126 856
rect 191294 800 191586 856
rect 191754 800 192046 856
rect 192214 800 192506 856
rect 192674 800 192966 856
rect 193134 800 193426 856
rect 193594 800 193794 856
rect 193962 800 194254 856
rect 194422 800 194714 856
rect 194882 800 195174 856
rect 195342 800 195634 856
rect 195802 800 196094 856
rect 196262 800 196554 856
rect 196722 800 197014 856
rect 197182 800 197474 856
rect 197642 800 197842 856
rect 198010 800 198302 856
rect 198470 800 198762 856
rect 198930 800 199222 856
rect 199390 800 199682 856
rect 199850 800 200142 856
rect 200310 800 200602 856
rect 200770 800 201062 856
rect 201230 800 201430 856
rect 201598 800 201890 856
rect 202058 800 202350 856
rect 202518 800 202810 856
rect 202978 800 203270 856
rect 203438 800 203730 856
rect 203898 800 204190 856
rect 204358 800 204650 856
rect 204818 800 205018 856
rect 205186 800 205478 856
rect 205646 800 205938 856
rect 206106 800 206398 856
rect 206566 800 206858 856
rect 207026 800 207318 856
rect 207486 800 207778 856
rect 207946 800 208238 856
rect 208406 800 208698 856
rect 208866 800 209066 856
rect 209234 800 209526 856
rect 209694 800 209986 856
rect 210154 800 210446 856
rect 210614 800 210906 856
rect 211074 800 211366 856
rect 211534 800 211826 856
rect 211994 800 212286 856
rect 212454 800 212654 856
rect 212822 800 213114 856
rect 213282 800 213574 856
rect 213742 800 214034 856
rect 214202 800 214494 856
rect 214662 800 214954 856
rect 215122 800 215414 856
rect 215582 800 215874 856
rect 216042 800 216242 856
rect 216410 800 216702 856
rect 216870 800 217162 856
rect 217330 800 217622 856
rect 217790 800 218082 856
rect 218250 800 218542 856
rect 218710 800 219002 856
rect 219170 800 219462 856
<< obsm3 >>
rect 1 851 215807 217633
<< metal4 >>
rect 4012 2128 4332 217648
rect 19372 2128 19692 217648
<< obsm4 >>
rect 9063 2128 19292 217648
rect 19772 2128 213737 217648
<< labels >>
rlabel metal2 s 742 219200 798 220000 6 io_in[0]
port 1 nsew default input
rlabel metal2 s 58610 219200 58666 220000 6 io_in[10]
port 2 nsew default input
rlabel metal2 s 64406 219200 64462 220000 6 io_in[11]
port 3 nsew default input
rlabel metal2 s 70202 219200 70258 220000 6 io_in[12]
port 4 nsew default input
rlabel metal2 s 75906 219200 75962 220000 6 io_in[13]
port 5 nsew default input
rlabel metal2 s 81702 219200 81758 220000 6 io_in[14]
port 6 nsew default input
rlabel metal2 s 87498 219200 87554 220000 6 io_in[15]
port 7 nsew default input
rlabel metal2 s 93294 219200 93350 220000 6 io_in[16]
port 8 nsew default input
rlabel metal2 s 99090 219200 99146 220000 6 io_in[17]
port 9 nsew default input
rlabel metal2 s 104886 219200 104942 220000 6 io_in[18]
port 10 nsew default input
rlabel metal2 s 110682 219200 110738 220000 6 io_in[19]
port 11 nsew default input
rlabel metal2 s 6446 219200 6502 220000 6 io_in[1]
port 12 nsew default input
rlabel metal2 s 116478 219200 116534 220000 6 io_in[20]
port 13 nsew default input
rlabel metal2 s 122274 219200 122330 220000 6 io_in[21]
port 14 nsew default input
rlabel metal2 s 128070 219200 128126 220000 6 io_in[22]
port 15 nsew default input
rlabel metal2 s 133866 219200 133922 220000 6 io_in[23]
port 16 nsew default input
rlabel metal2 s 139662 219200 139718 220000 6 io_in[24]
port 17 nsew default input
rlabel metal2 s 145458 219200 145514 220000 6 io_in[25]
port 18 nsew default input
rlabel metal2 s 151162 219200 151218 220000 6 io_in[26]
port 19 nsew default input
rlabel metal2 s 156958 219200 157014 220000 6 io_in[27]
port 20 nsew default input
rlabel metal2 s 162754 219200 162810 220000 6 io_in[28]
port 21 nsew default input
rlabel metal2 s 168550 219200 168606 220000 6 io_in[29]
port 22 nsew default input
rlabel metal2 s 12242 219200 12298 220000 6 io_in[2]
port 23 nsew default input
rlabel metal2 s 174346 219200 174402 220000 6 io_in[30]
port 24 nsew default input
rlabel metal2 s 180142 219200 180198 220000 6 io_in[31]
port 25 nsew default input
rlabel metal2 s 185938 219200 185994 220000 6 io_in[32]
port 26 nsew default input
rlabel metal2 s 191734 219200 191790 220000 6 io_in[33]
port 27 nsew default input
rlabel metal2 s 197530 219200 197586 220000 6 io_in[34]
port 28 nsew default input
rlabel metal2 s 203326 219200 203382 220000 6 io_in[35]
port 29 nsew default input
rlabel metal2 s 209122 219200 209178 220000 6 io_in[36]
port 30 nsew default input
rlabel metal2 s 214918 219200 214974 220000 6 io_in[37]
port 31 nsew default input
rlabel metal2 s 18038 219200 18094 220000 6 io_in[3]
port 32 nsew default input
rlabel metal2 s 23834 219200 23890 220000 6 io_in[4]
port 33 nsew default input
rlabel metal2 s 29630 219200 29686 220000 6 io_in[5]
port 34 nsew default input
rlabel metal2 s 35426 219200 35482 220000 6 io_in[6]
port 35 nsew default input
rlabel metal2 s 41222 219200 41278 220000 6 io_in[7]
port 36 nsew default input
rlabel metal2 s 47018 219200 47074 220000 6 io_in[8]
port 37 nsew default input
rlabel metal2 s 52814 219200 52870 220000 6 io_in[9]
port 38 nsew default input
rlabel metal2 s 2582 219200 2638 220000 6 io_oeb[0]
port 39 nsew default output
rlabel metal2 s 60542 219200 60598 220000 6 io_oeb[10]
port 40 nsew default output
rlabel metal2 s 66338 219200 66394 220000 6 io_oeb[11]
port 41 nsew default output
rlabel metal2 s 72134 219200 72190 220000 6 io_oeb[12]
port 42 nsew default output
rlabel metal2 s 77838 219200 77894 220000 6 io_oeb[13]
port 43 nsew default output
rlabel metal2 s 83634 219200 83690 220000 6 io_oeb[14]
port 44 nsew default output
rlabel metal2 s 89430 219200 89486 220000 6 io_oeb[15]
port 45 nsew default output
rlabel metal2 s 95226 219200 95282 220000 6 io_oeb[16]
port 46 nsew default output
rlabel metal2 s 101022 219200 101078 220000 6 io_oeb[17]
port 47 nsew default output
rlabel metal2 s 106818 219200 106874 220000 6 io_oeb[18]
port 48 nsew default output
rlabel metal2 s 112614 219200 112670 220000 6 io_oeb[19]
port 49 nsew default output
rlabel metal2 s 8378 219200 8434 220000 6 io_oeb[1]
port 50 nsew default output
rlabel metal2 s 118410 219200 118466 220000 6 io_oeb[20]
port 51 nsew default output
rlabel metal2 s 124206 219200 124262 220000 6 io_oeb[21]
port 52 nsew default output
rlabel metal2 s 130002 219200 130058 220000 6 io_oeb[22]
port 53 nsew default output
rlabel metal2 s 135798 219200 135854 220000 6 io_oeb[23]
port 54 nsew default output
rlabel metal2 s 141594 219200 141650 220000 6 io_oeb[24]
port 55 nsew default output
rlabel metal2 s 147390 219200 147446 220000 6 io_oeb[25]
port 56 nsew default output
rlabel metal2 s 153094 219200 153150 220000 6 io_oeb[26]
port 57 nsew default output
rlabel metal2 s 158890 219200 158946 220000 6 io_oeb[27]
port 58 nsew default output
rlabel metal2 s 164686 219200 164742 220000 6 io_oeb[28]
port 59 nsew default output
rlabel metal2 s 170482 219200 170538 220000 6 io_oeb[29]
port 60 nsew default output
rlabel metal2 s 14174 219200 14230 220000 6 io_oeb[2]
port 61 nsew default output
rlabel metal2 s 176278 219200 176334 220000 6 io_oeb[30]
port 62 nsew default output
rlabel metal2 s 182074 219200 182130 220000 6 io_oeb[31]
port 63 nsew default output
rlabel metal2 s 187870 219200 187926 220000 6 io_oeb[32]
port 64 nsew default output
rlabel metal2 s 193666 219200 193722 220000 6 io_oeb[33]
port 65 nsew default output
rlabel metal2 s 199462 219200 199518 220000 6 io_oeb[34]
port 66 nsew default output
rlabel metal2 s 205258 219200 205314 220000 6 io_oeb[35]
port 67 nsew default output
rlabel metal2 s 211054 219200 211110 220000 6 io_oeb[36]
port 68 nsew default output
rlabel metal2 s 216850 219200 216906 220000 6 io_oeb[37]
port 69 nsew default output
rlabel metal2 s 19970 219200 20026 220000 6 io_oeb[3]
port 70 nsew default output
rlabel metal2 s 25766 219200 25822 220000 6 io_oeb[4]
port 71 nsew default output
rlabel metal2 s 31562 219200 31618 220000 6 io_oeb[5]
port 72 nsew default output
rlabel metal2 s 37358 219200 37414 220000 6 io_oeb[6]
port 73 nsew default output
rlabel metal2 s 43154 219200 43210 220000 6 io_oeb[7]
port 74 nsew default output
rlabel metal2 s 48950 219200 49006 220000 6 io_oeb[8]
port 75 nsew default output
rlabel metal2 s 54746 219200 54802 220000 6 io_oeb[9]
port 76 nsew default output
rlabel metal2 s 4514 219200 4570 220000 6 io_out[0]
port 77 nsew default output
rlabel metal2 s 62474 219200 62530 220000 6 io_out[10]
port 78 nsew default output
rlabel metal2 s 68270 219200 68326 220000 6 io_out[11]
port 79 nsew default output
rlabel metal2 s 74066 219200 74122 220000 6 io_out[12]
port 80 nsew default output
rlabel metal2 s 79770 219200 79826 220000 6 io_out[13]
port 81 nsew default output
rlabel metal2 s 85566 219200 85622 220000 6 io_out[14]
port 82 nsew default output
rlabel metal2 s 91362 219200 91418 220000 6 io_out[15]
port 83 nsew default output
rlabel metal2 s 97158 219200 97214 220000 6 io_out[16]
port 84 nsew default output
rlabel metal2 s 102954 219200 103010 220000 6 io_out[17]
port 85 nsew default output
rlabel metal2 s 108750 219200 108806 220000 6 io_out[18]
port 86 nsew default output
rlabel metal2 s 114546 219200 114602 220000 6 io_out[19]
port 87 nsew default output
rlabel metal2 s 10310 219200 10366 220000 6 io_out[1]
port 88 nsew default output
rlabel metal2 s 120342 219200 120398 220000 6 io_out[20]
port 89 nsew default output
rlabel metal2 s 126138 219200 126194 220000 6 io_out[21]
port 90 nsew default output
rlabel metal2 s 131934 219200 131990 220000 6 io_out[22]
port 91 nsew default output
rlabel metal2 s 137730 219200 137786 220000 6 io_out[23]
port 92 nsew default output
rlabel metal2 s 143526 219200 143582 220000 6 io_out[24]
port 93 nsew default output
rlabel metal2 s 149230 219200 149286 220000 6 io_out[25]
port 94 nsew default output
rlabel metal2 s 155026 219200 155082 220000 6 io_out[26]
port 95 nsew default output
rlabel metal2 s 160822 219200 160878 220000 6 io_out[27]
port 96 nsew default output
rlabel metal2 s 166618 219200 166674 220000 6 io_out[28]
port 97 nsew default output
rlabel metal2 s 172414 219200 172470 220000 6 io_out[29]
port 98 nsew default output
rlabel metal2 s 16106 219200 16162 220000 6 io_out[2]
port 99 nsew default output
rlabel metal2 s 178210 219200 178266 220000 6 io_out[30]
port 100 nsew default output
rlabel metal2 s 184006 219200 184062 220000 6 io_out[31]
port 101 nsew default output
rlabel metal2 s 189802 219200 189858 220000 6 io_out[32]
port 102 nsew default output
rlabel metal2 s 195598 219200 195654 220000 6 io_out[33]
port 103 nsew default output
rlabel metal2 s 201394 219200 201450 220000 6 io_out[34]
port 104 nsew default output
rlabel metal2 s 207190 219200 207246 220000 6 io_out[35]
port 105 nsew default output
rlabel metal2 s 212986 219200 213042 220000 6 io_out[36]
port 106 nsew default output
rlabel metal2 s 218782 219200 218838 220000 6 io_out[37]
port 107 nsew default output
rlabel metal2 s 21902 219200 21958 220000 6 io_out[3]
port 108 nsew default output
rlabel metal2 s 27698 219200 27754 220000 6 io_out[4]
port 109 nsew default output
rlabel metal2 s 33494 219200 33550 220000 6 io_out[5]
port 110 nsew default output
rlabel metal2 s 39290 219200 39346 220000 6 io_out[6]
port 111 nsew default output
rlabel metal2 s 45086 219200 45142 220000 6 io_out[7]
port 112 nsew default output
rlabel metal2 s 50882 219200 50938 220000 6 io_out[8]
port 113 nsew default output
rlabel metal2 s 56678 219200 56734 220000 6 io_out[9]
port 114 nsew default output
rlabel metal2 s 47570 0 47626 800 6 la_data_in[0]
port 115 nsew default input
rlabel metal2 s 182258 0 182314 800 6 la_data_in[100]
port 116 nsew default input
rlabel metal2 s 183546 0 183602 800 6 la_data_in[101]
port 117 nsew default input
rlabel metal2 s 184926 0 184982 800 6 la_data_in[102]
port 118 nsew default input
rlabel metal2 s 186306 0 186362 800 6 la_data_in[103]
port 119 nsew default input
rlabel metal2 s 187594 0 187650 800 6 la_data_in[104]
port 120 nsew default input
rlabel metal2 s 188974 0 189030 800 6 la_data_in[105]
port 121 nsew default input
rlabel metal2 s 190262 0 190318 800 6 la_data_in[106]
port 122 nsew default input
rlabel metal2 s 191642 0 191698 800 6 la_data_in[107]
port 123 nsew default input
rlabel metal2 s 193022 0 193078 800 6 la_data_in[108]
port 124 nsew default input
rlabel metal2 s 194310 0 194366 800 6 la_data_in[109]
port 125 nsew default input
rlabel metal2 s 61002 0 61058 800 6 la_data_in[10]
port 126 nsew default input
rlabel metal2 s 195690 0 195746 800 6 la_data_in[110]
port 127 nsew default input
rlabel metal2 s 197070 0 197126 800 6 la_data_in[111]
port 128 nsew default input
rlabel metal2 s 198358 0 198414 800 6 la_data_in[112]
port 129 nsew default input
rlabel metal2 s 199738 0 199794 800 6 la_data_in[113]
port 130 nsew default input
rlabel metal2 s 201118 0 201174 800 6 la_data_in[114]
port 131 nsew default input
rlabel metal2 s 202406 0 202462 800 6 la_data_in[115]
port 132 nsew default input
rlabel metal2 s 203786 0 203842 800 6 la_data_in[116]
port 133 nsew default input
rlabel metal2 s 205074 0 205130 800 6 la_data_in[117]
port 134 nsew default input
rlabel metal2 s 206454 0 206510 800 6 la_data_in[118]
port 135 nsew default input
rlabel metal2 s 207834 0 207890 800 6 la_data_in[119]
port 136 nsew default input
rlabel metal2 s 62382 0 62438 800 6 la_data_in[11]
port 137 nsew default input
rlabel metal2 s 209122 0 209178 800 6 la_data_in[120]
port 138 nsew default input
rlabel metal2 s 210502 0 210558 800 6 la_data_in[121]
port 139 nsew default input
rlabel metal2 s 211882 0 211938 800 6 la_data_in[122]
port 140 nsew default input
rlabel metal2 s 213170 0 213226 800 6 la_data_in[123]
port 141 nsew default input
rlabel metal2 s 214550 0 214606 800 6 la_data_in[124]
port 142 nsew default input
rlabel metal2 s 215930 0 215986 800 6 la_data_in[125]
port 143 nsew default input
rlabel metal2 s 217218 0 217274 800 6 la_data_in[126]
port 144 nsew default input
rlabel metal2 s 218598 0 218654 800 6 la_data_in[127]
port 145 nsew default input
rlabel metal2 s 63670 0 63726 800 6 la_data_in[12]
port 146 nsew default input
rlabel metal2 s 65050 0 65106 800 6 la_data_in[13]
port 147 nsew default input
rlabel metal2 s 66430 0 66486 800 6 la_data_in[14]
port 148 nsew default input
rlabel metal2 s 67718 0 67774 800 6 la_data_in[15]
port 149 nsew default input
rlabel metal2 s 69098 0 69154 800 6 la_data_in[16]
port 150 nsew default input
rlabel metal2 s 70478 0 70534 800 6 la_data_in[17]
port 151 nsew default input
rlabel metal2 s 71766 0 71822 800 6 la_data_in[18]
port 152 nsew default input
rlabel metal2 s 73146 0 73202 800 6 la_data_in[19]
port 153 nsew default input
rlabel metal2 s 48858 0 48914 800 6 la_data_in[1]
port 154 nsew default input
rlabel metal2 s 74526 0 74582 800 6 la_data_in[20]
port 155 nsew default input
rlabel metal2 s 75814 0 75870 800 6 la_data_in[21]
port 156 nsew default input
rlabel metal2 s 77194 0 77250 800 6 la_data_in[22]
port 157 nsew default input
rlabel metal2 s 78482 0 78538 800 6 la_data_in[23]
port 158 nsew default input
rlabel metal2 s 79862 0 79918 800 6 la_data_in[24]
port 159 nsew default input
rlabel metal2 s 81242 0 81298 800 6 la_data_in[25]
port 160 nsew default input
rlabel metal2 s 82530 0 82586 800 6 la_data_in[26]
port 161 nsew default input
rlabel metal2 s 83910 0 83966 800 6 la_data_in[27]
port 162 nsew default input
rlabel metal2 s 85290 0 85346 800 6 la_data_in[28]
port 163 nsew default input
rlabel metal2 s 86578 0 86634 800 6 la_data_in[29]
port 164 nsew default input
rlabel metal2 s 50238 0 50294 800 6 la_data_in[2]
port 165 nsew default input
rlabel metal2 s 87958 0 88014 800 6 la_data_in[30]
port 166 nsew default input
rlabel metal2 s 89338 0 89394 800 6 la_data_in[31]
port 167 nsew default input
rlabel metal2 s 90626 0 90682 800 6 la_data_in[32]
port 168 nsew default input
rlabel metal2 s 92006 0 92062 800 6 la_data_in[33]
port 169 nsew default input
rlabel metal2 s 93294 0 93350 800 6 la_data_in[34]
port 170 nsew default input
rlabel metal2 s 94674 0 94730 800 6 la_data_in[35]
port 171 nsew default input
rlabel metal2 s 96054 0 96110 800 6 la_data_in[36]
port 172 nsew default input
rlabel metal2 s 97342 0 97398 800 6 la_data_in[37]
port 173 nsew default input
rlabel metal2 s 98722 0 98778 800 6 la_data_in[38]
port 174 nsew default input
rlabel metal2 s 100102 0 100158 800 6 la_data_in[39]
port 175 nsew default input
rlabel metal2 s 51618 0 51674 800 6 la_data_in[3]
port 176 nsew default input
rlabel metal2 s 101390 0 101446 800 6 la_data_in[40]
port 177 nsew default input
rlabel metal2 s 102770 0 102826 800 6 la_data_in[41]
port 178 nsew default input
rlabel metal2 s 104150 0 104206 800 6 la_data_in[42]
port 179 nsew default input
rlabel metal2 s 105438 0 105494 800 6 la_data_in[43]
port 180 nsew default input
rlabel metal2 s 106818 0 106874 800 6 la_data_in[44]
port 181 nsew default input
rlabel metal2 s 108106 0 108162 800 6 la_data_in[45]
port 182 nsew default input
rlabel metal2 s 109486 0 109542 800 6 la_data_in[46]
port 183 nsew default input
rlabel metal2 s 110866 0 110922 800 6 la_data_in[47]
port 184 nsew default input
rlabel metal2 s 112154 0 112210 800 6 la_data_in[48]
port 185 nsew default input
rlabel metal2 s 113534 0 113590 800 6 la_data_in[49]
port 186 nsew default input
rlabel metal2 s 52906 0 52962 800 6 la_data_in[4]
port 187 nsew default input
rlabel metal2 s 114914 0 114970 800 6 la_data_in[50]
port 188 nsew default input
rlabel metal2 s 116202 0 116258 800 6 la_data_in[51]
port 189 nsew default input
rlabel metal2 s 117582 0 117638 800 6 la_data_in[52]
port 190 nsew default input
rlabel metal2 s 118962 0 119018 800 6 la_data_in[53]
port 191 nsew default input
rlabel metal2 s 120250 0 120306 800 6 la_data_in[54]
port 192 nsew default input
rlabel metal2 s 121630 0 121686 800 6 la_data_in[55]
port 193 nsew default input
rlabel metal2 s 123010 0 123066 800 6 la_data_in[56]
port 194 nsew default input
rlabel metal2 s 124298 0 124354 800 6 la_data_in[57]
port 195 nsew default input
rlabel metal2 s 125678 0 125734 800 6 la_data_in[58]
port 196 nsew default input
rlabel metal2 s 126966 0 127022 800 6 la_data_in[59]
port 197 nsew default input
rlabel metal2 s 54286 0 54342 800 6 la_data_in[5]
port 198 nsew default input
rlabel metal2 s 128346 0 128402 800 6 la_data_in[60]
port 199 nsew default input
rlabel metal2 s 129726 0 129782 800 6 la_data_in[61]
port 200 nsew default input
rlabel metal2 s 131014 0 131070 800 6 la_data_in[62]
port 201 nsew default input
rlabel metal2 s 132394 0 132450 800 6 la_data_in[63]
port 202 nsew default input
rlabel metal2 s 133774 0 133830 800 6 la_data_in[64]
port 203 nsew default input
rlabel metal2 s 135062 0 135118 800 6 la_data_in[65]
port 204 nsew default input
rlabel metal2 s 136442 0 136498 800 6 la_data_in[66]
port 205 nsew default input
rlabel metal2 s 137822 0 137878 800 6 la_data_in[67]
port 206 nsew default input
rlabel metal2 s 139110 0 139166 800 6 la_data_in[68]
port 207 nsew default input
rlabel metal2 s 140490 0 140546 800 6 la_data_in[69]
port 208 nsew default input
rlabel metal2 s 55666 0 55722 800 6 la_data_in[6]
port 209 nsew default input
rlabel metal2 s 141778 0 141834 800 6 la_data_in[70]
port 210 nsew default input
rlabel metal2 s 143158 0 143214 800 6 la_data_in[71]
port 211 nsew default input
rlabel metal2 s 144538 0 144594 800 6 la_data_in[72]
port 212 nsew default input
rlabel metal2 s 145826 0 145882 800 6 la_data_in[73]
port 213 nsew default input
rlabel metal2 s 147206 0 147262 800 6 la_data_in[74]
port 214 nsew default input
rlabel metal2 s 148586 0 148642 800 6 la_data_in[75]
port 215 nsew default input
rlabel metal2 s 149874 0 149930 800 6 la_data_in[76]
port 216 nsew default input
rlabel metal2 s 151254 0 151310 800 6 la_data_in[77]
port 217 nsew default input
rlabel metal2 s 152634 0 152690 800 6 la_data_in[78]
port 218 nsew default input
rlabel metal2 s 153922 0 153978 800 6 la_data_in[79]
port 219 nsew default input
rlabel metal2 s 56954 0 57010 800 6 la_data_in[7]
port 220 nsew default input
rlabel metal2 s 155302 0 155358 800 6 la_data_in[80]
port 221 nsew default input
rlabel metal2 s 156590 0 156646 800 6 la_data_in[81]
port 222 nsew default input
rlabel metal2 s 157970 0 158026 800 6 la_data_in[82]
port 223 nsew default input
rlabel metal2 s 159350 0 159406 800 6 la_data_in[83]
port 224 nsew default input
rlabel metal2 s 160638 0 160694 800 6 la_data_in[84]
port 225 nsew default input
rlabel metal2 s 162018 0 162074 800 6 la_data_in[85]
port 226 nsew default input
rlabel metal2 s 163398 0 163454 800 6 la_data_in[86]
port 227 nsew default input
rlabel metal2 s 164686 0 164742 800 6 la_data_in[87]
port 228 nsew default input
rlabel metal2 s 166066 0 166122 800 6 la_data_in[88]
port 229 nsew default input
rlabel metal2 s 167446 0 167502 800 6 la_data_in[89]
port 230 nsew default input
rlabel metal2 s 58334 0 58390 800 6 la_data_in[8]
port 231 nsew default input
rlabel metal2 s 168734 0 168790 800 6 la_data_in[90]
port 232 nsew default input
rlabel metal2 s 170114 0 170170 800 6 la_data_in[91]
port 233 nsew default input
rlabel metal2 s 171494 0 171550 800 6 la_data_in[92]
port 234 nsew default input
rlabel metal2 s 172782 0 172838 800 6 la_data_in[93]
port 235 nsew default input
rlabel metal2 s 174162 0 174218 800 6 la_data_in[94]
port 236 nsew default input
rlabel metal2 s 175450 0 175506 800 6 la_data_in[95]
port 237 nsew default input
rlabel metal2 s 176830 0 176886 800 6 la_data_in[96]
port 238 nsew default input
rlabel metal2 s 178210 0 178266 800 6 la_data_in[97]
port 239 nsew default input
rlabel metal2 s 179498 0 179554 800 6 la_data_in[98]
port 240 nsew default input
rlabel metal2 s 180878 0 180934 800 6 la_data_in[99]
port 241 nsew default input
rlabel metal2 s 59622 0 59678 800 6 la_data_in[9]
port 242 nsew default input
rlabel metal2 s 48030 0 48086 800 6 la_data_out[0]
port 243 nsew default output
rlabel metal2 s 182626 0 182682 800 6 la_data_out[100]
port 244 nsew default output
rlabel metal2 s 184006 0 184062 800 6 la_data_out[101]
port 245 nsew default output
rlabel metal2 s 185386 0 185442 800 6 la_data_out[102]
port 246 nsew default output
rlabel metal2 s 186674 0 186730 800 6 la_data_out[103]
port 247 nsew default output
rlabel metal2 s 188054 0 188110 800 6 la_data_out[104]
port 248 nsew default output
rlabel metal2 s 189434 0 189490 800 6 la_data_out[105]
port 249 nsew default output
rlabel metal2 s 190722 0 190778 800 6 la_data_out[106]
port 250 nsew default output
rlabel metal2 s 192102 0 192158 800 6 la_data_out[107]
port 251 nsew default output
rlabel metal2 s 193482 0 193538 800 6 la_data_out[108]
port 252 nsew default output
rlabel metal2 s 194770 0 194826 800 6 la_data_out[109]
port 253 nsew default output
rlabel metal2 s 61462 0 61518 800 6 la_data_out[10]
port 254 nsew default output
rlabel metal2 s 196150 0 196206 800 6 la_data_out[110]
port 255 nsew default output
rlabel metal2 s 197530 0 197586 800 6 la_data_out[111]
port 256 nsew default output
rlabel metal2 s 198818 0 198874 800 6 la_data_out[112]
port 257 nsew default output
rlabel metal2 s 200198 0 200254 800 6 la_data_out[113]
port 258 nsew default output
rlabel metal2 s 201486 0 201542 800 6 la_data_out[114]
port 259 nsew default output
rlabel metal2 s 202866 0 202922 800 6 la_data_out[115]
port 260 nsew default output
rlabel metal2 s 204246 0 204302 800 6 la_data_out[116]
port 261 nsew default output
rlabel metal2 s 205534 0 205590 800 6 la_data_out[117]
port 262 nsew default output
rlabel metal2 s 206914 0 206970 800 6 la_data_out[118]
port 263 nsew default output
rlabel metal2 s 208294 0 208350 800 6 la_data_out[119]
port 264 nsew default output
rlabel metal2 s 62842 0 62898 800 6 la_data_out[11]
port 265 nsew default output
rlabel metal2 s 209582 0 209638 800 6 la_data_out[120]
port 266 nsew default output
rlabel metal2 s 210962 0 211018 800 6 la_data_out[121]
port 267 nsew default output
rlabel metal2 s 212342 0 212398 800 6 la_data_out[122]
port 268 nsew default output
rlabel metal2 s 213630 0 213686 800 6 la_data_out[123]
port 269 nsew default output
rlabel metal2 s 215010 0 215066 800 6 la_data_out[124]
port 270 nsew default output
rlabel metal2 s 216298 0 216354 800 6 la_data_out[125]
port 271 nsew default output
rlabel metal2 s 217678 0 217734 800 6 la_data_out[126]
port 272 nsew default output
rlabel metal2 s 219058 0 219114 800 6 la_data_out[127]
port 273 nsew default output
rlabel metal2 s 64130 0 64186 800 6 la_data_out[12]
port 274 nsew default output
rlabel metal2 s 65510 0 65566 800 6 la_data_out[13]
port 275 nsew default output
rlabel metal2 s 66890 0 66946 800 6 la_data_out[14]
port 276 nsew default output
rlabel metal2 s 68178 0 68234 800 6 la_data_out[15]
port 277 nsew default output
rlabel metal2 s 69558 0 69614 800 6 la_data_out[16]
port 278 nsew default output
rlabel metal2 s 70846 0 70902 800 6 la_data_out[17]
port 279 nsew default output
rlabel metal2 s 72226 0 72282 800 6 la_data_out[18]
port 280 nsew default output
rlabel metal2 s 73606 0 73662 800 6 la_data_out[19]
port 281 nsew default output
rlabel metal2 s 49318 0 49374 800 6 la_data_out[1]
port 282 nsew default output
rlabel metal2 s 74894 0 74950 800 6 la_data_out[20]
port 283 nsew default output
rlabel metal2 s 76274 0 76330 800 6 la_data_out[21]
port 284 nsew default output
rlabel metal2 s 77654 0 77710 800 6 la_data_out[22]
port 285 nsew default output
rlabel metal2 s 78942 0 78998 800 6 la_data_out[23]
port 286 nsew default output
rlabel metal2 s 80322 0 80378 800 6 la_data_out[24]
port 287 nsew default output
rlabel metal2 s 81702 0 81758 800 6 la_data_out[25]
port 288 nsew default output
rlabel metal2 s 82990 0 83046 800 6 la_data_out[26]
port 289 nsew default output
rlabel metal2 s 84370 0 84426 800 6 la_data_out[27]
port 290 nsew default output
rlabel metal2 s 85750 0 85806 800 6 la_data_out[28]
port 291 nsew default output
rlabel metal2 s 87038 0 87094 800 6 la_data_out[29]
port 292 nsew default output
rlabel metal2 s 50698 0 50754 800 6 la_data_out[2]
port 293 nsew default output
rlabel metal2 s 88418 0 88474 800 6 la_data_out[30]
port 294 nsew default output
rlabel metal2 s 89706 0 89762 800 6 la_data_out[31]
port 295 nsew default output
rlabel metal2 s 91086 0 91142 800 6 la_data_out[32]
port 296 nsew default output
rlabel metal2 s 92466 0 92522 800 6 la_data_out[33]
port 297 nsew default output
rlabel metal2 s 93754 0 93810 800 6 la_data_out[34]
port 298 nsew default output
rlabel metal2 s 95134 0 95190 800 6 la_data_out[35]
port 299 nsew default output
rlabel metal2 s 96514 0 96570 800 6 la_data_out[36]
port 300 nsew default output
rlabel metal2 s 97802 0 97858 800 6 la_data_out[37]
port 301 nsew default output
rlabel metal2 s 99182 0 99238 800 6 la_data_out[38]
port 302 nsew default output
rlabel metal2 s 100562 0 100618 800 6 la_data_out[39]
port 303 nsew default output
rlabel metal2 s 52078 0 52134 800 6 la_data_out[3]
port 304 nsew default output
rlabel metal2 s 101850 0 101906 800 6 la_data_out[40]
port 305 nsew default output
rlabel metal2 s 103230 0 103286 800 6 la_data_out[41]
port 306 nsew default output
rlabel metal2 s 104518 0 104574 800 6 la_data_out[42]
port 307 nsew default output
rlabel metal2 s 105898 0 105954 800 6 la_data_out[43]
port 308 nsew default output
rlabel metal2 s 107278 0 107334 800 6 la_data_out[44]
port 309 nsew default output
rlabel metal2 s 108566 0 108622 800 6 la_data_out[45]
port 310 nsew default output
rlabel metal2 s 109946 0 110002 800 6 la_data_out[46]
port 311 nsew default output
rlabel metal2 s 111326 0 111382 800 6 la_data_out[47]
port 312 nsew default output
rlabel metal2 s 112614 0 112670 800 6 la_data_out[48]
port 313 nsew default output
rlabel metal2 s 113994 0 114050 800 6 la_data_out[49]
port 314 nsew default output
rlabel metal2 s 53366 0 53422 800 6 la_data_out[4]
port 315 nsew default output
rlabel metal2 s 115374 0 115430 800 6 la_data_out[50]
port 316 nsew default output
rlabel metal2 s 116662 0 116718 800 6 la_data_out[51]
port 317 nsew default output
rlabel metal2 s 118042 0 118098 800 6 la_data_out[52]
port 318 nsew default output
rlabel metal2 s 119330 0 119386 800 6 la_data_out[53]
port 319 nsew default output
rlabel metal2 s 120710 0 120766 800 6 la_data_out[54]
port 320 nsew default output
rlabel metal2 s 122090 0 122146 800 6 la_data_out[55]
port 321 nsew default output
rlabel metal2 s 123378 0 123434 800 6 la_data_out[56]
port 322 nsew default output
rlabel metal2 s 124758 0 124814 800 6 la_data_out[57]
port 323 nsew default output
rlabel metal2 s 126138 0 126194 800 6 la_data_out[58]
port 324 nsew default output
rlabel metal2 s 127426 0 127482 800 6 la_data_out[59]
port 325 nsew default output
rlabel metal2 s 54746 0 54802 800 6 la_data_out[5]
port 326 nsew default output
rlabel metal2 s 128806 0 128862 800 6 la_data_out[60]
port 327 nsew default output
rlabel metal2 s 130186 0 130242 800 6 la_data_out[61]
port 328 nsew default output
rlabel metal2 s 131474 0 131530 800 6 la_data_out[62]
port 329 nsew default output
rlabel metal2 s 132854 0 132910 800 6 la_data_out[63]
port 330 nsew default output
rlabel metal2 s 134142 0 134198 800 6 la_data_out[64]
port 331 nsew default output
rlabel metal2 s 135522 0 135578 800 6 la_data_out[65]
port 332 nsew default output
rlabel metal2 s 136902 0 136958 800 6 la_data_out[66]
port 333 nsew default output
rlabel metal2 s 138190 0 138246 800 6 la_data_out[67]
port 334 nsew default output
rlabel metal2 s 139570 0 139626 800 6 la_data_out[68]
port 335 nsew default output
rlabel metal2 s 140950 0 141006 800 6 la_data_out[69]
port 336 nsew default output
rlabel metal2 s 56034 0 56090 800 6 la_data_out[6]
port 337 nsew default output
rlabel metal2 s 142238 0 142294 800 6 la_data_out[70]
port 338 nsew default output
rlabel metal2 s 143618 0 143674 800 6 la_data_out[71]
port 339 nsew default output
rlabel metal2 s 144998 0 145054 800 6 la_data_out[72]
port 340 nsew default output
rlabel metal2 s 146286 0 146342 800 6 la_data_out[73]
port 341 nsew default output
rlabel metal2 s 147666 0 147722 800 6 la_data_out[74]
port 342 nsew default output
rlabel metal2 s 149046 0 149102 800 6 la_data_out[75]
port 343 nsew default output
rlabel metal2 s 150334 0 150390 800 6 la_data_out[76]
port 344 nsew default output
rlabel metal2 s 151714 0 151770 800 6 la_data_out[77]
port 345 nsew default output
rlabel metal2 s 153002 0 153058 800 6 la_data_out[78]
port 346 nsew default output
rlabel metal2 s 154382 0 154438 800 6 la_data_out[79]
port 347 nsew default output
rlabel metal2 s 57414 0 57470 800 6 la_data_out[7]
port 348 nsew default output
rlabel metal2 s 155762 0 155818 800 6 la_data_out[80]
port 349 nsew default output
rlabel metal2 s 157050 0 157106 800 6 la_data_out[81]
port 350 nsew default output
rlabel metal2 s 158430 0 158486 800 6 la_data_out[82]
port 351 nsew default output
rlabel metal2 s 159810 0 159866 800 6 la_data_out[83]
port 352 nsew default output
rlabel metal2 s 161098 0 161154 800 6 la_data_out[84]
port 353 nsew default output
rlabel metal2 s 162478 0 162534 800 6 la_data_out[85]
port 354 nsew default output
rlabel metal2 s 163858 0 163914 800 6 la_data_out[86]
port 355 nsew default output
rlabel metal2 s 165146 0 165202 800 6 la_data_out[87]
port 356 nsew default output
rlabel metal2 s 166526 0 166582 800 6 la_data_out[88]
port 357 nsew default output
rlabel metal2 s 167814 0 167870 800 6 la_data_out[89]
port 358 nsew default output
rlabel metal2 s 58794 0 58850 800 6 la_data_out[8]
port 359 nsew default output
rlabel metal2 s 169194 0 169250 800 6 la_data_out[90]
port 360 nsew default output
rlabel metal2 s 170574 0 170630 800 6 la_data_out[91]
port 361 nsew default output
rlabel metal2 s 171862 0 171918 800 6 la_data_out[92]
port 362 nsew default output
rlabel metal2 s 173242 0 173298 800 6 la_data_out[93]
port 363 nsew default output
rlabel metal2 s 174622 0 174678 800 6 la_data_out[94]
port 364 nsew default output
rlabel metal2 s 175910 0 175966 800 6 la_data_out[95]
port 365 nsew default output
rlabel metal2 s 177290 0 177346 800 6 la_data_out[96]
port 366 nsew default output
rlabel metal2 s 178670 0 178726 800 6 la_data_out[97]
port 367 nsew default output
rlabel metal2 s 179958 0 180014 800 6 la_data_out[98]
port 368 nsew default output
rlabel metal2 s 181338 0 181394 800 6 la_data_out[99]
port 369 nsew default output
rlabel metal2 s 60082 0 60138 800 6 la_data_out[9]
port 370 nsew default output
rlabel metal2 s 48398 0 48454 800 6 la_oen[0]
port 371 nsew default input
rlabel metal2 s 183086 0 183142 800 6 la_oen[100]
port 372 nsew default input
rlabel metal2 s 184466 0 184522 800 6 la_oen[101]
port 373 nsew default input
rlabel metal2 s 185846 0 185902 800 6 la_oen[102]
port 374 nsew default input
rlabel metal2 s 187134 0 187190 800 6 la_oen[103]
port 375 nsew default input
rlabel metal2 s 188514 0 188570 800 6 la_oen[104]
port 376 nsew default input
rlabel metal2 s 189894 0 189950 800 6 la_oen[105]
port 377 nsew default input
rlabel metal2 s 191182 0 191238 800 6 la_oen[106]
port 378 nsew default input
rlabel metal2 s 192562 0 192618 800 6 la_oen[107]
port 379 nsew default input
rlabel metal2 s 193850 0 193906 800 6 la_oen[108]
port 380 nsew default input
rlabel metal2 s 195230 0 195286 800 6 la_oen[109]
port 381 nsew default input
rlabel metal2 s 61922 0 61978 800 6 la_oen[10]
port 382 nsew default input
rlabel metal2 s 196610 0 196666 800 6 la_oen[110]
port 383 nsew default input
rlabel metal2 s 197898 0 197954 800 6 la_oen[111]
port 384 nsew default input
rlabel metal2 s 199278 0 199334 800 6 la_oen[112]
port 385 nsew default input
rlabel metal2 s 200658 0 200714 800 6 la_oen[113]
port 386 nsew default input
rlabel metal2 s 201946 0 202002 800 6 la_oen[114]
port 387 nsew default input
rlabel metal2 s 203326 0 203382 800 6 la_oen[115]
port 388 nsew default input
rlabel metal2 s 204706 0 204762 800 6 la_oen[116]
port 389 nsew default input
rlabel metal2 s 205994 0 206050 800 6 la_oen[117]
port 390 nsew default input
rlabel metal2 s 207374 0 207430 800 6 la_oen[118]
port 391 nsew default input
rlabel metal2 s 208754 0 208810 800 6 la_oen[119]
port 392 nsew default input
rlabel metal2 s 63302 0 63358 800 6 la_oen[11]
port 393 nsew default input
rlabel metal2 s 210042 0 210098 800 6 la_oen[120]
port 394 nsew default input
rlabel metal2 s 211422 0 211478 800 6 la_oen[121]
port 395 nsew default input
rlabel metal2 s 212710 0 212766 800 6 la_oen[122]
port 396 nsew default input
rlabel metal2 s 214090 0 214146 800 6 la_oen[123]
port 397 nsew default input
rlabel metal2 s 215470 0 215526 800 6 la_oen[124]
port 398 nsew default input
rlabel metal2 s 216758 0 216814 800 6 la_oen[125]
port 399 nsew default input
rlabel metal2 s 218138 0 218194 800 6 la_oen[126]
port 400 nsew default input
rlabel metal2 s 219518 0 219574 800 6 la_oen[127]
port 401 nsew default input
rlabel metal2 s 64590 0 64646 800 6 la_oen[12]
port 402 nsew default input
rlabel metal2 s 65970 0 66026 800 6 la_oen[13]
port 403 nsew default input
rlabel metal2 s 67258 0 67314 800 6 la_oen[14]
port 404 nsew default input
rlabel metal2 s 68638 0 68694 800 6 la_oen[15]
port 405 nsew default input
rlabel metal2 s 70018 0 70074 800 6 la_oen[16]
port 406 nsew default input
rlabel metal2 s 71306 0 71362 800 6 la_oen[17]
port 407 nsew default input
rlabel metal2 s 72686 0 72742 800 6 la_oen[18]
port 408 nsew default input
rlabel metal2 s 74066 0 74122 800 6 la_oen[19]
port 409 nsew default input
rlabel metal2 s 49778 0 49834 800 6 la_oen[1]
port 410 nsew default input
rlabel metal2 s 75354 0 75410 800 6 la_oen[20]
port 411 nsew default input
rlabel metal2 s 76734 0 76790 800 6 la_oen[21]
port 412 nsew default input
rlabel metal2 s 78114 0 78170 800 6 la_oen[22]
port 413 nsew default input
rlabel metal2 s 79402 0 79458 800 6 la_oen[23]
port 414 nsew default input
rlabel metal2 s 80782 0 80838 800 6 la_oen[24]
port 415 nsew default input
rlabel metal2 s 82070 0 82126 800 6 la_oen[25]
port 416 nsew default input
rlabel metal2 s 83450 0 83506 800 6 la_oen[26]
port 417 nsew default input
rlabel metal2 s 84830 0 84886 800 6 la_oen[27]
port 418 nsew default input
rlabel metal2 s 86118 0 86174 800 6 la_oen[28]
port 419 nsew default input
rlabel metal2 s 87498 0 87554 800 6 la_oen[29]
port 420 nsew default input
rlabel metal2 s 51158 0 51214 800 6 la_oen[2]
port 421 nsew default input
rlabel metal2 s 88878 0 88934 800 6 la_oen[30]
port 422 nsew default input
rlabel metal2 s 90166 0 90222 800 6 la_oen[31]
port 423 nsew default input
rlabel metal2 s 91546 0 91602 800 6 la_oen[32]
port 424 nsew default input
rlabel metal2 s 92926 0 92982 800 6 la_oen[33]
port 425 nsew default input
rlabel metal2 s 94214 0 94270 800 6 la_oen[34]
port 426 nsew default input
rlabel metal2 s 95594 0 95650 800 6 la_oen[35]
port 427 nsew default input
rlabel metal2 s 96882 0 96938 800 6 la_oen[36]
port 428 nsew default input
rlabel metal2 s 98262 0 98318 800 6 la_oen[37]
port 429 nsew default input
rlabel metal2 s 99642 0 99698 800 6 la_oen[38]
port 430 nsew default input
rlabel metal2 s 100930 0 100986 800 6 la_oen[39]
port 431 nsew default input
rlabel metal2 s 52446 0 52502 800 6 la_oen[3]
port 432 nsew default input
rlabel metal2 s 102310 0 102366 800 6 la_oen[40]
port 433 nsew default input
rlabel metal2 s 103690 0 103746 800 6 la_oen[41]
port 434 nsew default input
rlabel metal2 s 104978 0 105034 800 6 la_oen[42]
port 435 nsew default input
rlabel metal2 s 106358 0 106414 800 6 la_oen[43]
port 436 nsew default input
rlabel metal2 s 107738 0 107794 800 6 la_oen[44]
port 437 nsew default input
rlabel metal2 s 109026 0 109082 800 6 la_oen[45]
port 438 nsew default input
rlabel metal2 s 110406 0 110462 800 6 la_oen[46]
port 439 nsew default input
rlabel metal2 s 111786 0 111842 800 6 la_oen[47]
port 440 nsew default input
rlabel metal2 s 113074 0 113130 800 6 la_oen[48]
port 441 nsew default input
rlabel metal2 s 114454 0 114510 800 6 la_oen[49]
port 442 nsew default input
rlabel metal2 s 53826 0 53882 800 6 la_oen[4]
port 443 nsew default input
rlabel metal2 s 115742 0 115798 800 6 la_oen[50]
port 444 nsew default input
rlabel metal2 s 117122 0 117178 800 6 la_oen[51]
port 445 nsew default input
rlabel metal2 s 118502 0 118558 800 6 la_oen[52]
port 446 nsew default input
rlabel metal2 s 119790 0 119846 800 6 la_oen[53]
port 447 nsew default input
rlabel metal2 s 121170 0 121226 800 6 la_oen[54]
port 448 nsew default input
rlabel metal2 s 122550 0 122606 800 6 la_oen[55]
port 449 nsew default input
rlabel metal2 s 123838 0 123894 800 6 la_oen[56]
port 450 nsew default input
rlabel metal2 s 125218 0 125274 800 6 la_oen[57]
port 451 nsew default input
rlabel metal2 s 126598 0 126654 800 6 la_oen[58]
port 452 nsew default input
rlabel metal2 s 127886 0 127942 800 6 la_oen[59]
port 453 nsew default input
rlabel metal2 s 55206 0 55262 800 6 la_oen[5]
port 454 nsew default input
rlabel metal2 s 129266 0 129322 800 6 la_oen[60]
port 455 nsew default input
rlabel metal2 s 130554 0 130610 800 6 la_oen[61]
port 456 nsew default input
rlabel metal2 s 131934 0 131990 800 6 la_oen[62]
port 457 nsew default input
rlabel metal2 s 133314 0 133370 800 6 la_oen[63]
port 458 nsew default input
rlabel metal2 s 134602 0 134658 800 6 la_oen[64]
port 459 nsew default input
rlabel metal2 s 135982 0 136038 800 6 la_oen[65]
port 460 nsew default input
rlabel metal2 s 137362 0 137418 800 6 la_oen[66]
port 461 nsew default input
rlabel metal2 s 138650 0 138706 800 6 la_oen[67]
port 462 nsew default input
rlabel metal2 s 140030 0 140086 800 6 la_oen[68]
port 463 nsew default input
rlabel metal2 s 141410 0 141466 800 6 la_oen[69]
port 464 nsew default input
rlabel metal2 s 56494 0 56550 800 6 la_oen[6]
port 465 nsew default input
rlabel metal2 s 142698 0 142754 800 6 la_oen[70]
port 466 nsew default input
rlabel metal2 s 144078 0 144134 800 6 la_oen[71]
port 467 nsew default input
rlabel metal2 s 145366 0 145422 800 6 la_oen[72]
port 468 nsew default input
rlabel metal2 s 146746 0 146802 800 6 la_oen[73]
port 469 nsew default input
rlabel metal2 s 148126 0 148182 800 6 la_oen[74]
port 470 nsew default input
rlabel metal2 s 149414 0 149470 800 6 la_oen[75]
port 471 nsew default input
rlabel metal2 s 150794 0 150850 800 6 la_oen[76]
port 472 nsew default input
rlabel metal2 s 152174 0 152230 800 6 la_oen[77]
port 473 nsew default input
rlabel metal2 s 153462 0 153518 800 6 la_oen[78]
port 474 nsew default input
rlabel metal2 s 154842 0 154898 800 6 la_oen[79]
port 475 nsew default input
rlabel metal2 s 57874 0 57930 800 6 la_oen[7]
port 476 nsew default input
rlabel metal2 s 156222 0 156278 800 6 la_oen[80]
port 477 nsew default input
rlabel metal2 s 157510 0 157566 800 6 la_oen[81]
port 478 nsew default input
rlabel metal2 s 158890 0 158946 800 6 la_oen[82]
port 479 nsew default input
rlabel metal2 s 160270 0 160326 800 6 la_oen[83]
port 480 nsew default input
rlabel metal2 s 161558 0 161614 800 6 la_oen[84]
port 481 nsew default input
rlabel metal2 s 162938 0 162994 800 6 la_oen[85]
port 482 nsew default input
rlabel metal2 s 164226 0 164282 800 6 la_oen[86]
port 483 nsew default input
rlabel metal2 s 165606 0 165662 800 6 la_oen[87]
port 484 nsew default input
rlabel metal2 s 166986 0 167042 800 6 la_oen[88]
port 485 nsew default input
rlabel metal2 s 168274 0 168330 800 6 la_oen[89]
port 486 nsew default input
rlabel metal2 s 59254 0 59310 800 6 la_oen[8]
port 487 nsew default input
rlabel metal2 s 169654 0 169710 800 6 la_oen[90]
port 488 nsew default input
rlabel metal2 s 171034 0 171090 800 6 la_oen[91]
port 489 nsew default input
rlabel metal2 s 172322 0 172378 800 6 la_oen[92]
port 490 nsew default input
rlabel metal2 s 173702 0 173758 800 6 la_oen[93]
port 491 nsew default input
rlabel metal2 s 175082 0 175138 800 6 la_oen[94]
port 492 nsew default input
rlabel metal2 s 176370 0 176426 800 6 la_oen[95]
port 493 nsew default input
rlabel metal2 s 177750 0 177806 800 6 la_oen[96]
port 494 nsew default input
rlabel metal2 s 179038 0 179094 800 6 la_oen[97]
port 495 nsew default input
rlabel metal2 s 180418 0 180474 800 6 la_oen[98]
port 496 nsew default input
rlabel metal2 s 181798 0 181854 800 6 la_oen[99]
port 497 nsew default input
rlabel metal2 s 60542 0 60598 800 6 la_oen[9]
port 498 nsew default input
rlabel metal2 s 6 0 62 800 6 wb_clk_i
port 499 nsew default input
rlabel metal2 s 374 0 430 800 6 wb_rst_i
port 500 nsew default input
rlabel metal2 s 834 0 890 800 6 wbs_ack_o
port 501 nsew default output
rlabel metal2 s 2674 0 2730 800 6 wbs_adr_i[0]
port 502 nsew default input
rlabel metal2 s 17946 0 18002 800 6 wbs_adr_i[10]
port 503 nsew default input
rlabel metal2 s 19234 0 19290 800 6 wbs_adr_i[11]
port 504 nsew default input
rlabel metal2 s 20614 0 20670 800 6 wbs_adr_i[12]
port 505 nsew default input
rlabel metal2 s 21994 0 22050 800 6 wbs_adr_i[13]
port 506 nsew default input
rlabel metal2 s 23282 0 23338 800 6 wbs_adr_i[14]
port 507 nsew default input
rlabel metal2 s 24662 0 24718 800 6 wbs_adr_i[15]
port 508 nsew default input
rlabel metal2 s 26042 0 26098 800 6 wbs_adr_i[16]
port 509 nsew default input
rlabel metal2 s 27330 0 27386 800 6 wbs_adr_i[17]
port 510 nsew default input
rlabel metal2 s 28710 0 28766 800 6 wbs_adr_i[18]
port 511 nsew default input
rlabel metal2 s 29998 0 30054 800 6 wbs_adr_i[19]
port 512 nsew default input
rlabel metal2 s 4422 0 4478 800 6 wbs_adr_i[1]
port 513 nsew default input
rlabel metal2 s 31378 0 31434 800 6 wbs_adr_i[20]
port 514 nsew default input
rlabel metal2 s 32758 0 32814 800 6 wbs_adr_i[21]
port 515 nsew default input
rlabel metal2 s 34046 0 34102 800 6 wbs_adr_i[22]
port 516 nsew default input
rlabel metal2 s 35426 0 35482 800 6 wbs_adr_i[23]
port 517 nsew default input
rlabel metal2 s 36806 0 36862 800 6 wbs_adr_i[24]
port 518 nsew default input
rlabel metal2 s 38094 0 38150 800 6 wbs_adr_i[25]
port 519 nsew default input
rlabel metal2 s 39474 0 39530 800 6 wbs_adr_i[26]
port 520 nsew default input
rlabel metal2 s 40854 0 40910 800 6 wbs_adr_i[27]
port 521 nsew default input
rlabel metal2 s 42142 0 42198 800 6 wbs_adr_i[28]
port 522 nsew default input
rlabel metal2 s 43522 0 43578 800 6 wbs_adr_i[29]
port 523 nsew default input
rlabel metal2 s 6262 0 6318 800 6 wbs_adr_i[2]
port 524 nsew default input
rlabel metal2 s 44810 0 44866 800 6 wbs_adr_i[30]
port 525 nsew default input
rlabel metal2 s 46190 0 46246 800 6 wbs_adr_i[31]
port 526 nsew default input
rlabel metal2 s 8010 0 8066 800 6 wbs_adr_i[3]
port 527 nsew default input
rlabel metal2 s 9850 0 9906 800 6 wbs_adr_i[4]
port 528 nsew default input
rlabel metal2 s 11138 0 11194 800 6 wbs_adr_i[5]
port 529 nsew default input
rlabel metal2 s 12518 0 12574 800 6 wbs_adr_i[6]
port 530 nsew default input
rlabel metal2 s 13898 0 13954 800 6 wbs_adr_i[7]
port 531 nsew default input
rlabel metal2 s 15186 0 15242 800 6 wbs_adr_i[8]
port 532 nsew default input
rlabel metal2 s 16566 0 16622 800 6 wbs_adr_i[9]
port 533 nsew default input
rlabel metal2 s 1294 0 1350 800 6 wbs_cyc_i
port 534 nsew default input
rlabel metal2 s 3134 0 3190 800 6 wbs_dat_i[0]
port 535 nsew default input
rlabel metal2 s 18406 0 18462 800 6 wbs_dat_i[10]
port 536 nsew default input
rlabel metal2 s 19694 0 19750 800 6 wbs_dat_i[11]
port 537 nsew default input
rlabel metal2 s 21074 0 21130 800 6 wbs_dat_i[12]
port 538 nsew default input
rlabel metal2 s 22362 0 22418 800 6 wbs_dat_i[13]
port 539 nsew default input
rlabel metal2 s 23742 0 23798 800 6 wbs_dat_i[14]
port 540 nsew default input
rlabel metal2 s 25122 0 25178 800 6 wbs_dat_i[15]
port 541 nsew default input
rlabel metal2 s 26410 0 26466 800 6 wbs_dat_i[16]
port 542 nsew default input
rlabel metal2 s 27790 0 27846 800 6 wbs_dat_i[17]
port 543 nsew default input
rlabel metal2 s 29170 0 29226 800 6 wbs_dat_i[18]
port 544 nsew default input
rlabel metal2 s 30458 0 30514 800 6 wbs_dat_i[19]
port 545 nsew default input
rlabel metal2 s 4882 0 4938 800 6 wbs_dat_i[1]
port 546 nsew default input
rlabel metal2 s 31838 0 31894 800 6 wbs_dat_i[20]
port 547 nsew default input
rlabel metal2 s 33218 0 33274 800 6 wbs_dat_i[21]
port 548 nsew default input
rlabel metal2 s 34506 0 34562 800 6 wbs_dat_i[22]
port 549 nsew default input
rlabel metal2 s 35886 0 35942 800 6 wbs_dat_i[23]
port 550 nsew default input
rlabel metal2 s 37266 0 37322 800 6 wbs_dat_i[24]
port 551 nsew default input
rlabel metal2 s 38554 0 38610 800 6 wbs_dat_i[25]
port 552 nsew default input
rlabel metal2 s 39934 0 39990 800 6 wbs_dat_i[26]
port 553 nsew default input
rlabel metal2 s 41222 0 41278 800 6 wbs_dat_i[27]
port 554 nsew default input
rlabel metal2 s 42602 0 42658 800 6 wbs_dat_i[28]
port 555 nsew default input
rlabel metal2 s 43982 0 44038 800 6 wbs_dat_i[29]
port 556 nsew default input
rlabel metal2 s 6722 0 6778 800 6 wbs_dat_i[2]
port 557 nsew default input
rlabel metal2 s 45270 0 45326 800 6 wbs_dat_i[30]
port 558 nsew default input
rlabel metal2 s 46650 0 46706 800 6 wbs_dat_i[31]
port 559 nsew default input
rlabel metal2 s 8470 0 8526 800 6 wbs_dat_i[3]
port 560 nsew default input
rlabel metal2 s 10310 0 10366 800 6 wbs_dat_i[4]
port 561 nsew default input
rlabel metal2 s 11598 0 11654 800 6 wbs_dat_i[5]
port 562 nsew default input
rlabel metal2 s 12978 0 13034 800 6 wbs_dat_i[6]
port 563 nsew default input
rlabel metal2 s 14358 0 14414 800 6 wbs_dat_i[7]
port 564 nsew default input
rlabel metal2 s 15646 0 15702 800 6 wbs_dat_i[8]
port 565 nsew default input
rlabel metal2 s 17026 0 17082 800 6 wbs_dat_i[9]
port 566 nsew default input
rlabel metal2 s 3594 0 3650 800 6 wbs_dat_o[0]
port 567 nsew default output
rlabel metal2 s 18774 0 18830 800 6 wbs_dat_o[10]
port 568 nsew default output
rlabel metal2 s 20154 0 20210 800 6 wbs_dat_o[11]
port 569 nsew default output
rlabel metal2 s 21534 0 21590 800 6 wbs_dat_o[12]
port 570 nsew default output
rlabel metal2 s 22822 0 22878 800 6 wbs_dat_o[13]
port 571 nsew default output
rlabel metal2 s 24202 0 24258 800 6 wbs_dat_o[14]
port 572 nsew default output
rlabel metal2 s 25582 0 25638 800 6 wbs_dat_o[15]
port 573 nsew default output
rlabel metal2 s 26870 0 26926 800 6 wbs_dat_o[16]
port 574 nsew default output
rlabel metal2 s 28250 0 28306 800 6 wbs_dat_o[17]
port 575 nsew default output
rlabel metal2 s 29630 0 29686 800 6 wbs_dat_o[18]
port 576 nsew default output
rlabel metal2 s 30918 0 30974 800 6 wbs_dat_o[19]
port 577 nsew default output
rlabel metal2 s 5342 0 5398 800 6 wbs_dat_o[1]
port 578 nsew default output
rlabel metal2 s 32298 0 32354 800 6 wbs_dat_o[20]
port 579 nsew default output
rlabel metal2 s 33586 0 33642 800 6 wbs_dat_o[21]
port 580 nsew default output
rlabel metal2 s 34966 0 35022 800 6 wbs_dat_o[22]
port 581 nsew default output
rlabel metal2 s 36346 0 36402 800 6 wbs_dat_o[23]
port 582 nsew default output
rlabel metal2 s 37634 0 37690 800 6 wbs_dat_o[24]
port 583 nsew default output
rlabel metal2 s 39014 0 39070 800 6 wbs_dat_o[25]
port 584 nsew default output
rlabel metal2 s 40394 0 40450 800 6 wbs_dat_o[26]
port 585 nsew default output
rlabel metal2 s 41682 0 41738 800 6 wbs_dat_o[27]
port 586 nsew default output
rlabel metal2 s 43062 0 43118 800 6 wbs_dat_o[28]
port 587 nsew default output
rlabel metal2 s 44442 0 44498 800 6 wbs_dat_o[29]
port 588 nsew default output
rlabel metal2 s 7182 0 7238 800 6 wbs_dat_o[2]
port 589 nsew default output
rlabel metal2 s 45730 0 45786 800 6 wbs_dat_o[30]
port 590 nsew default output
rlabel metal2 s 47110 0 47166 800 6 wbs_dat_o[31]
port 591 nsew default output
rlabel metal2 s 8930 0 8986 800 6 wbs_dat_o[3]
port 592 nsew default output
rlabel metal2 s 10770 0 10826 800 6 wbs_dat_o[4]
port 593 nsew default output
rlabel metal2 s 12058 0 12114 800 6 wbs_dat_o[5]
port 594 nsew default output
rlabel metal2 s 13438 0 13494 800 6 wbs_dat_o[6]
port 595 nsew default output
rlabel metal2 s 14818 0 14874 800 6 wbs_dat_o[7]
port 596 nsew default output
rlabel metal2 s 16106 0 16162 800 6 wbs_dat_o[8]
port 597 nsew default output
rlabel metal2 s 17486 0 17542 800 6 wbs_dat_o[9]
port 598 nsew default output
rlabel metal2 s 3962 0 4018 800 6 wbs_sel_i[0]
port 599 nsew default input
rlabel metal2 s 5802 0 5858 800 6 wbs_sel_i[1]
port 600 nsew default input
rlabel metal2 s 7550 0 7606 800 6 wbs_sel_i[2]
port 601 nsew default input
rlabel metal2 s 9390 0 9446 800 6 wbs_sel_i[3]
port 602 nsew default input
rlabel metal2 s 1754 0 1810 800 6 wbs_stb_i
port 603 nsew default input
rlabel metal2 s 2214 0 2270 800 6 wbs_we_i
port 604 nsew default input
rlabel metal4 s 4012 2128 4332 217648 6 VPWR
port 605 nsew power input
rlabel metal4 s 19372 2128 19692 217648 6 VGND
port 606 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 1 0 219578 220000
string LEFview TRUE
<< end >>
