VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2700.000 BY 3700.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 3203.520 2700.000 3204.120 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.280 2.400 369.880 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2686.030 0.000 2686.310 2.400 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 3269.480 2700.000 3270.080 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2691.550 0.000 2691.830 2.400 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 319.330 3697.600 319.610 3700.000 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 3336.120 2700.000 3336.720 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 3402.080 2700.000 3402.680 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.960 2.400 302.560 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 3468.040 2700.000 3468.640 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 248.490 3697.600 248.770 3700.000 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 571.240 2.400 571.840 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 234.640 2.400 235.240 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.320 2.400 167.920 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 2.400 100.600 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 2.400 33.960 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 3534.000 2700.000 3534.600 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 177.190 3697.600 177.470 3700.000 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 106.350 3697.600 106.630 3700.000 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 3599.960 2700.000 3600.560 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 3665.920 2700.000 3666.520 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 35.510 3697.600 35.790 3700.000 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.920 2.400 504.520 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2697.070 0.000 2697.350 2.400 ;
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 674.910 3697.600 675.190 3700.000 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 603.610 3697.600 603.890 3700.000 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 436.600 2.400 437.200 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2680.510 0.000 2680.790 2.400 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 532.770 3697.600 533.050 3700.000 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 461.470 3697.600 461.750 3700.000 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 390.630 3697.600 390.910 3700.000 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 32.680 2700.000 33.280 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 2146.800 2700.000 2147.400 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 2344.680 2700.000 2345.280 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 2543.240 2700.000 2543.840 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 2741.120 2700.000 2741.720 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 3005.640 2700.000 3006.240 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2664.410 3697.600 2664.690 3700.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2380.130 3697.600 2380.410 3700.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2167.150 3697.600 2167.430 3700.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1953.710 3697.600 1953.990 3700.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1740.730 3697.600 1741.010 3700.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 230.560 2700.000 231.160 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1527.290 3697.600 1527.570 3700.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1314.310 3697.600 1314.590 3700.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1101.330 3697.600 1101.610 3700.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 887.890 3697.600 888.170 3700.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3665.920 2.400 3666.520 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3329.320 2.400 3329.920 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3127.360 2.400 3127.960 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2925.400 2.400 2926.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2724.120 2.400 2724.720 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2522.160 2.400 2522.760 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 428.440 2700.000 429.040 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2320.200 2.400 2320.800 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2118.240 2.400 2118.840 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1782.320 2.400 1782.920 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1580.360 2.400 1580.960 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1378.400 2.400 1379.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1176.440 2.400 1177.040 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 974.480 2.400 975.080 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 773.200 2.400 773.800 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 627.000 2700.000 627.600 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 824.880 2700.000 825.480 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 1023.440 2700.000 1024.040 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 1221.320 2700.000 1221.920 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 1551.800 2700.000 1552.400 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 1750.360 2700.000 1750.960 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 1948.240 2700.000 1948.840 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 164.600 2700.000 165.200 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 2278.720 2700.000 2279.320 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 2476.600 2700.000 2477.200 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 2675.160 2700.000 2675.760 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 2873.040 2700.000 2873.640 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 3137.560 2700.000 3138.160 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2522.270 3697.600 2522.550 3700.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2237.990 3697.600 2238.270 3700.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2025.010 3697.600 2025.290 3700.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1811.570 3697.600 1811.850 3700.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1598.590 3697.600 1598.870 3700.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 362.480 2700.000 363.080 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1385.610 3697.600 1385.890 3700.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1172.170 3697.600 1172.450 3700.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 959.190 3697.600 959.470 3700.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 745.750 3697.600 746.030 3700.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 3531.280 2.400 3531.880 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 3194.680 2.400 3195.280 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2992.720 2.400 2993.320 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2791.440 2.400 2792.040 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2589.480 2.400 2590.080 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2387.520 2.400 2388.120 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 561.040 2700.000 561.640 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2185.560 2.400 2186.160 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1983.600 2.400 1984.200 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1647.680 2.400 1648.280 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1445.720 2.400 1446.320 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1243.760 2.400 1244.360 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1041.800 2.400 1042.400 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 840.520 2.400 841.120 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 638.560 2.400 639.160 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 758.920 2700.000 759.520 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 957.480 2700.000 958.080 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 1155.360 2700.000 1155.960 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 1353.920 2700.000 1354.520 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 1684.400 2700.000 1685.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 1882.280 2700.000 1882.880 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 2080.160 2700.000 2080.760 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 98.640 2700.000 99.240 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 2212.760 2700.000 2213.360 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 2410.640 2700.000 2411.240 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 2609.200 2700.000 2609.800 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 2807.080 2700.000 2807.680 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 3071.600 2700.000 3072.200 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2593.570 3697.600 2593.850 3700.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2309.290 3697.600 2309.570 3700.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2095.850 3697.600 2096.130 3700.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1882.870 3697.600 1883.150 3700.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1669.430 3697.600 1669.710 3700.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 296.520 2700.000 297.120 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1456.450 3697.600 1456.730 3700.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1243.470 3697.600 1243.750 3700.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1030.030 3697.600 1030.310 3700.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 817.050 3697.600 817.330 3700.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 3598.600 2.400 3599.200 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 3262.000 2.400 3262.600 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 3060.040 2.400 3060.640 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2858.080 2.400 2858.680 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2656.800 2.400 2657.400 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2454.840 2.400 2455.440 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 495.080 2700.000 495.680 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2252.880 2.400 2253.480 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2050.920 2.400 2051.520 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1715.000 2.400 1715.600 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1513.040 2.400 1513.640 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1311.080 2.400 1311.680 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1109.120 2.400 1109.720 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 907.840 2.400 908.440 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 705.880 2.400 706.480 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 692.960 2700.000 693.560 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 891.520 2700.000 892.120 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 1089.400 2700.000 1090.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 1287.960 2700.000 1288.560 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 1617.760 2700.000 1618.360 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 1816.320 2700.000 1816.920 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 2014.200 2700.000 2014.800 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 580.610 0.000 580.890 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2216.830 0.000 2217.110 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2233.390 0.000 2233.670 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2249.490 0.000 2249.770 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2266.050 0.000 2266.330 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2282.150 0.000 2282.430 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2298.710 0.000 2298.990 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2315.270 0.000 2315.550 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2331.370 0.000 2331.650 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2347.930 0.000 2348.210 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2364.030 0.000 2364.310 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 743.910 0.000 744.190 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2380.590 0.000 2380.870 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2396.690 0.000 2396.970 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2413.250 0.000 2413.530 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2429.810 0.000 2430.090 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2445.910 0.000 2446.190 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2462.470 0.000 2462.750 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2478.570 0.000 2478.850 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2495.130 0.000 2495.410 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2511.230 0.000 2511.510 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2527.790 0.000 2528.070 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 760.470 0.000 760.750 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2544.350 0.000 2544.630 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2560.450 0.000 2560.730 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2577.010 0.000 2577.290 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2593.110 0.000 2593.390 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2609.670 0.000 2609.950 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2625.770 0.000 2626.050 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2642.330 0.000 2642.610 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2658.890 0.000 2659.170 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 776.570 0.000 776.850 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 793.130 0.000 793.410 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 809.690 0.000 809.970 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 825.790 0.000 826.070 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 842.350 0.000 842.630 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 858.450 0.000 858.730 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 875.010 0.000 875.290 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 891.110 0.000 891.390 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 596.710 0.000 596.990 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 907.670 0.000 907.950 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 924.230 0.000 924.510 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 940.330 0.000 940.610 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 956.890 0.000 957.170 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 972.990 0.000 973.270 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 989.550 0.000 989.830 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1005.650 0.000 1005.930 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1022.210 0.000 1022.490 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1038.770 0.000 1039.050 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1054.870 0.000 1055.150 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 613.270 0.000 613.550 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1071.430 0.000 1071.710 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1087.530 0.000 1087.810 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1104.090 0.000 1104.370 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1120.650 0.000 1120.930 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1136.750 0.000 1137.030 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1153.310 0.000 1153.590 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1169.410 0.000 1169.690 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1185.970 0.000 1186.250 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1202.070 0.000 1202.350 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1218.630 0.000 1218.910 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 629.370 0.000 629.650 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1235.190 0.000 1235.470 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1251.290 0.000 1251.570 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1267.850 0.000 1268.130 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1283.950 0.000 1284.230 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1300.510 0.000 1300.790 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1316.610 0.000 1316.890 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1333.170 0.000 1333.450 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1349.730 0.000 1350.010 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1365.830 0.000 1366.110 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1382.390 0.000 1382.670 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 645.930 0.000 646.210 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1398.490 0.000 1398.770 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1415.050 0.000 1415.330 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1431.150 0.000 1431.430 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1447.710 0.000 1447.990 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1464.270 0.000 1464.550 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1480.370 0.000 1480.650 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1496.930 0.000 1497.210 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1513.030 0.000 1513.310 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1529.590 0.000 1529.870 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1545.690 0.000 1545.970 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 662.030 0.000 662.310 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1562.250 0.000 1562.530 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1578.810 0.000 1579.090 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1594.910 0.000 1595.190 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1611.470 0.000 1611.750 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1627.570 0.000 1627.850 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1644.130 0.000 1644.410 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1660.690 0.000 1660.970 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1676.790 0.000 1677.070 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1693.350 0.000 1693.630 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1709.450 0.000 1709.730 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 678.590 0.000 678.870 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1726.010 0.000 1726.290 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1742.110 0.000 1742.390 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1758.670 0.000 1758.950 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1775.230 0.000 1775.510 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1791.330 0.000 1791.610 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1807.890 0.000 1808.170 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1823.990 0.000 1824.270 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1840.550 0.000 1840.830 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1856.650 0.000 1856.930 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1873.210 0.000 1873.490 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 695.150 0.000 695.430 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1889.770 0.000 1890.050 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1905.870 0.000 1906.150 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1922.430 0.000 1922.710 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1938.530 0.000 1938.810 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1955.090 0.000 1955.370 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1971.190 0.000 1971.470 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1987.750 0.000 1988.030 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2004.310 0.000 2004.590 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2020.410 0.000 2020.690 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2036.970 0.000 2037.250 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 711.250 0.000 711.530 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2053.070 0.000 2053.350 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2069.630 0.000 2069.910 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2085.730 0.000 2086.010 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2102.290 0.000 2102.570 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2118.850 0.000 2119.130 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2134.950 0.000 2135.230 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2151.510 0.000 2151.790 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2167.610 0.000 2167.890 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2184.170 0.000 2184.450 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2200.730 0.000 2201.010 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 727.810 0.000 728.090 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 585.670 0.000 585.950 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2222.350 0.000 2222.630 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2238.910 0.000 2239.190 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2255.010 0.000 2255.290 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2271.570 0.000 2271.850 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2287.670 0.000 2287.950 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2304.230 0.000 2304.510 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2320.330 0.000 2320.610 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2336.890 0.000 2337.170 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2353.450 0.000 2353.730 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2369.550 0.000 2369.830 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 749.430 0.000 749.710 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2386.110 0.000 2386.390 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2402.210 0.000 2402.490 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2418.770 0.000 2419.050 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2434.870 0.000 2435.150 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2451.430 0.000 2451.710 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2467.990 0.000 2468.270 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2484.090 0.000 2484.370 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2500.650 0.000 2500.930 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2516.750 0.000 2517.030 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2533.310 0.000 2533.590 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 765.990 0.000 766.270 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2549.410 0.000 2549.690 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2565.970 0.000 2566.250 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2582.530 0.000 2582.810 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2598.630 0.000 2598.910 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2615.190 0.000 2615.470 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2631.290 0.000 2631.570 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2647.850 0.000 2648.130 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2663.950 0.000 2664.230 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 782.090 0.000 782.370 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 798.650 0.000 798.930 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 814.750 0.000 815.030 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 831.310 0.000 831.590 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 847.870 0.000 848.150 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 863.970 0.000 864.250 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 880.530 0.000 880.810 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 896.630 0.000 896.910 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 602.230 0.000 602.510 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 913.190 0.000 913.470 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 929.290 0.000 929.570 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 945.850 0.000 946.130 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 962.410 0.000 962.690 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 978.510 0.000 978.790 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 995.070 0.000 995.350 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1011.170 0.000 1011.450 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1027.730 0.000 1028.010 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1043.830 0.000 1044.110 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1060.390 0.000 1060.670 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 618.790 0.000 619.070 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1076.950 0.000 1077.230 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1093.050 0.000 1093.330 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1109.610 0.000 1109.890 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1125.710 0.000 1125.990 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1142.270 0.000 1142.550 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1158.830 0.000 1159.110 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1174.930 0.000 1175.210 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1191.490 0.000 1191.770 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1207.590 0.000 1207.870 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1224.150 0.000 1224.430 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 634.890 0.000 635.170 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1240.250 0.000 1240.530 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1256.810 0.000 1257.090 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1273.370 0.000 1273.650 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1289.470 0.000 1289.750 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1306.030 0.000 1306.310 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1322.130 0.000 1322.410 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1338.690 0.000 1338.970 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1354.790 0.000 1355.070 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1371.350 0.000 1371.630 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1387.910 0.000 1388.190 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 651.450 0.000 651.730 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1404.010 0.000 1404.290 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1420.570 0.000 1420.850 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1436.670 0.000 1436.950 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1453.230 0.000 1453.510 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1469.330 0.000 1469.610 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1485.890 0.000 1486.170 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1502.450 0.000 1502.730 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1518.550 0.000 1518.830 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1535.110 0.000 1535.390 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1551.210 0.000 1551.490 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 667.550 0.000 667.830 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1567.770 0.000 1568.050 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1583.870 0.000 1584.150 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1600.430 0.000 1600.710 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1616.990 0.000 1617.270 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1633.090 0.000 1633.370 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1649.650 0.000 1649.930 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1665.750 0.000 1666.030 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1682.310 0.000 1682.590 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1698.870 0.000 1699.150 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1714.970 0.000 1715.250 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 684.110 0.000 684.390 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1731.530 0.000 1731.810 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1747.630 0.000 1747.910 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1764.190 0.000 1764.470 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1780.290 0.000 1780.570 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1796.850 0.000 1797.130 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1813.410 0.000 1813.690 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1829.510 0.000 1829.790 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1846.070 0.000 1846.350 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1862.170 0.000 1862.450 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1878.730 0.000 1879.010 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 700.210 0.000 700.490 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1894.830 0.000 1895.110 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1911.390 0.000 1911.670 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1927.950 0.000 1928.230 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1944.050 0.000 1944.330 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1960.610 0.000 1960.890 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1976.710 0.000 1976.990 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1993.270 0.000 1993.550 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2009.370 0.000 2009.650 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2025.930 0.000 2026.210 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2042.490 0.000 2042.770 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 716.770 0.000 717.050 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2058.590 0.000 2058.870 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2075.150 0.000 2075.430 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2091.250 0.000 2091.530 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2107.810 0.000 2108.090 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2123.910 0.000 2124.190 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2140.470 0.000 2140.750 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2157.030 0.000 2157.310 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2173.130 0.000 2173.410 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2189.690 0.000 2189.970 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2205.790 0.000 2206.070 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 733.330 0.000 733.610 2.400 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 591.190 0.000 591.470 2.400 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2227.870 0.000 2228.150 2.400 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2243.970 0.000 2244.250 2.400 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2260.530 0.000 2260.810 2.400 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2277.090 0.000 2277.370 2.400 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2293.190 0.000 2293.470 2.400 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2309.750 0.000 2310.030 2.400 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2325.850 0.000 2326.130 2.400 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2342.410 0.000 2342.690 2.400 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2358.510 0.000 2358.790 2.400 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2375.070 0.000 2375.350 2.400 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 754.950 0.000 755.230 2.400 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2391.630 0.000 2391.910 2.400 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2407.730 0.000 2408.010 2.400 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2424.290 0.000 2424.570 2.400 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2440.390 0.000 2440.670 2.400 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2456.950 0.000 2457.230 2.400 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2473.050 0.000 2473.330 2.400 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2489.610 0.000 2489.890 2.400 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2506.170 0.000 2506.450 2.400 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2522.270 0.000 2522.550 2.400 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2538.830 0.000 2539.110 2.400 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 771.510 0.000 771.790 2.400 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2554.930 0.000 2555.210 2.400 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2571.490 0.000 2571.770 2.400 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2587.590 0.000 2587.870 2.400 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2604.150 0.000 2604.430 2.400 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2620.710 0.000 2620.990 2.400 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2636.810 0.000 2637.090 2.400 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2653.370 0.000 2653.650 2.400 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2669.470 0.000 2669.750 2.400 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 787.610 0.000 787.890 2.400 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 804.170 0.000 804.450 2.400 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 820.270 0.000 820.550 2.400 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 836.830 0.000 837.110 2.400 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 852.930 0.000 853.210 2.400 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 869.490 0.000 869.770 2.400 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 886.050 0.000 886.330 2.400 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 902.150 0.000 902.430 2.400 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 607.750 0.000 608.030 2.400 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 918.710 0.000 918.990 2.400 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 934.810 0.000 935.090 2.400 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 951.370 0.000 951.650 2.400 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 967.470 0.000 967.750 2.400 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 984.030 0.000 984.310 2.400 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1000.590 0.000 1000.870 2.400 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1016.690 0.000 1016.970 2.400 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1033.250 0.000 1033.530 2.400 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1049.350 0.000 1049.630 2.400 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1065.910 0.000 1066.190 2.400 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 623.850 0.000 624.130 2.400 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1082.470 0.000 1082.750 2.400 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1098.570 0.000 1098.850 2.400 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1115.130 0.000 1115.410 2.400 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1131.230 0.000 1131.510 2.400 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1147.790 0.000 1148.070 2.400 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1163.890 0.000 1164.170 2.400 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1180.450 0.000 1180.730 2.400 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1197.010 0.000 1197.290 2.400 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1213.110 0.000 1213.390 2.400 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1229.670 0.000 1229.950 2.400 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 640.410 0.000 640.690 2.400 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1245.770 0.000 1246.050 2.400 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1262.330 0.000 1262.610 2.400 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1278.430 0.000 1278.710 2.400 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1294.990 0.000 1295.270 2.400 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1311.550 0.000 1311.830 2.400 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1327.650 0.000 1327.930 2.400 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1344.210 0.000 1344.490 2.400 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1360.310 0.000 1360.590 2.400 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1376.870 0.000 1377.150 2.400 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1392.970 0.000 1393.250 2.400 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 656.970 0.000 657.250 2.400 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1409.530 0.000 1409.810 2.400 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1426.090 0.000 1426.370 2.400 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1442.190 0.000 1442.470 2.400 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1458.750 0.000 1459.030 2.400 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1474.850 0.000 1475.130 2.400 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1491.410 0.000 1491.690 2.400 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1507.510 0.000 1507.790 2.400 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1524.070 0.000 1524.350 2.400 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1540.630 0.000 1540.910 2.400 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1556.730 0.000 1557.010 2.400 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 673.070 0.000 673.350 2.400 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1573.290 0.000 1573.570 2.400 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1589.390 0.000 1589.670 2.400 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1605.950 0.000 1606.230 2.400 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1622.510 0.000 1622.790 2.400 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1638.610 0.000 1638.890 2.400 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1655.170 0.000 1655.450 2.400 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1671.270 0.000 1671.550 2.400 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1687.830 0.000 1688.110 2.400 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1703.930 0.000 1704.210 2.400 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1720.490 0.000 1720.770 2.400 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 689.630 0.000 689.910 2.400 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1737.050 0.000 1737.330 2.400 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1753.150 0.000 1753.430 2.400 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1769.710 0.000 1769.990 2.400 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1785.810 0.000 1786.090 2.400 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1802.370 0.000 1802.650 2.400 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1818.470 0.000 1818.750 2.400 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1835.030 0.000 1835.310 2.400 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1851.590 0.000 1851.870 2.400 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1867.690 0.000 1867.970 2.400 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1884.250 0.000 1884.530 2.400 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 705.730 0.000 706.010 2.400 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1900.350 0.000 1900.630 2.400 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1916.910 0.000 1917.190 2.400 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1933.010 0.000 1933.290 2.400 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1949.570 0.000 1949.850 2.400 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1966.130 0.000 1966.410 2.400 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1982.230 0.000 1982.510 2.400 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1998.790 0.000 1999.070 2.400 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2014.890 0.000 2015.170 2.400 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2031.450 0.000 2031.730 2.400 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2047.550 0.000 2047.830 2.400 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 722.290 0.000 722.570 2.400 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2064.110 0.000 2064.390 2.400 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2080.670 0.000 2080.950 2.400 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2096.770 0.000 2097.050 2.400 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2113.330 0.000 2113.610 2.400 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2129.430 0.000 2129.710 2.400 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2145.990 0.000 2146.270 2.400 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2162.550 0.000 2162.830 2.400 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2178.650 0.000 2178.930 2.400 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2195.210 0.000 2195.490 2.400 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2211.310 0.000 2211.590 2.400 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 738.390 0.000 738.670 2.400 ;
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2674.990 0.000 2675.270 2.400 ;
    END
  END user_clock2
  PIN vccd1
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 2939.680 2700.000 2940.280 ;
    END
  END vccd1
  PIN vccd2
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3463.960 2.400 3464.560 ;
    END
  END vccd2
  PIN vdda1
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 1485.840 2700.000 1486.440 ;
    END
  END vdda1
  PIN vdda2
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1916.280 2.400 1916.880 ;
    END
  END vdda2
  PIN vssa1
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2451.430 3697.600 2451.710 3700.000 ;
    END
  END vssa1
  PIN vssa2
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3396.640 2.400 3397.240 ;
    END
  END vssa2
  PIN vssd1
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 1419.880 2700.000 1420.480 ;
    END
  END vssd1
  PIN vssd2
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1849.640 2.400 1850.240 ;
    END
  END vssd2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 220.430 0.000 220.710 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 236.530 0.000 236.810 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 253.090 0.000 253.370 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 269.650 0.000 269.930 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 285.750 0.000 286.030 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 302.310 0.000 302.590 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 318.410 0.000 318.690 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 334.970 0.000 335.250 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 351.070 0.000 351.350 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 367.630 0.000 367.910 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.670 0.000 56.950 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 384.190 0.000 384.470 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 400.290 0.000 400.570 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 416.850 0.000 417.130 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 432.950 0.000 433.230 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 449.510 0.000 449.790 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 465.610 0.000 465.890 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 482.170 0.000 482.450 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 498.730 0.000 499.010 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 514.830 0.000 515.110 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 531.390 0.000 531.670 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 78.750 0.000 79.030 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 547.490 0.000 547.770 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 564.050 0.000 564.330 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 100.370 0.000 100.650 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 121.990 0.000 122.270 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 155.110 0.000 155.390 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 171.210 0.000 171.490 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 187.770 0.000 188.050 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 203.870 0.000 204.150 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 225.950 0.000 226.230 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 242.050 0.000 242.330 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 258.610 0.000 258.890 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 274.710 0.000 274.990 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 291.270 0.000 291.550 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 307.830 0.000 308.110 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 323.930 0.000 324.210 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 340.490 0.000 340.770 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 356.590 0.000 356.870 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 373.150 0.000 373.430 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 62.190 0.000 62.470 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 389.250 0.000 389.530 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 405.810 0.000 406.090 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 422.370 0.000 422.650 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 438.470 0.000 438.750 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 455.030 0.000 455.310 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 471.130 0.000 471.410 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 487.690 0.000 487.970 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 503.790 0.000 504.070 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 520.350 0.000 520.630 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 536.910 0.000 537.190 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 553.010 0.000 553.290 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 569.570 0.000 569.850 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 105.890 0.000 106.170 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 127.510 0.000 127.790 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 144.070 0.000 144.350 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 160.170 0.000 160.450 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 176.730 0.000 177.010 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 45.630 0.000 45.910 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 231.470 0.000 231.750 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 247.570 0.000 247.850 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 280.230 0.000 280.510 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 296.790 0.000 297.070 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 312.890 0.000 313.170 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 329.450 0.000 329.730 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 346.010 0.000 346.290 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 362.110 0.000 362.390 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 378.670 0.000 378.950 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 394.770 0.000 395.050 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 411.330 0.000 411.610 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 427.430 0.000 427.710 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 443.990 0.000 444.270 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 460.550 0.000 460.830 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 476.650 0.000 476.930 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 493.210 0.000 493.490 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 509.310 0.000 509.590 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 525.870 0.000 526.150 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 542.430 0.000 542.710 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 89.330 0.000 89.610 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 558.530 0.000 558.810 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 575.090 0.000 575.370 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 111.410 0.000 111.690 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 133.030 0.000 133.310 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 149.590 0.000 149.870 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 165.690 0.000 165.970 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 182.250 0.000 182.530 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 198.350 0.000 198.630 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 214.910 0.000 215.190 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 51.150 0.000 51.430 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 73.230 0.000 73.510 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 94.850 0.000 95.130 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 116.930 0.000 117.210 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.010 0.000 24.290 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 29.530 0.000 29.810 2.400 ;
    END
  END wbs_we_i
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.490 2694.220 28.090 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 103.080 2694.220 104.680 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2694.220 3688.405 ;
      LAYER met1 ;
        RECT 2.370 2.760 2694.220 3688.560 ;
      LAYER met2 ;
        RECT 2.400 3697.320 35.230 3698.250 ;
        RECT 36.070 3697.320 106.070 3698.250 ;
        RECT 106.910 3697.320 176.910 3698.250 ;
        RECT 177.750 3697.320 248.210 3698.250 ;
        RECT 249.050 3697.320 319.050 3698.250 ;
        RECT 319.890 3697.320 390.350 3698.250 ;
        RECT 391.190 3697.320 461.190 3698.250 ;
        RECT 462.030 3697.320 532.490 3698.250 ;
        RECT 533.330 3697.320 603.330 3698.250 ;
        RECT 604.170 3697.320 674.630 3698.250 ;
        RECT 675.470 3697.320 745.470 3698.250 ;
        RECT 746.310 3697.320 816.770 3698.250 ;
        RECT 817.610 3697.320 887.610 3698.250 ;
        RECT 888.450 3697.320 958.910 3698.250 ;
        RECT 959.750 3697.320 1029.750 3698.250 ;
        RECT 1030.590 3697.320 1101.050 3698.250 ;
        RECT 1101.890 3697.320 1171.890 3698.250 ;
        RECT 1172.730 3697.320 1243.190 3698.250 ;
        RECT 1244.030 3697.320 1314.030 3698.250 ;
        RECT 1314.870 3697.320 1385.330 3698.250 ;
        RECT 1386.170 3697.320 1456.170 3698.250 ;
        RECT 1457.010 3697.320 1527.010 3698.250 ;
        RECT 1527.850 3697.320 1598.310 3698.250 ;
        RECT 1599.150 3697.320 1669.150 3698.250 ;
        RECT 1669.990 3697.320 1740.450 3698.250 ;
        RECT 1741.290 3697.320 1811.290 3698.250 ;
        RECT 1812.130 3697.320 1882.590 3698.250 ;
        RECT 1883.430 3697.320 1953.430 3698.250 ;
        RECT 1954.270 3697.320 2024.730 3698.250 ;
        RECT 2025.570 3697.320 2095.570 3698.250 ;
        RECT 2096.410 3697.320 2166.870 3698.250 ;
        RECT 2167.710 3697.320 2237.710 3698.250 ;
        RECT 2238.550 3697.320 2309.010 3698.250 ;
        RECT 2309.850 3697.320 2379.850 3698.250 ;
        RECT 2380.690 3697.320 2451.150 3698.250 ;
        RECT 2451.990 3697.320 2521.990 3698.250 ;
        RECT 2522.830 3697.320 2593.290 3698.250 ;
        RECT 2594.130 3697.320 2664.130 3698.250 ;
        RECT 2664.970 3697.320 2689.070 3698.250 ;
        RECT 2.400 2.680 2689.070 3697.320 ;
        RECT 2.950 2.400 7.170 2.680 ;
        RECT 8.010 2.400 12.690 2.680 ;
        RECT 13.530 2.400 18.210 2.680 ;
        RECT 19.050 2.400 23.730 2.680 ;
        RECT 24.570 2.400 29.250 2.680 ;
        RECT 30.090 2.400 34.770 2.680 ;
        RECT 35.610 2.400 40.290 2.680 ;
        RECT 41.130 2.400 45.350 2.680 ;
        RECT 46.190 2.400 50.870 2.680 ;
        RECT 51.710 2.400 56.390 2.680 ;
        RECT 57.230 2.400 61.910 2.680 ;
        RECT 62.750 2.400 67.430 2.680 ;
        RECT 68.270 2.400 72.950 2.680 ;
        RECT 73.790 2.400 78.470 2.680 ;
        RECT 79.310 2.400 83.530 2.680 ;
        RECT 84.370 2.400 89.050 2.680 ;
        RECT 89.890 2.400 94.570 2.680 ;
        RECT 95.410 2.400 100.090 2.680 ;
        RECT 100.930 2.400 105.610 2.680 ;
        RECT 106.450 2.400 111.130 2.680 ;
        RECT 111.970 2.400 116.650 2.680 ;
        RECT 117.490 2.400 121.710 2.680 ;
        RECT 122.550 2.400 127.230 2.680 ;
        RECT 128.070 2.400 132.750 2.680 ;
        RECT 133.590 2.400 138.270 2.680 ;
        RECT 139.110 2.400 143.790 2.680 ;
        RECT 144.630 2.400 149.310 2.680 ;
        RECT 150.150 2.400 154.830 2.680 ;
        RECT 155.670 2.400 159.890 2.680 ;
        RECT 160.730 2.400 165.410 2.680 ;
        RECT 166.250 2.400 170.930 2.680 ;
        RECT 171.770 2.400 176.450 2.680 ;
        RECT 177.290 2.400 181.970 2.680 ;
        RECT 182.810 2.400 187.490 2.680 ;
        RECT 188.330 2.400 193.010 2.680 ;
        RECT 193.850 2.400 198.070 2.680 ;
        RECT 198.910 2.400 203.590 2.680 ;
        RECT 204.430 2.400 209.110 2.680 ;
        RECT 209.950 2.400 214.630 2.680 ;
        RECT 215.470 2.400 220.150 2.680 ;
        RECT 220.990 2.400 225.670 2.680 ;
        RECT 226.510 2.400 231.190 2.680 ;
        RECT 232.030 2.400 236.250 2.680 ;
        RECT 237.090 2.400 241.770 2.680 ;
        RECT 242.610 2.400 247.290 2.680 ;
        RECT 248.130 2.400 252.810 2.680 ;
        RECT 253.650 2.400 258.330 2.680 ;
        RECT 259.170 2.400 263.850 2.680 ;
        RECT 264.690 2.400 269.370 2.680 ;
        RECT 270.210 2.400 274.430 2.680 ;
        RECT 275.270 2.400 279.950 2.680 ;
        RECT 280.790 2.400 285.470 2.680 ;
        RECT 286.310 2.400 290.990 2.680 ;
        RECT 291.830 2.400 296.510 2.680 ;
        RECT 297.350 2.400 302.030 2.680 ;
        RECT 302.870 2.400 307.550 2.680 ;
        RECT 308.390 2.400 312.610 2.680 ;
        RECT 313.450 2.400 318.130 2.680 ;
        RECT 318.970 2.400 323.650 2.680 ;
        RECT 324.490 2.400 329.170 2.680 ;
        RECT 330.010 2.400 334.690 2.680 ;
        RECT 335.530 2.400 340.210 2.680 ;
        RECT 341.050 2.400 345.730 2.680 ;
        RECT 346.570 2.400 350.790 2.680 ;
        RECT 351.630 2.400 356.310 2.680 ;
        RECT 357.150 2.400 361.830 2.680 ;
        RECT 362.670 2.400 367.350 2.680 ;
        RECT 368.190 2.400 372.870 2.680 ;
        RECT 373.710 2.400 378.390 2.680 ;
        RECT 379.230 2.400 383.910 2.680 ;
        RECT 384.750 2.400 388.970 2.680 ;
        RECT 389.810 2.400 394.490 2.680 ;
        RECT 395.330 2.400 400.010 2.680 ;
        RECT 400.850 2.400 405.530 2.680 ;
        RECT 406.370 2.400 411.050 2.680 ;
        RECT 411.890 2.400 416.570 2.680 ;
        RECT 417.410 2.400 422.090 2.680 ;
        RECT 422.930 2.400 427.150 2.680 ;
        RECT 427.990 2.400 432.670 2.680 ;
        RECT 433.510 2.400 438.190 2.680 ;
        RECT 439.030 2.400 443.710 2.680 ;
        RECT 444.550 2.400 449.230 2.680 ;
        RECT 450.070 2.400 454.750 2.680 ;
        RECT 455.590 2.400 460.270 2.680 ;
        RECT 461.110 2.400 465.330 2.680 ;
        RECT 466.170 2.400 470.850 2.680 ;
        RECT 471.690 2.400 476.370 2.680 ;
        RECT 477.210 2.400 481.890 2.680 ;
        RECT 482.730 2.400 487.410 2.680 ;
        RECT 488.250 2.400 492.930 2.680 ;
        RECT 493.770 2.400 498.450 2.680 ;
        RECT 499.290 2.400 503.510 2.680 ;
        RECT 504.350 2.400 509.030 2.680 ;
        RECT 509.870 2.400 514.550 2.680 ;
        RECT 515.390 2.400 520.070 2.680 ;
        RECT 520.910 2.400 525.590 2.680 ;
        RECT 526.430 2.400 531.110 2.680 ;
        RECT 531.950 2.400 536.630 2.680 ;
        RECT 537.470 2.400 542.150 2.680 ;
        RECT 542.990 2.400 547.210 2.680 ;
        RECT 548.050 2.400 552.730 2.680 ;
        RECT 553.570 2.400 558.250 2.680 ;
        RECT 559.090 2.400 563.770 2.680 ;
        RECT 564.610 2.400 569.290 2.680 ;
        RECT 570.130 2.400 574.810 2.680 ;
        RECT 575.650 2.400 580.330 2.680 ;
        RECT 581.170 2.400 585.390 2.680 ;
        RECT 586.230 2.400 590.910 2.680 ;
        RECT 591.750 2.400 596.430 2.680 ;
        RECT 597.270 2.400 601.950 2.680 ;
        RECT 602.790 2.400 607.470 2.680 ;
        RECT 608.310 2.400 612.990 2.680 ;
        RECT 613.830 2.400 618.510 2.680 ;
        RECT 619.350 2.400 623.570 2.680 ;
        RECT 624.410 2.400 629.090 2.680 ;
        RECT 629.930 2.400 634.610 2.680 ;
        RECT 635.450 2.400 640.130 2.680 ;
        RECT 640.970 2.400 645.650 2.680 ;
        RECT 646.490 2.400 651.170 2.680 ;
        RECT 652.010 2.400 656.690 2.680 ;
        RECT 657.530 2.400 661.750 2.680 ;
        RECT 662.590 2.400 667.270 2.680 ;
        RECT 668.110 2.400 672.790 2.680 ;
        RECT 673.630 2.400 678.310 2.680 ;
        RECT 679.150 2.400 683.830 2.680 ;
        RECT 684.670 2.400 689.350 2.680 ;
        RECT 690.190 2.400 694.870 2.680 ;
        RECT 695.710 2.400 699.930 2.680 ;
        RECT 700.770 2.400 705.450 2.680 ;
        RECT 706.290 2.400 710.970 2.680 ;
        RECT 711.810 2.400 716.490 2.680 ;
        RECT 717.330 2.400 722.010 2.680 ;
        RECT 722.850 2.400 727.530 2.680 ;
        RECT 728.370 2.400 733.050 2.680 ;
        RECT 733.890 2.400 738.110 2.680 ;
        RECT 738.950 2.400 743.630 2.680 ;
        RECT 744.470 2.400 749.150 2.680 ;
        RECT 749.990 2.400 754.670 2.680 ;
        RECT 755.510 2.400 760.190 2.680 ;
        RECT 761.030 2.400 765.710 2.680 ;
        RECT 766.550 2.400 771.230 2.680 ;
        RECT 772.070 2.400 776.290 2.680 ;
        RECT 777.130 2.400 781.810 2.680 ;
        RECT 782.650 2.400 787.330 2.680 ;
        RECT 788.170 2.400 792.850 2.680 ;
        RECT 793.690 2.400 798.370 2.680 ;
        RECT 799.210 2.400 803.890 2.680 ;
        RECT 804.730 2.400 809.410 2.680 ;
        RECT 810.250 2.400 814.470 2.680 ;
        RECT 815.310 2.400 819.990 2.680 ;
        RECT 820.830 2.400 825.510 2.680 ;
        RECT 826.350 2.400 831.030 2.680 ;
        RECT 831.870 2.400 836.550 2.680 ;
        RECT 837.390 2.400 842.070 2.680 ;
        RECT 842.910 2.400 847.590 2.680 ;
        RECT 848.430 2.400 852.650 2.680 ;
        RECT 853.490 2.400 858.170 2.680 ;
        RECT 859.010 2.400 863.690 2.680 ;
        RECT 864.530 2.400 869.210 2.680 ;
        RECT 870.050 2.400 874.730 2.680 ;
        RECT 875.570 2.400 880.250 2.680 ;
        RECT 881.090 2.400 885.770 2.680 ;
        RECT 886.610 2.400 890.830 2.680 ;
        RECT 891.670 2.400 896.350 2.680 ;
        RECT 897.190 2.400 901.870 2.680 ;
        RECT 902.710 2.400 907.390 2.680 ;
        RECT 908.230 2.400 912.910 2.680 ;
        RECT 913.750 2.400 918.430 2.680 ;
        RECT 919.270 2.400 923.950 2.680 ;
        RECT 924.790 2.400 929.010 2.680 ;
        RECT 929.850 2.400 934.530 2.680 ;
        RECT 935.370 2.400 940.050 2.680 ;
        RECT 940.890 2.400 945.570 2.680 ;
        RECT 946.410 2.400 951.090 2.680 ;
        RECT 951.930 2.400 956.610 2.680 ;
        RECT 957.450 2.400 962.130 2.680 ;
        RECT 962.970 2.400 967.190 2.680 ;
        RECT 968.030 2.400 972.710 2.680 ;
        RECT 973.550 2.400 978.230 2.680 ;
        RECT 979.070 2.400 983.750 2.680 ;
        RECT 984.590 2.400 989.270 2.680 ;
        RECT 990.110 2.400 994.790 2.680 ;
        RECT 995.630 2.400 1000.310 2.680 ;
        RECT 1001.150 2.400 1005.370 2.680 ;
        RECT 1006.210 2.400 1010.890 2.680 ;
        RECT 1011.730 2.400 1016.410 2.680 ;
        RECT 1017.250 2.400 1021.930 2.680 ;
        RECT 1022.770 2.400 1027.450 2.680 ;
        RECT 1028.290 2.400 1032.970 2.680 ;
        RECT 1033.810 2.400 1038.490 2.680 ;
        RECT 1039.330 2.400 1043.550 2.680 ;
        RECT 1044.390 2.400 1049.070 2.680 ;
        RECT 1049.910 2.400 1054.590 2.680 ;
        RECT 1055.430 2.400 1060.110 2.680 ;
        RECT 1060.950 2.400 1065.630 2.680 ;
        RECT 1066.470 2.400 1071.150 2.680 ;
        RECT 1071.990 2.400 1076.670 2.680 ;
        RECT 1077.510 2.400 1082.190 2.680 ;
        RECT 1083.030 2.400 1087.250 2.680 ;
        RECT 1088.090 2.400 1092.770 2.680 ;
        RECT 1093.610 2.400 1098.290 2.680 ;
        RECT 1099.130 2.400 1103.810 2.680 ;
        RECT 1104.650 2.400 1109.330 2.680 ;
        RECT 1110.170 2.400 1114.850 2.680 ;
        RECT 1115.690 2.400 1120.370 2.680 ;
        RECT 1121.210 2.400 1125.430 2.680 ;
        RECT 1126.270 2.400 1130.950 2.680 ;
        RECT 1131.790 2.400 1136.470 2.680 ;
        RECT 1137.310 2.400 1141.990 2.680 ;
        RECT 1142.830 2.400 1147.510 2.680 ;
        RECT 1148.350 2.400 1153.030 2.680 ;
        RECT 1153.870 2.400 1158.550 2.680 ;
        RECT 1159.390 2.400 1163.610 2.680 ;
        RECT 1164.450 2.400 1169.130 2.680 ;
        RECT 1169.970 2.400 1174.650 2.680 ;
        RECT 1175.490 2.400 1180.170 2.680 ;
        RECT 1181.010 2.400 1185.690 2.680 ;
        RECT 1186.530 2.400 1191.210 2.680 ;
        RECT 1192.050 2.400 1196.730 2.680 ;
        RECT 1197.570 2.400 1201.790 2.680 ;
        RECT 1202.630 2.400 1207.310 2.680 ;
        RECT 1208.150 2.400 1212.830 2.680 ;
        RECT 1213.670 2.400 1218.350 2.680 ;
        RECT 1219.190 2.400 1223.870 2.680 ;
        RECT 1224.710 2.400 1229.390 2.680 ;
        RECT 1230.230 2.400 1234.910 2.680 ;
        RECT 1235.750 2.400 1239.970 2.680 ;
        RECT 1240.810 2.400 1245.490 2.680 ;
        RECT 1246.330 2.400 1251.010 2.680 ;
        RECT 1251.850 2.400 1256.530 2.680 ;
        RECT 1257.370 2.400 1262.050 2.680 ;
        RECT 1262.890 2.400 1267.570 2.680 ;
        RECT 1268.410 2.400 1273.090 2.680 ;
        RECT 1273.930 2.400 1278.150 2.680 ;
        RECT 1278.990 2.400 1283.670 2.680 ;
        RECT 1284.510 2.400 1289.190 2.680 ;
        RECT 1290.030 2.400 1294.710 2.680 ;
        RECT 1295.550 2.400 1300.230 2.680 ;
        RECT 1301.070 2.400 1305.750 2.680 ;
        RECT 1306.590 2.400 1311.270 2.680 ;
        RECT 1312.110 2.400 1316.330 2.680 ;
        RECT 1317.170 2.400 1321.850 2.680 ;
        RECT 1322.690 2.400 1327.370 2.680 ;
        RECT 1328.210 2.400 1332.890 2.680 ;
        RECT 1333.730 2.400 1338.410 2.680 ;
        RECT 1339.250 2.400 1343.930 2.680 ;
        RECT 1344.770 2.400 1349.450 2.680 ;
        RECT 1350.290 2.400 1354.510 2.680 ;
        RECT 1355.350 2.400 1360.030 2.680 ;
        RECT 1360.870 2.400 1365.550 2.680 ;
        RECT 1366.390 2.400 1371.070 2.680 ;
        RECT 1371.910 2.400 1376.590 2.680 ;
        RECT 1377.430 2.400 1382.110 2.680 ;
        RECT 1382.950 2.400 1387.630 2.680 ;
        RECT 1388.470 2.400 1392.690 2.680 ;
        RECT 1393.530 2.400 1398.210 2.680 ;
        RECT 1399.050 2.400 1403.730 2.680 ;
        RECT 1404.570 2.400 1409.250 2.680 ;
        RECT 1410.090 2.400 1414.770 2.680 ;
        RECT 1415.610 2.400 1420.290 2.680 ;
        RECT 1421.130 2.400 1425.810 2.680 ;
        RECT 1426.650 2.400 1430.870 2.680 ;
        RECT 1431.710 2.400 1436.390 2.680 ;
        RECT 1437.230 2.400 1441.910 2.680 ;
        RECT 1442.750 2.400 1447.430 2.680 ;
        RECT 1448.270 2.400 1452.950 2.680 ;
        RECT 1453.790 2.400 1458.470 2.680 ;
        RECT 1459.310 2.400 1463.990 2.680 ;
        RECT 1464.830 2.400 1469.050 2.680 ;
        RECT 1469.890 2.400 1474.570 2.680 ;
        RECT 1475.410 2.400 1480.090 2.680 ;
        RECT 1480.930 2.400 1485.610 2.680 ;
        RECT 1486.450 2.400 1491.130 2.680 ;
        RECT 1491.970 2.400 1496.650 2.680 ;
        RECT 1497.490 2.400 1502.170 2.680 ;
        RECT 1503.010 2.400 1507.230 2.680 ;
        RECT 1508.070 2.400 1512.750 2.680 ;
        RECT 1513.590 2.400 1518.270 2.680 ;
        RECT 1519.110 2.400 1523.790 2.680 ;
        RECT 1524.630 2.400 1529.310 2.680 ;
        RECT 1530.150 2.400 1534.830 2.680 ;
        RECT 1535.670 2.400 1540.350 2.680 ;
        RECT 1541.190 2.400 1545.410 2.680 ;
        RECT 1546.250 2.400 1550.930 2.680 ;
        RECT 1551.770 2.400 1556.450 2.680 ;
        RECT 1557.290 2.400 1561.970 2.680 ;
        RECT 1562.810 2.400 1567.490 2.680 ;
        RECT 1568.330 2.400 1573.010 2.680 ;
        RECT 1573.850 2.400 1578.530 2.680 ;
        RECT 1579.370 2.400 1583.590 2.680 ;
        RECT 1584.430 2.400 1589.110 2.680 ;
        RECT 1589.950 2.400 1594.630 2.680 ;
        RECT 1595.470 2.400 1600.150 2.680 ;
        RECT 1600.990 2.400 1605.670 2.680 ;
        RECT 1606.510 2.400 1611.190 2.680 ;
        RECT 1612.030 2.400 1616.710 2.680 ;
        RECT 1617.550 2.400 1622.230 2.680 ;
        RECT 1623.070 2.400 1627.290 2.680 ;
        RECT 1628.130 2.400 1632.810 2.680 ;
        RECT 1633.650 2.400 1638.330 2.680 ;
        RECT 1639.170 2.400 1643.850 2.680 ;
        RECT 1644.690 2.400 1649.370 2.680 ;
        RECT 1650.210 2.400 1654.890 2.680 ;
        RECT 1655.730 2.400 1660.410 2.680 ;
        RECT 1661.250 2.400 1665.470 2.680 ;
        RECT 1666.310 2.400 1670.990 2.680 ;
        RECT 1671.830 2.400 1676.510 2.680 ;
        RECT 1677.350 2.400 1682.030 2.680 ;
        RECT 1682.870 2.400 1687.550 2.680 ;
        RECT 1688.390 2.400 1693.070 2.680 ;
        RECT 1693.910 2.400 1698.590 2.680 ;
        RECT 1699.430 2.400 1703.650 2.680 ;
        RECT 1704.490 2.400 1709.170 2.680 ;
        RECT 1710.010 2.400 1714.690 2.680 ;
        RECT 1715.530 2.400 1720.210 2.680 ;
        RECT 1721.050 2.400 1725.730 2.680 ;
        RECT 1726.570 2.400 1731.250 2.680 ;
        RECT 1732.090 2.400 1736.770 2.680 ;
        RECT 1737.610 2.400 1741.830 2.680 ;
        RECT 1742.670 2.400 1747.350 2.680 ;
        RECT 1748.190 2.400 1752.870 2.680 ;
        RECT 1753.710 2.400 1758.390 2.680 ;
        RECT 1759.230 2.400 1763.910 2.680 ;
        RECT 1764.750 2.400 1769.430 2.680 ;
        RECT 1770.270 2.400 1774.950 2.680 ;
        RECT 1775.790 2.400 1780.010 2.680 ;
        RECT 1780.850 2.400 1785.530 2.680 ;
        RECT 1786.370 2.400 1791.050 2.680 ;
        RECT 1791.890 2.400 1796.570 2.680 ;
        RECT 1797.410 2.400 1802.090 2.680 ;
        RECT 1802.930 2.400 1807.610 2.680 ;
        RECT 1808.450 2.400 1813.130 2.680 ;
        RECT 1813.970 2.400 1818.190 2.680 ;
        RECT 1819.030 2.400 1823.710 2.680 ;
        RECT 1824.550 2.400 1829.230 2.680 ;
        RECT 1830.070 2.400 1834.750 2.680 ;
        RECT 1835.590 2.400 1840.270 2.680 ;
        RECT 1841.110 2.400 1845.790 2.680 ;
        RECT 1846.630 2.400 1851.310 2.680 ;
        RECT 1852.150 2.400 1856.370 2.680 ;
        RECT 1857.210 2.400 1861.890 2.680 ;
        RECT 1862.730 2.400 1867.410 2.680 ;
        RECT 1868.250 2.400 1872.930 2.680 ;
        RECT 1873.770 2.400 1878.450 2.680 ;
        RECT 1879.290 2.400 1883.970 2.680 ;
        RECT 1884.810 2.400 1889.490 2.680 ;
        RECT 1890.330 2.400 1894.550 2.680 ;
        RECT 1895.390 2.400 1900.070 2.680 ;
        RECT 1900.910 2.400 1905.590 2.680 ;
        RECT 1906.430 2.400 1911.110 2.680 ;
        RECT 1911.950 2.400 1916.630 2.680 ;
        RECT 1917.470 2.400 1922.150 2.680 ;
        RECT 1922.990 2.400 1927.670 2.680 ;
        RECT 1928.510 2.400 1932.730 2.680 ;
        RECT 1933.570 2.400 1938.250 2.680 ;
        RECT 1939.090 2.400 1943.770 2.680 ;
        RECT 1944.610 2.400 1949.290 2.680 ;
        RECT 1950.130 2.400 1954.810 2.680 ;
        RECT 1955.650 2.400 1960.330 2.680 ;
        RECT 1961.170 2.400 1965.850 2.680 ;
        RECT 1966.690 2.400 1970.910 2.680 ;
        RECT 1971.750 2.400 1976.430 2.680 ;
        RECT 1977.270 2.400 1981.950 2.680 ;
        RECT 1982.790 2.400 1987.470 2.680 ;
        RECT 1988.310 2.400 1992.990 2.680 ;
        RECT 1993.830 2.400 1998.510 2.680 ;
        RECT 1999.350 2.400 2004.030 2.680 ;
        RECT 2004.870 2.400 2009.090 2.680 ;
        RECT 2009.930 2.400 2014.610 2.680 ;
        RECT 2015.450 2.400 2020.130 2.680 ;
        RECT 2020.970 2.400 2025.650 2.680 ;
        RECT 2026.490 2.400 2031.170 2.680 ;
        RECT 2032.010 2.400 2036.690 2.680 ;
        RECT 2037.530 2.400 2042.210 2.680 ;
        RECT 2043.050 2.400 2047.270 2.680 ;
        RECT 2048.110 2.400 2052.790 2.680 ;
        RECT 2053.630 2.400 2058.310 2.680 ;
        RECT 2059.150 2.400 2063.830 2.680 ;
        RECT 2064.670 2.400 2069.350 2.680 ;
        RECT 2070.190 2.400 2074.870 2.680 ;
        RECT 2075.710 2.400 2080.390 2.680 ;
        RECT 2081.230 2.400 2085.450 2.680 ;
        RECT 2086.290 2.400 2090.970 2.680 ;
        RECT 2091.810 2.400 2096.490 2.680 ;
        RECT 2097.330 2.400 2102.010 2.680 ;
        RECT 2102.850 2.400 2107.530 2.680 ;
        RECT 2108.370 2.400 2113.050 2.680 ;
        RECT 2113.890 2.400 2118.570 2.680 ;
        RECT 2119.410 2.400 2123.630 2.680 ;
        RECT 2124.470 2.400 2129.150 2.680 ;
        RECT 2129.990 2.400 2134.670 2.680 ;
        RECT 2135.510 2.400 2140.190 2.680 ;
        RECT 2141.030 2.400 2145.710 2.680 ;
        RECT 2146.550 2.400 2151.230 2.680 ;
        RECT 2152.070 2.400 2156.750 2.680 ;
        RECT 2157.590 2.400 2162.270 2.680 ;
        RECT 2163.110 2.400 2167.330 2.680 ;
        RECT 2168.170 2.400 2172.850 2.680 ;
        RECT 2173.690 2.400 2178.370 2.680 ;
        RECT 2179.210 2.400 2183.890 2.680 ;
        RECT 2184.730 2.400 2189.410 2.680 ;
        RECT 2190.250 2.400 2194.930 2.680 ;
        RECT 2195.770 2.400 2200.450 2.680 ;
        RECT 2201.290 2.400 2205.510 2.680 ;
        RECT 2206.350 2.400 2211.030 2.680 ;
        RECT 2211.870 2.400 2216.550 2.680 ;
        RECT 2217.390 2.400 2222.070 2.680 ;
        RECT 2222.910 2.400 2227.590 2.680 ;
        RECT 2228.430 2.400 2233.110 2.680 ;
        RECT 2233.950 2.400 2238.630 2.680 ;
        RECT 2239.470 2.400 2243.690 2.680 ;
        RECT 2244.530 2.400 2249.210 2.680 ;
        RECT 2250.050 2.400 2254.730 2.680 ;
        RECT 2255.570 2.400 2260.250 2.680 ;
        RECT 2261.090 2.400 2265.770 2.680 ;
        RECT 2266.610 2.400 2271.290 2.680 ;
        RECT 2272.130 2.400 2276.810 2.680 ;
        RECT 2277.650 2.400 2281.870 2.680 ;
        RECT 2282.710 2.400 2287.390 2.680 ;
        RECT 2288.230 2.400 2292.910 2.680 ;
        RECT 2293.750 2.400 2298.430 2.680 ;
        RECT 2299.270 2.400 2303.950 2.680 ;
        RECT 2304.790 2.400 2309.470 2.680 ;
        RECT 2310.310 2.400 2314.990 2.680 ;
        RECT 2315.830 2.400 2320.050 2.680 ;
        RECT 2320.890 2.400 2325.570 2.680 ;
        RECT 2326.410 2.400 2331.090 2.680 ;
        RECT 2331.930 2.400 2336.610 2.680 ;
        RECT 2337.450 2.400 2342.130 2.680 ;
        RECT 2342.970 2.400 2347.650 2.680 ;
        RECT 2348.490 2.400 2353.170 2.680 ;
        RECT 2354.010 2.400 2358.230 2.680 ;
        RECT 2359.070 2.400 2363.750 2.680 ;
        RECT 2364.590 2.400 2369.270 2.680 ;
        RECT 2370.110 2.400 2374.790 2.680 ;
        RECT 2375.630 2.400 2380.310 2.680 ;
        RECT 2381.150 2.400 2385.830 2.680 ;
        RECT 2386.670 2.400 2391.350 2.680 ;
        RECT 2392.190 2.400 2396.410 2.680 ;
        RECT 2397.250 2.400 2401.930 2.680 ;
        RECT 2402.770 2.400 2407.450 2.680 ;
        RECT 2408.290 2.400 2412.970 2.680 ;
        RECT 2413.810 2.400 2418.490 2.680 ;
        RECT 2419.330 2.400 2424.010 2.680 ;
        RECT 2424.850 2.400 2429.530 2.680 ;
        RECT 2430.370 2.400 2434.590 2.680 ;
        RECT 2435.430 2.400 2440.110 2.680 ;
        RECT 2440.950 2.400 2445.630 2.680 ;
        RECT 2446.470 2.400 2451.150 2.680 ;
        RECT 2451.990 2.400 2456.670 2.680 ;
        RECT 2457.510 2.400 2462.190 2.680 ;
        RECT 2463.030 2.400 2467.710 2.680 ;
        RECT 2468.550 2.400 2472.770 2.680 ;
        RECT 2473.610 2.400 2478.290 2.680 ;
        RECT 2479.130 2.400 2483.810 2.680 ;
        RECT 2484.650 2.400 2489.330 2.680 ;
        RECT 2490.170 2.400 2494.850 2.680 ;
        RECT 2495.690 2.400 2500.370 2.680 ;
        RECT 2501.210 2.400 2505.890 2.680 ;
        RECT 2506.730 2.400 2510.950 2.680 ;
        RECT 2511.790 2.400 2516.470 2.680 ;
        RECT 2517.310 2.400 2521.990 2.680 ;
        RECT 2522.830 2.400 2527.510 2.680 ;
        RECT 2528.350 2.400 2533.030 2.680 ;
        RECT 2533.870 2.400 2538.550 2.680 ;
        RECT 2539.390 2.400 2544.070 2.680 ;
        RECT 2544.910 2.400 2549.130 2.680 ;
        RECT 2549.970 2.400 2554.650 2.680 ;
        RECT 2555.490 2.400 2560.170 2.680 ;
        RECT 2561.010 2.400 2565.690 2.680 ;
        RECT 2566.530 2.400 2571.210 2.680 ;
        RECT 2572.050 2.400 2576.730 2.680 ;
        RECT 2577.570 2.400 2582.250 2.680 ;
        RECT 2583.090 2.400 2587.310 2.680 ;
        RECT 2588.150 2.400 2592.830 2.680 ;
        RECT 2593.670 2.400 2598.350 2.680 ;
        RECT 2599.190 2.400 2603.870 2.680 ;
        RECT 2604.710 2.400 2609.390 2.680 ;
        RECT 2610.230 2.400 2614.910 2.680 ;
        RECT 2615.750 2.400 2620.430 2.680 ;
        RECT 2621.270 2.400 2625.490 2.680 ;
        RECT 2626.330 2.400 2631.010 2.680 ;
        RECT 2631.850 2.400 2636.530 2.680 ;
        RECT 2637.370 2.400 2642.050 2.680 ;
        RECT 2642.890 2.400 2647.570 2.680 ;
        RECT 2648.410 2.400 2653.090 2.680 ;
        RECT 2653.930 2.400 2658.610 2.680 ;
        RECT 2659.450 2.400 2663.670 2.680 ;
        RECT 2664.510 2.400 2669.190 2.680 ;
        RECT 2670.030 2.400 2674.710 2.680 ;
        RECT 2675.550 2.400 2680.230 2.680 ;
        RECT 2681.070 2.400 2685.750 2.680 ;
        RECT 2686.590 2.400 2689.070 2.680 ;
      LAYER met3 ;
        RECT 2.400 3666.920 2697.600 3697.665 ;
        RECT 2.800 3665.520 2697.200 3666.920 ;
        RECT 2.400 3600.960 2697.600 3665.520 ;
        RECT 2.400 3599.600 2697.200 3600.960 ;
        RECT 2.800 3599.560 2697.200 3599.600 ;
        RECT 2.800 3598.200 2697.600 3599.560 ;
        RECT 2.400 3535.000 2697.600 3598.200 ;
        RECT 2.400 3533.600 2697.200 3535.000 ;
        RECT 2.400 3532.280 2697.600 3533.600 ;
        RECT 2.800 3530.880 2697.600 3532.280 ;
        RECT 2.400 3469.040 2697.600 3530.880 ;
        RECT 2.400 3467.640 2697.200 3469.040 ;
        RECT 2.400 3464.960 2697.600 3467.640 ;
        RECT 2.800 3463.560 2697.600 3464.960 ;
        RECT 2.400 3403.080 2697.600 3463.560 ;
        RECT 2.400 3401.680 2697.200 3403.080 ;
        RECT 2.400 3397.640 2697.600 3401.680 ;
        RECT 2.800 3396.240 2697.600 3397.640 ;
        RECT 2.400 3337.120 2697.600 3396.240 ;
        RECT 2.400 3335.720 2697.200 3337.120 ;
        RECT 2.400 3330.320 2697.600 3335.720 ;
        RECT 2.800 3328.920 2697.600 3330.320 ;
        RECT 2.400 3270.480 2697.600 3328.920 ;
        RECT 2.400 3269.080 2697.200 3270.480 ;
        RECT 2.400 3263.000 2697.600 3269.080 ;
        RECT 2.800 3261.600 2697.600 3263.000 ;
        RECT 2.400 3204.520 2697.600 3261.600 ;
        RECT 2.400 3203.120 2697.200 3204.520 ;
        RECT 2.400 3195.680 2697.600 3203.120 ;
        RECT 2.800 3194.280 2697.600 3195.680 ;
        RECT 2.400 3138.560 2697.600 3194.280 ;
        RECT 2.400 3137.160 2697.200 3138.560 ;
        RECT 2.400 3128.360 2697.600 3137.160 ;
        RECT 2.800 3126.960 2697.600 3128.360 ;
        RECT 2.400 3072.600 2697.600 3126.960 ;
        RECT 2.400 3071.200 2697.200 3072.600 ;
        RECT 2.400 3061.040 2697.600 3071.200 ;
        RECT 2.800 3059.640 2697.600 3061.040 ;
        RECT 2.400 3006.640 2697.600 3059.640 ;
        RECT 2.400 3005.240 2697.200 3006.640 ;
        RECT 2.400 2993.720 2697.600 3005.240 ;
        RECT 2.800 2992.320 2697.600 2993.720 ;
        RECT 2.400 2940.680 2697.600 2992.320 ;
        RECT 2.400 2939.280 2697.200 2940.680 ;
        RECT 2.400 2926.400 2697.600 2939.280 ;
        RECT 2.800 2925.000 2697.600 2926.400 ;
        RECT 2.400 2874.040 2697.600 2925.000 ;
        RECT 2.400 2872.640 2697.200 2874.040 ;
        RECT 2.400 2859.080 2697.600 2872.640 ;
        RECT 2.800 2857.680 2697.600 2859.080 ;
        RECT 2.400 2808.080 2697.600 2857.680 ;
        RECT 2.400 2806.680 2697.200 2808.080 ;
        RECT 2.400 2792.440 2697.600 2806.680 ;
        RECT 2.800 2791.040 2697.600 2792.440 ;
        RECT 2.400 2742.120 2697.600 2791.040 ;
        RECT 2.400 2740.720 2697.200 2742.120 ;
        RECT 2.400 2725.120 2697.600 2740.720 ;
        RECT 2.800 2723.720 2697.600 2725.120 ;
        RECT 2.400 2676.160 2697.600 2723.720 ;
        RECT 2.400 2674.760 2697.200 2676.160 ;
        RECT 2.400 2657.800 2697.600 2674.760 ;
        RECT 2.800 2656.400 2697.600 2657.800 ;
        RECT 2.400 2610.200 2697.600 2656.400 ;
        RECT 2.400 2608.800 2697.200 2610.200 ;
        RECT 2.400 2590.480 2697.600 2608.800 ;
        RECT 2.800 2589.080 2697.600 2590.480 ;
        RECT 2.400 2544.240 2697.600 2589.080 ;
        RECT 2.400 2542.840 2697.200 2544.240 ;
        RECT 2.400 2523.160 2697.600 2542.840 ;
        RECT 2.800 2521.760 2697.600 2523.160 ;
        RECT 2.400 2477.600 2697.600 2521.760 ;
        RECT 2.400 2476.200 2697.200 2477.600 ;
        RECT 2.400 2455.840 2697.600 2476.200 ;
        RECT 2.800 2454.440 2697.600 2455.840 ;
        RECT 2.400 2411.640 2697.600 2454.440 ;
        RECT 2.400 2410.240 2697.200 2411.640 ;
        RECT 2.400 2388.520 2697.600 2410.240 ;
        RECT 2.800 2387.120 2697.600 2388.520 ;
        RECT 2.400 2345.680 2697.600 2387.120 ;
        RECT 2.400 2344.280 2697.200 2345.680 ;
        RECT 2.400 2321.200 2697.600 2344.280 ;
        RECT 2.800 2319.800 2697.600 2321.200 ;
        RECT 2.400 2279.720 2697.600 2319.800 ;
        RECT 2.400 2278.320 2697.200 2279.720 ;
        RECT 2.400 2253.880 2697.600 2278.320 ;
        RECT 2.800 2252.480 2697.600 2253.880 ;
        RECT 2.400 2213.760 2697.600 2252.480 ;
        RECT 2.400 2212.360 2697.200 2213.760 ;
        RECT 2.400 2186.560 2697.600 2212.360 ;
        RECT 2.800 2185.160 2697.600 2186.560 ;
        RECT 2.400 2147.800 2697.600 2185.160 ;
        RECT 2.400 2146.400 2697.200 2147.800 ;
        RECT 2.400 2119.240 2697.600 2146.400 ;
        RECT 2.800 2117.840 2697.600 2119.240 ;
        RECT 2.400 2081.160 2697.600 2117.840 ;
        RECT 2.400 2079.760 2697.200 2081.160 ;
        RECT 2.400 2051.920 2697.600 2079.760 ;
        RECT 2.800 2050.520 2697.600 2051.920 ;
        RECT 2.400 2015.200 2697.600 2050.520 ;
        RECT 2.400 2013.800 2697.200 2015.200 ;
        RECT 2.400 1984.600 2697.600 2013.800 ;
        RECT 2.800 1983.200 2697.600 1984.600 ;
        RECT 2.400 1949.240 2697.600 1983.200 ;
        RECT 2.400 1947.840 2697.200 1949.240 ;
        RECT 2.400 1917.280 2697.600 1947.840 ;
        RECT 2.800 1915.880 2697.600 1917.280 ;
        RECT 2.400 1883.280 2697.600 1915.880 ;
        RECT 2.400 1881.880 2697.200 1883.280 ;
        RECT 2.400 1850.640 2697.600 1881.880 ;
        RECT 2.800 1849.240 2697.600 1850.640 ;
        RECT 2.400 1817.320 2697.600 1849.240 ;
        RECT 2.400 1815.920 2697.200 1817.320 ;
        RECT 2.400 1783.320 2697.600 1815.920 ;
        RECT 2.800 1781.920 2697.600 1783.320 ;
        RECT 2.400 1751.360 2697.600 1781.920 ;
        RECT 2.400 1749.960 2697.200 1751.360 ;
        RECT 2.400 1716.000 2697.600 1749.960 ;
        RECT 2.800 1714.600 2697.600 1716.000 ;
        RECT 2.400 1685.400 2697.600 1714.600 ;
        RECT 2.400 1684.000 2697.200 1685.400 ;
        RECT 2.400 1648.680 2697.600 1684.000 ;
        RECT 2.800 1647.280 2697.600 1648.680 ;
        RECT 2.400 1618.760 2697.600 1647.280 ;
        RECT 2.400 1617.360 2697.200 1618.760 ;
        RECT 2.400 1581.360 2697.600 1617.360 ;
        RECT 2.800 1579.960 2697.600 1581.360 ;
        RECT 2.400 1552.800 2697.600 1579.960 ;
        RECT 2.400 1551.400 2697.200 1552.800 ;
        RECT 2.400 1514.040 2697.600 1551.400 ;
        RECT 2.800 1512.640 2697.600 1514.040 ;
        RECT 2.400 1486.840 2697.600 1512.640 ;
        RECT 2.400 1485.440 2697.200 1486.840 ;
        RECT 2.400 1446.720 2697.600 1485.440 ;
        RECT 2.800 1445.320 2697.600 1446.720 ;
        RECT 2.400 1420.880 2697.600 1445.320 ;
        RECT 2.400 1419.480 2697.200 1420.880 ;
        RECT 2.400 1379.400 2697.600 1419.480 ;
        RECT 2.800 1378.000 2697.600 1379.400 ;
        RECT 2.400 1354.920 2697.600 1378.000 ;
        RECT 2.400 1353.520 2697.200 1354.920 ;
        RECT 2.400 1312.080 2697.600 1353.520 ;
        RECT 2.800 1310.680 2697.600 1312.080 ;
        RECT 2.400 1288.960 2697.600 1310.680 ;
        RECT 2.400 1287.560 2697.200 1288.960 ;
        RECT 2.400 1244.760 2697.600 1287.560 ;
        RECT 2.800 1243.360 2697.600 1244.760 ;
        RECT 2.400 1222.320 2697.600 1243.360 ;
        RECT 2.400 1220.920 2697.200 1222.320 ;
        RECT 2.400 1177.440 2697.600 1220.920 ;
        RECT 2.800 1176.040 2697.600 1177.440 ;
        RECT 2.400 1156.360 2697.600 1176.040 ;
        RECT 2.400 1154.960 2697.200 1156.360 ;
        RECT 2.400 1110.120 2697.600 1154.960 ;
        RECT 2.800 1108.720 2697.600 1110.120 ;
        RECT 2.400 1090.400 2697.600 1108.720 ;
        RECT 2.400 1089.000 2697.200 1090.400 ;
        RECT 2.400 1042.800 2697.600 1089.000 ;
        RECT 2.800 1041.400 2697.600 1042.800 ;
        RECT 2.400 1024.440 2697.600 1041.400 ;
        RECT 2.400 1023.040 2697.200 1024.440 ;
        RECT 2.400 975.480 2697.600 1023.040 ;
        RECT 2.800 974.080 2697.600 975.480 ;
        RECT 2.400 958.480 2697.600 974.080 ;
        RECT 2.400 957.080 2697.200 958.480 ;
        RECT 2.400 908.840 2697.600 957.080 ;
        RECT 2.800 907.440 2697.600 908.840 ;
        RECT 2.400 892.520 2697.600 907.440 ;
        RECT 2.400 891.120 2697.200 892.520 ;
        RECT 2.400 841.520 2697.600 891.120 ;
        RECT 2.800 840.120 2697.600 841.520 ;
        RECT 2.400 825.880 2697.600 840.120 ;
        RECT 2.400 824.480 2697.200 825.880 ;
        RECT 2.400 774.200 2697.600 824.480 ;
        RECT 2.800 772.800 2697.600 774.200 ;
        RECT 2.400 759.920 2697.600 772.800 ;
        RECT 2.400 758.520 2697.200 759.920 ;
        RECT 2.400 706.880 2697.600 758.520 ;
        RECT 2.800 705.480 2697.600 706.880 ;
        RECT 2.400 693.960 2697.600 705.480 ;
        RECT 2.400 692.560 2697.200 693.960 ;
        RECT 2.400 639.560 2697.600 692.560 ;
        RECT 2.800 638.160 2697.600 639.560 ;
        RECT 2.400 628.000 2697.600 638.160 ;
        RECT 2.400 626.600 2697.200 628.000 ;
        RECT 2.400 572.240 2697.600 626.600 ;
        RECT 2.800 570.840 2697.600 572.240 ;
        RECT 2.400 562.040 2697.600 570.840 ;
        RECT 2.400 560.640 2697.200 562.040 ;
        RECT 2.400 504.920 2697.600 560.640 ;
        RECT 2.800 503.520 2697.600 504.920 ;
        RECT 2.400 496.080 2697.600 503.520 ;
        RECT 2.400 494.680 2697.200 496.080 ;
        RECT 2.400 437.600 2697.600 494.680 ;
        RECT 2.800 436.200 2697.600 437.600 ;
        RECT 2.400 429.440 2697.600 436.200 ;
        RECT 2.400 428.040 2697.200 429.440 ;
        RECT 2.400 370.280 2697.600 428.040 ;
        RECT 2.800 368.880 2697.600 370.280 ;
        RECT 2.400 363.480 2697.600 368.880 ;
        RECT 2.400 362.080 2697.200 363.480 ;
        RECT 2.400 302.960 2697.600 362.080 ;
        RECT 2.800 301.560 2697.600 302.960 ;
        RECT 2.400 297.520 2697.600 301.560 ;
        RECT 2.400 296.120 2697.200 297.520 ;
        RECT 2.400 235.640 2697.600 296.120 ;
        RECT 2.800 234.240 2697.600 235.640 ;
        RECT 2.400 231.560 2697.600 234.240 ;
        RECT 2.400 230.160 2697.200 231.560 ;
        RECT 2.400 168.320 2697.600 230.160 ;
        RECT 2.800 166.920 2697.600 168.320 ;
        RECT 2.400 165.600 2697.600 166.920 ;
        RECT 2.400 164.200 2697.200 165.600 ;
        RECT 2.400 101.000 2697.600 164.200 ;
        RECT 2.800 99.640 2697.600 101.000 ;
        RECT 2.800 99.600 2697.200 99.640 ;
        RECT 2.400 98.240 2697.200 99.600 ;
        RECT 2.400 34.360 2697.600 98.240 ;
        RECT 2.800 33.680 2697.600 34.360 ;
        RECT 2.800 32.960 2697.200 33.680 ;
        RECT 2.400 32.280 2697.200 32.960 ;
        RECT 2.400 10.715 2697.600 32.280 ;
      LAYER met4 ;
        RECT 17.775 10.640 2633.840 3688.560 ;
      LAYER met5 ;
        RECT 5.520 179.670 2694.220 3627.820 ;
  END
END user_project_wrapper
END LIBRARY

