magic
tech sky130A
magscale 1 2
timestamp 1607892876
<< locali >>
rect 429577 666587 429611 684437
rect 494069 666587 494103 676141
rect 559297 666587 559331 684437
rect 429393 601715 429427 608549
rect 559113 601715 559147 608549
rect 429577 589339 429611 598893
rect 559297 589339 559331 598893
rect 429485 569959 429519 579581
rect 494069 569959 494103 579581
rect 559297 569959 559331 579581
rect 303997 562955 304031 563057
rect 306941 562955 306975 562989
rect 306941 562921 307125 562955
rect 310471 562921 311817 562955
rect 395353 561051 395387 562105
rect 400263 560881 400413 560915
rect 400355 560813 400505 560847
rect 400355 560677 400505 560711
rect 400263 560609 400413 560643
rect 287805 560235 287839 560609
rect 372203 560541 372353 560575
rect 400355 560541 400505 560575
rect 372295 560473 372445 560507
rect 400263 560473 400413 560507
rect 372387 560405 372537 560439
rect 400355 560405 400505 560439
rect 372387 560269 372537 560303
rect 400355 560269 400505 560303
rect 372203 560201 372261 560235
rect 400355 560133 400505 560167
rect 400355 559997 400505 560031
rect 372203 559929 372721 559963
rect 390603 559861 390753 559895
rect 419583 559861 419641 559895
rect 372203 559793 372537 559827
rect 390695 559793 390845 559827
rect 400263 559793 400413 559827
rect 372295 559725 372445 559759
rect 390695 559657 390845 559691
rect 390603 559589 390753 559623
rect 372295 559521 372353 559555
rect 229753 559283 229787 559453
rect 234629 559419 234663 559521
rect 236745 559351 236779 559453
rect 236653 559283 236687 559317
rect 236837 559283 236871 559385
rect 385325 559351 385359 559385
rect 396273 559385 396457 559419
rect 408359 559385 408509 559419
rect 396273 559351 396307 559385
rect 415869 559351 415903 559385
rect 301731 559317 301881 559351
rect 321051 559317 321201 559351
rect 340371 559317 340521 559351
rect 369811 559317 370053 559351
rect 385325 559317 385509 559351
rect 408451 559317 408601 559351
rect 415869 559317 416053 559351
rect 236653 559249 236871 559283
rect 9689 559011 9723 559113
rect 19257 559011 19291 559181
rect 20453 559079 20487 559181
rect 41521 559147 41555 559181
rect 41371 559113 41555 559147
rect 29009 558943 29043 559045
rect 38577 558943 38611 559113
rect 48329 559011 48363 559181
rect 60841 559147 60875 559181
rect 60691 559113 60875 559147
rect 57897 559011 57931 559113
rect 67649 559011 67683 559181
rect 80161 559147 80195 559181
rect 80011 559113 80195 559147
rect 77217 559011 77251 559113
rect 86969 559011 87003 559181
rect 99481 559147 99515 559181
rect 99331 559113 99515 559147
rect 96537 559011 96571 559113
rect 106289 559011 106323 559181
rect 118801 559147 118835 559181
rect 118651 559113 118835 559147
rect 115857 559011 115891 559113
rect 125609 559011 125643 559181
rect 138121 559147 138155 559181
rect 137971 559113 138155 559147
rect 135177 559011 135211 559113
rect 144929 559011 144963 559181
rect 157441 559147 157475 559181
rect 157291 559113 157475 559147
rect 154497 559011 154531 559113
rect 164249 559011 164283 559181
rect 176761 559147 176795 559181
rect 176611 559113 176795 559147
rect 173817 559011 173851 559113
rect 183569 559011 183603 559181
rect 196081 559147 196115 559181
rect 195931 559113 196115 559147
rect 193137 559011 193171 559113
rect 202889 559011 202923 559181
rect 212457 559011 212491 559113
rect 229845 337535 229879 337705
rect 229937 337467 229971 337705
rect 229695 337433 229971 337467
rect 253857 337467 253891 337773
rect 259377 337739 259411 337841
rect 259469 337807 259503 337977
rect 259595 337569 259745 337603
rect 287713 337331 287747 337637
rect 89637 337127 89671 337297
rect 99389 336923 99423 337297
rect 108957 336923 108991 337297
rect 118709 336787 118743 337297
rect 128277 336719 128311 337297
rect 233525 328491 233559 334441
rect 235089 327131 235123 331925
rect 234813 317475 234847 327029
rect 239137 318835 239171 336685
rect 267013 328491 267047 337229
rect 287437 327131 287471 334305
rect 294061 329443 294095 337977
rect 297373 337331 297407 337909
rect 302157 337875 302191 338045
rect 299397 337059 299431 337229
rect 299489 337059 299523 337229
rect 303445 337195 303479 338045
rect 326261 337399 326295 337637
rect 326169 337331 326203 337365
rect 326445 337331 326479 337569
rect 326169 337297 326479 337331
rect 326203 337161 326353 337195
rect 336565 337059 336599 337977
rect 337945 337331 337979 337773
rect 340061 337399 340095 337705
rect 340245 337331 340279 337569
rect 326445 336787 326479 337025
rect 336657 336923 336691 337025
rect 341717 336991 341751 337841
rect 341809 336923 341843 337297
rect 345489 336787 345523 337365
rect 345581 337059 345615 337501
rect 345673 337399 345707 337705
rect 319177 328491 319211 334169
rect 324697 328355 324731 336685
rect 327457 328491 327491 331177
rect 343833 328491 343867 335529
rect 347973 328491 348007 338045
rect 352849 337875 352883 337977
rect 353033 337535 353067 338045
rect 353493 337535 353527 337705
rect 355149 337535 355183 337909
rect 356621 337467 356655 337705
rect 381829 337535 381863 337977
rect 383577 337807 383611 337977
rect 383853 337195 383887 337705
rect 385969 337263 386003 337841
rect 388545 337195 388579 337841
rect 390569 337739 390603 338045
rect 393237 337331 393271 337501
rect 396917 337467 396951 337977
rect 425621 337739 425655 338113
rect 417065 337467 417099 337637
rect 394559 337365 394801 337399
rect 427001 337331 427035 338045
rect 432429 337943 432463 338045
rect 427093 337263 427127 337909
rect 432521 337875 432555 338045
rect 362877 336991 362911 337161
rect 407773 336787 407807 337093
rect 417433 336991 417467 337229
rect 428105 336719 428139 337433
rect 428289 337399 428323 337501
rect 432705 337467 432739 337841
rect 433349 337671 433383 337773
rect 433441 337671 433475 338181
rect 435281 336515 435315 337569
rect 437029 337467 437063 337705
rect 437305 336651 437339 337841
rect 442181 337535 442215 337841
rect 442273 337467 442307 337841
rect 442917 337535 442951 337705
rect 444941 337535 444975 337637
rect 444791 337501 444975 337535
rect 445677 337399 445711 337637
rect 446965 336787 446999 337705
rect 450001 336787 450035 337569
rect 437615 336753 437765 336787
rect 446965 336753 447057 336787
rect 347973 318835 348007 328321
rect 363245 318835 363279 328389
rect 229293 298163 229327 299557
rect 234905 298163 234939 307717
rect 235089 299523 235123 309077
rect 248797 299523 248831 311933
rect 250085 299523 250119 315945
rect 262689 312171 262723 318733
rect 287345 311831 287379 317373
rect 267013 299523 267047 309009
rect 290105 307819 290139 315877
rect 292865 309179 292899 318733
rect 298477 307819 298511 317373
rect 327457 309179 327491 318733
rect 342545 309179 342579 318733
rect 345213 309179 345247 318733
rect 235089 280211 235123 298061
rect 240425 288439 240459 298061
rect 241897 288439 241931 298061
rect 262597 289935 262631 299421
rect 287345 289867 287379 299421
rect 229385 273139 229419 280109
rect 229385 263483 229419 270453
rect 235089 260899 235123 278681
rect 239321 267767 239355 274057
rect 244289 260899 244323 270453
rect 245945 260899 245979 270453
rect 251465 260899 251499 273853
rect 254225 270555 254259 280109
rect 262505 278851 262539 288337
rect 288725 282863 288759 289697
rect 291485 288439 291519 298061
rect 298477 289867 298511 299421
rect 305469 298163 305503 307717
rect 316325 298163 316359 307717
rect 310805 296735 310839 298129
rect 324605 289935 324639 299421
rect 342453 298163 342487 307717
rect 347973 299591 348007 309009
rect 434269 299523 434303 309077
rect 325985 289867 326019 294661
rect 316233 287079 316267 288473
rect 327273 288439 327307 298061
rect 345213 280279 345247 289765
rect 434269 280211 434303 289765
rect 255605 260899 255639 270385
rect 262505 263483 262539 278681
rect 287345 270555 287379 280109
rect 290105 273003 290139 280109
rect 298477 270623 298511 280109
rect 288725 263551 288759 270385
rect 229385 253827 229419 260797
rect 235089 241519 235123 259369
rect 239137 240159 239171 249849
rect 244289 241519 244323 251141
rect 245945 241519 245979 251141
rect 251465 251107 251499 259369
rect 254225 251243 254259 260797
rect 255605 251243 255639 260729
rect 262597 251243 262631 260797
rect 287345 251243 287379 260797
rect 290105 252875 290139 260797
rect 291485 251311 291519 260797
rect 298477 251311 298511 260797
rect 307953 258111 307987 270453
rect 309425 267767 309459 273173
rect 310713 267835 310747 273377
rect 324513 263483 324547 278681
rect 342545 270555 342579 280109
rect 363153 270555 363187 280109
rect 345213 260967 345247 270453
rect 347973 260967 348007 270453
rect 434269 260899 434303 270453
rect 291485 241519 291519 251141
rect 298477 241519 298511 251141
rect 305193 241519 305227 251141
rect 307953 244239 307987 251141
rect 251465 240159 251499 241485
rect 234905 230503 234939 240057
rect 251465 230503 251499 239989
rect 288725 231863 288759 240057
rect 310805 240023 310839 256649
rect 324605 251243 324639 260797
rect 342545 251243 342579 260797
rect 363153 251243 363187 260797
rect 435281 251311 435315 260797
rect 327273 242675 327307 251141
rect 345213 241519 345247 251141
rect 347973 241519 348007 251141
rect 434269 241519 434303 251141
rect 435097 241519 435131 251141
rect 435097 222207 435131 224961
rect 229293 215271 229327 220745
rect 235089 211191 235123 220745
rect 267013 212551 267047 215305
rect 288725 212551 288759 215305
rect 239137 202827 239171 211089
rect 267013 202827 267047 211089
rect 288817 202895 288851 205649
rect 291393 202963 291427 220745
rect 308045 212551 308079 217413
rect 310897 214591 310931 219385
rect 434269 215271 434303 220745
rect 305285 202895 305319 205649
rect 343741 202827 343775 211089
rect 234813 192287 234847 201433
rect 238861 198067 238895 198441
rect 240425 193171 240459 201433
rect 255605 186303 255639 191777
rect 262597 183515 262631 191777
rect 267013 190519 267047 200073
rect 288725 193239 288759 195993
rect 298477 193239 298511 196061
rect 305285 195959 305319 201433
rect 308045 193239 308079 195993
rect 288817 183583 288851 186337
rect 310805 185623 310839 200073
rect 345029 192763 345063 201433
rect 434453 193239 434487 195993
rect 316233 190519 316267 191845
rect 239137 173859 239171 182121
rect 241805 173927 241839 178789
rect 255605 172567 255639 182121
rect 234905 140879 234939 161313
rect 234997 151827 235031 161381
rect 238861 159375 238895 159681
rect 239045 151827 239079 154649
rect 240425 153323 240459 154581
rect 241897 153255 241931 162809
rect 251373 161483 251407 171037
rect 310805 169779 310839 179333
rect 327365 171139 327399 180761
rect 261309 153255 261343 162809
rect 262505 153255 262539 162809
rect 287345 154615 287379 164169
rect 288725 153867 288759 161381
rect 305285 153255 305319 162809
rect 313565 161483 313599 171037
rect 240333 143599 240367 153153
rect 234813 134623 234847 140709
rect 239137 132515 239171 142069
rect 240333 132515 240367 142069
rect 251557 135235 251591 143497
rect 233433 131155 233467 132481
rect 233433 121499 233467 125477
rect 235089 122859 235123 128333
rect 241897 125647 241931 135201
rect 251465 124219 251499 133841
rect 262689 129795 262723 139349
rect 287253 137819 287287 143497
rect 288817 139519 288851 149005
rect 305285 142171 305319 153085
rect 308045 151827 308079 161381
rect 324605 154615 324639 164169
rect 313657 150467 313691 150569
rect 309517 139451 309551 149005
rect 327365 147611 327399 153493
rect 343925 153255 343959 162809
rect 267105 128299 267139 135201
rect 229293 106335 229327 115889
rect 234905 100759 234939 120037
rect 240333 104907 240367 122757
rect 241897 114563 241931 124117
rect 254225 115991 254259 125545
rect 261217 118643 261251 124117
rect 291577 121499 291611 124185
rect 305377 122859 305411 132413
rect 310805 124219 310839 133841
rect 316325 132515 316359 142069
rect 343833 135303 343867 148325
rect 345213 144959 345247 162809
rect 434453 154615 434487 159137
rect 444113 157335 444147 164169
rect 444113 145027 444147 154513
rect 434453 137955 434487 143497
rect 327365 128299 327399 135201
rect 444113 128299 444147 143497
rect 245945 106335 245979 115889
rect 255605 104907 255639 114461
rect 229293 87023 229327 96577
rect 234813 92055 234847 100725
rect 241805 95251 241839 104805
rect 251465 95319 251499 104805
rect 262689 102187 262723 120037
rect 328469 118643 328503 125545
rect 287345 104907 287379 114461
rect 288725 104907 288759 114461
rect 298477 108851 298511 115889
rect 240517 84235 240551 93789
rect 244473 85595 244507 94605
rect 248705 85595 248739 94605
rect 255697 93891 255731 98685
rect 255697 84235 255731 93721
rect 262505 86955 262539 99433
rect 234813 74579 234847 84133
rect 267013 82875 267047 102085
rect 280537 95251 280571 104805
rect 305285 102187 305319 106233
rect 309333 102459 309367 115209
rect 345213 114563 345247 124117
rect 347973 116059 348007 125545
rect 444205 118643 444239 125545
rect 313657 102459 313691 113101
rect 324697 104907 324731 106301
rect 342545 104975 342579 114461
rect 288633 86139 288667 99433
rect 327365 95251 327399 104805
rect 342545 95251 342579 104805
rect 345213 98719 345247 104805
rect 347973 96747 348007 106233
rect 434361 95251 434395 104805
rect 444113 99331 444147 106233
rect 309425 85595 309459 89777
rect 229293 64991 229327 74477
rect 240517 66351 240551 75837
rect 234813 55267 234847 64821
rect 239045 51051 239079 57885
rect 240333 55267 240367 64821
rect 244289 57987 244323 67541
rect 248797 66283 248831 75837
rect 262781 66283 262815 75837
rect 267105 67643 267139 77945
rect 255605 64719 255639 66181
rect 245945 48331 245979 57885
rect 267013 56627 267047 61081
rect 288725 57987 288759 73797
rect 291485 66283 291519 79305
rect 307953 74579 307987 84133
rect 313657 74579 313691 84133
rect 327365 77299 327399 86853
rect 343741 76007 343775 85493
rect 345213 75939 345247 93789
rect 434361 87159 434395 91749
rect 362969 77299 363003 86921
rect 305285 64923 305319 74409
rect 327365 66283 327399 67609
rect 343741 66283 343775 75837
rect 308045 64923 308079 66249
rect 254133 46971 254167 56525
rect 255605 45679 255639 55165
rect 261217 48331 261251 53125
rect 229293 38743 229327 41429
rect 234813 35955 234847 45509
rect 241805 29019 241839 44081
rect 245945 29019 245979 38573
rect 262873 37315 262907 46869
rect 267105 38675 267139 48229
rect 290013 45611 290047 55097
rect 324605 53091 324639 66181
rect 299857 48331 299891 51153
rect 336933 48331 336967 57885
rect 345213 56627 345247 66181
rect 347973 64923 348007 74477
rect 362969 70295 363003 77129
rect 435189 75939 435223 85493
rect 444113 77299 444147 86921
rect 434269 66351 434303 75837
rect 342545 46971 342579 51153
rect 261217 27659 261251 31773
rect 267013 27659 267047 37213
rect 280537 28883 280571 44489
rect 229201 8347 229235 17901
rect 231317 9707 231351 12529
rect 234721 11203 234755 12461
rect 234813 8959 234847 26197
rect 234905 16643 234939 26197
rect 238953 8347 238987 26197
rect 251373 18003 251407 27557
rect 290013 26299 290047 35853
rect 292773 26299 292807 30685
rect 305377 24871 305411 35853
rect 240241 8347 240275 17901
rect 241621 8347 241655 17901
rect 252753 9707 252787 22729
rect 254133 9707 254167 22729
rect 262597 19363 262631 24157
rect 299857 15215 299891 16677
rect 308137 12971 308171 19465
rect 324605 19363 324639 28917
rect 328561 27659 328595 31841
rect 345213 29019 345247 46869
rect 346593 45611 346627 51153
rect 347881 45679 347915 55165
rect 363153 48331 363187 57885
rect 435189 51051 435223 66181
rect 435281 38675 435315 48229
rect 444113 38675 444147 48229
rect 363153 29019 363187 38573
rect 434453 29087 434487 35037
rect 444113 29019 444147 31841
rect 290105 12223 290139 12461
rect 327273 9707 327307 19261
rect 328469 12359 328503 22729
rect 342453 9707 342487 27557
rect 345213 9707 345247 27557
rect 346409 16643 346443 26197
rect 363245 9707 363279 19261
rect 434637 18003 434671 27557
rect 435281 19363 435315 28917
rect 251189 8007 251223 8245
rect 254593 8007 254627 8245
rect 227637 6919 227671 7565
rect 2789 4743 2823 4845
rect 12449 4743 12483 4845
rect 19349 4743 19383 4845
rect 31769 4743 31803 4845
rect 41429 4743 41463 4845
rect 51089 4743 51123 4845
rect 60749 4743 60783 4845
rect 128369 4743 128403 4845
rect 138029 4743 138063 4845
rect 147689 4743 147723 4845
rect 157349 4743 157383 4845
rect 167009 4743 167043 4845
rect 173909 4743 173943 4845
rect 186329 4743 186363 4845
rect 195989 4743 196023 4845
rect 205649 4607 205683 4845
rect 215217 4607 215251 4845
rect 224233 4811 224267 4913
rect 306849 4777 307067 4811
rect 224141 4267 224175 4777
rect 306849 4743 306883 4777
rect 304825 4709 305101 4743
rect 304825 4607 304859 4709
rect 306941 4403 306975 4709
rect 307033 4471 307067 4777
rect 307033 4437 307125 4471
rect 284677 3927 284711 4097
rect 263609 3451 263643 3485
rect 263551 3417 263643 3451
rect 270543 3417 270601 3451
rect 280077 3247 280111 3417
rect 82921 2975 82955 3145
rect 280169 3111 280203 3281
rect 289737 3111 289771 3417
rect 290933 3383 290967 3485
rect 292439 3417 292589 3451
rect 302249 2975 302283 3417
rect 321569 3383 321603 3961
rect 326353 3383 326387 3485
rect 326445 3247 326479 3689
rect 330585 3519 330619 3757
rect 331263 3417 331413 3451
rect 326353 2975 326387 3213
rect 102793 2771 102827 2941
rect 326537 2907 326571 3009
rect 326629 2839 326663 2873
rect 326387 2805 326663 2839
rect 335277 2839 335311 3961
rect 344569 3587 344603 3893
rect 349905 3859 349939 4097
rect 393731 3893 393973 3927
rect 387165 3383 387199 3485
rect 388361 3247 388395 3893
rect 394065 3655 394099 4029
rect 394341 3383 394375 3757
rect 394433 3519 394467 3689
rect 394525 3451 394559 3757
rect 394341 3349 394433 3383
rect 400321 2975 400355 3417
rect 404921 3179 404955 3349
rect 422309 2975 422343 3213
rect 422401 2907 422435 3349
rect 427185 3247 427219 3349
rect 427093 3043 427127 3213
rect 432521 2907 432555 3213
rect 432613 3043 432647 3213
rect 441997 2975 442031 3213
rect 442181 2907 442215 3417
rect 442273 3247 442307 3553
rect 446689 2975 446723 3485
rect 456165 2907 456199 3485
rect 446321 2771 446355 2873
<< viali >>
rect 429577 684437 429611 684471
rect 559297 684437 559331 684471
rect 429577 666553 429611 666587
rect 494069 676141 494103 676175
rect 494069 666553 494103 666587
rect 559297 666553 559331 666587
rect 429393 608549 429427 608583
rect 429393 601681 429427 601715
rect 559113 608549 559147 608583
rect 559113 601681 559147 601715
rect 429577 598893 429611 598927
rect 429577 589305 429611 589339
rect 559297 598893 559331 598927
rect 559297 589305 559331 589339
rect 429485 579581 429519 579615
rect 429485 569925 429519 569959
rect 494069 579581 494103 579615
rect 494069 569925 494103 569959
rect 559297 579581 559331 579615
rect 559297 569925 559331 569959
rect 303997 563057 304031 563091
rect 303997 562921 304031 562955
rect 306941 562989 306975 563023
rect 307125 562921 307159 562955
rect 310437 562921 310471 562955
rect 311817 562921 311851 562955
rect 395353 562105 395387 562139
rect 395353 561017 395387 561051
rect 400229 560881 400263 560915
rect 400413 560881 400447 560915
rect 400321 560813 400355 560847
rect 400505 560813 400539 560847
rect 400321 560677 400355 560711
rect 400505 560677 400539 560711
rect 287805 560609 287839 560643
rect 400229 560609 400263 560643
rect 400413 560609 400447 560643
rect 372169 560541 372203 560575
rect 372353 560541 372387 560575
rect 400321 560541 400355 560575
rect 400505 560541 400539 560575
rect 372261 560473 372295 560507
rect 372445 560473 372479 560507
rect 400229 560473 400263 560507
rect 400413 560473 400447 560507
rect 372353 560405 372387 560439
rect 372537 560405 372571 560439
rect 400321 560405 400355 560439
rect 400505 560405 400539 560439
rect 372353 560269 372387 560303
rect 372537 560269 372571 560303
rect 400321 560269 400355 560303
rect 400505 560269 400539 560303
rect 287805 560201 287839 560235
rect 372169 560201 372203 560235
rect 372261 560201 372295 560235
rect 400321 560133 400355 560167
rect 400505 560133 400539 560167
rect 400321 559997 400355 560031
rect 400505 559997 400539 560031
rect 372169 559929 372203 559963
rect 372721 559929 372755 559963
rect 390569 559861 390603 559895
rect 390753 559861 390787 559895
rect 419549 559861 419583 559895
rect 419641 559861 419675 559895
rect 372169 559793 372203 559827
rect 372537 559793 372571 559827
rect 390661 559793 390695 559827
rect 390845 559793 390879 559827
rect 400229 559793 400263 559827
rect 400413 559793 400447 559827
rect 372261 559725 372295 559759
rect 372445 559725 372479 559759
rect 390661 559657 390695 559691
rect 390845 559657 390879 559691
rect 390569 559589 390603 559623
rect 390753 559589 390787 559623
rect 234629 559521 234663 559555
rect 372261 559521 372295 559555
rect 372353 559521 372387 559555
rect 229753 559453 229787 559487
rect 234629 559385 234663 559419
rect 236745 559453 236779 559487
rect 229753 559249 229787 559283
rect 236653 559317 236687 559351
rect 236745 559317 236779 559351
rect 236837 559385 236871 559419
rect 385325 559385 385359 559419
rect 396457 559385 396491 559419
rect 408325 559385 408359 559419
rect 408509 559385 408543 559419
rect 415869 559385 415903 559419
rect 301697 559317 301731 559351
rect 301881 559317 301915 559351
rect 321017 559317 321051 559351
rect 321201 559317 321235 559351
rect 340337 559317 340371 559351
rect 340521 559317 340555 559351
rect 369777 559317 369811 559351
rect 370053 559317 370087 559351
rect 385509 559317 385543 559351
rect 396273 559317 396307 559351
rect 408417 559317 408451 559351
rect 408601 559317 408635 559351
rect 416053 559317 416087 559351
rect 19257 559181 19291 559215
rect 9689 559113 9723 559147
rect 9689 558977 9723 559011
rect 20453 559181 20487 559215
rect 41521 559181 41555 559215
rect 38577 559113 38611 559147
rect 41337 559113 41371 559147
rect 48329 559181 48363 559215
rect 20453 559045 20487 559079
rect 29009 559045 29043 559079
rect 19257 558977 19291 559011
rect 29009 558909 29043 558943
rect 60841 559181 60875 559215
rect 48329 558977 48363 559011
rect 57897 559113 57931 559147
rect 60657 559113 60691 559147
rect 67649 559181 67683 559215
rect 57897 558977 57931 559011
rect 80161 559181 80195 559215
rect 67649 558977 67683 559011
rect 77217 559113 77251 559147
rect 79977 559113 80011 559147
rect 86969 559181 87003 559215
rect 77217 558977 77251 559011
rect 99481 559181 99515 559215
rect 86969 558977 87003 559011
rect 96537 559113 96571 559147
rect 99297 559113 99331 559147
rect 106289 559181 106323 559215
rect 96537 558977 96571 559011
rect 118801 559181 118835 559215
rect 106289 558977 106323 559011
rect 115857 559113 115891 559147
rect 118617 559113 118651 559147
rect 125609 559181 125643 559215
rect 115857 558977 115891 559011
rect 138121 559181 138155 559215
rect 125609 558977 125643 559011
rect 135177 559113 135211 559147
rect 137937 559113 137971 559147
rect 144929 559181 144963 559215
rect 135177 558977 135211 559011
rect 157441 559181 157475 559215
rect 144929 558977 144963 559011
rect 154497 559113 154531 559147
rect 157257 559113 157291 559147
rect 164249 559181 164283 559215
rect 154497 558977 154531 559011
rect 176761 559181 176795 559215
rect 164249 558977 164283 559011
rect 173817 559113 173851 559147
rect 176577 559113 176611 559147
rect 183569 559181 183603 559215
rect 173817 558977 173851 559011
rect 196081 559181 196115 559215
rect 183569 558977 183603 559011
rect 193137 559113 193171 559147
rect 195897 559113 195931 559147
rect 202889 559181 202923 559215
rect 193137 558977 193171 559011
rect 202889 558977 202923 559011
rect 212457 559113 212491 559147
rect 212457 558977 212491 559011
rect 38577 558909 38611 558943
rect 433441 338181 433475 338215
rect 425621 338113 425655 338147
rect 302157 338045 302191 338079
rect 259469 337977 259503 338011
rect 259377 337841 259411 337875
rect 253857 337773 253891 337807
rect 229845 337705 229879 337739
rect 229845 337501 229879 337535
rect 229937 337705 229971 337739
rect 229661 337433 229695 337467
rect 259469 337773 259503 337807
rect 294061 337977 294095 338011
rect 259377 337705 259411 337739
rect 287713 337637 287747 337671
rect 259561 337569 259595 337603
rect 259745 337569 259779 337603
rect 253857 337433 253891 337467
rect 89637 337297 89671 337331
rect 89637 337093 89671 337127
rect 99389 337297 99423 337331
rect 99389 336889 99423 336923
rect 108957 337297 108991 337331
rect 108957 336889 108991 336923
rect 118709 337297 118743 337331
rect 118709 336753 118743 336787
rect 128277 337297 128311 337331
rect 287713 337297 287747 337331
rect 267013 337229 267047 337263
rect 128277 336685 128311 336719
rect 239137 336685 239171 336719
rect 233525 334441 233559 334475
rect 233525 328457 233559 328491
rect 235089 331925 235123 331959
rect 235089 327097 235123 327131
rect 234813 327029 234847 327063
rect 267013 328457 267047 328491
rect 287437 334305 287471 334339
rect 297373 337909 297407 337943
rect 302157 337841 302191 337875
rect 303445 338045 303479 338079
rect 297373 337297 297407 337331
rect 299397 337229 299431 337263
rect 299397 337025 299431 337059
rect 299489 337229 299523 337263
rect 347973 338045 348007 338079
rect 336565 337977 336599 338011
rect 326261 337637 326295 337671
rect 326169 337365 326203 337399
rect 326261 337365 326295 337399
rect 326445 337569 326479 337603
rect 303445 337161 303479 337195
rect 326169 337161 326203 337195
rect 326353 337161 326387 337195
rect 341717 337841 341751 337875
rect 337945 337773 337979 337807
rect 340061 337705 340095 337739
rect 340061 337365 340095 337399
rect 340245 337569 340279 337603
rect 337945 337297 337979 337331
rect 340245 337297 340279 337331
rect 299489 337025 299523 337059
rect 326445 337025 326479 337059
rect 336565 337025 336599 337059
rect 336657 337025 336691 337059
rect 345673 337705 345707 337739
rect 345581 337501 345615 337535
rect 345489 337365 345523 337399
rect 341717 336957 341751 336991
rect 341809 337297 341843 337331
rect 336657 336889 336691 336923
rect 341809 336889 341843 336923
rect 326445 336753 326479 336787
rect 345673 337365 345707 337399
rect 345581 337025 345615 337059
rect 345489 336753 345523 336787
rect 324697 336685 324731 336719
rect 294061 329409 294095 329443
rect 319177 334169 319211 334203
rect 319177 328457 319211 328491
rect 343833 335529 343867 335563
rect 327457 331177 327491 331211
rect 327457 328457 327491 328491
rect 343833 328457 343867 328491
rect 353033 338045 353067 338079
rect 352849 337977 352883 338011
rect 352849 337841 352883 337875
rect 390569 338045 390603 338079
rect 381829 337977 381863 338011
rect 355149 337909 355183 337943
rect 353033 337501 353067 337535
rect 353493 337705 353527 337739
rect 353493 337501 353527 337535
rect 355149 337501 355183 337535
rect 356621 337705 356655 337739
rect 383577 337977 383611 338011
rect 383577 337773 383611 337807
rect 385969 337841 386003 337875
rect 381829 337501 381863 337535
rect 383853 337705 383887 337739
rect 356621 337433 356655 337467
rect 385969 337229 386003 337263
rect 388545 337841 388579 337875
rect 362877 337161 362911 337195
rect 383853 337161 383887 337195
rect 390569 337705 390603 337739
rect 396917 337977 396951 338011
rect 393237 337501 393271 337535
rect 425621 337705 425655 337739
rect 427001 338045 427035 338079
rect 396917 337433 396951 337467
rect 417065 337637 417099 337671
rect 417065 337433 417099 337467
rect 394525 337365 394559 337399
rect 394801 337365 394835 337399
rect 393237 337297 393271 337331
rect 432429 338045 432463 338079
rect 427001 337297 427035 337331
rect 427093 337909 427127 337943
rect 432429 337909 432463 337943
rect 432521 338045 432555 338079
rect 432521 337841 432555 337875
rect 432705 337841 432739 337875
rect 428289 337501 428323 337535
rect 388545 337161 388579 337195
rect 417433 337229 417467 337263
rect 427093 337229 427127 337263
rect 428105 337433 428139 337467
rect 362877 336957 362911 336991
rect 407773 337093 407807 337127
rect 417433 336957 417467 336991
rect 407773 336753 407807 336787
rect 433349 337773 433383 337807
rect 433349 337637 433383 337671
rect 437305 337841 437339 337875
rect 433441 337637 433475 337671
rect 437029 337705 437063 337739
rect 432705 337433 432739 337467
rect 435281 337569 435315 337603
rect 428289 337365 428323 337399
rect 428105 336685 428139 336719
rect 437029 337433 437063 337467
rect 442181 337841 442215 337875
rect 442181 337501 442215 337535
rect 442273 337841 442307 337875
rect 442917 337705 442951 337739
rect 446965 337705 446999 337739
rect 444941 337637 444975 337671
rect 442917 337501 442951 337535
rect 444757 337501 444791 337535
rect 445677 337637 445711 337671
rect 442273 337433 442307 337467
rect 445677 337365 445711 337399
rect 450001 337569 450035 337603
rect 437581 336753 437615 336787
rect 437765 336753 437799 336787
rect 447057 336753 447091 336787
rect 450001 336753 450035 336787
rect 437305 336617 437339 336651
rect 435281 336481 435315 336515
rect 347973 328457 348007 328491
rect 363245 328389 363279 328423
rect 324697 328321 324731 328355
rect 347973 328321 348007 328355
rect 287437 327097 287471 327131
rect 239137 318801 239171 318835
rect 347973 318801 348007 318835
rect 363245 318801 363279 318835
rect 234813 317441 234847 317475
rect 262689 318733 262723 318767
rect 250085 315945 250119 315979
rect 248797 311933 248831 311967
rect 235089 309077 235123 309111
rect 234905 307717 234939 307751
rect 229293 299557 229327 299591
rect 229293 298129 229327 298163
rect 235089 299489 235123 299523
rect 248797 299489 248831 299523
rect 292865 318733 292899 318767
rect 262689 312137 262723 312171
rect 287345 317373 287379 317407
rect 287345 311797 287379 311831
rect 290105 315877 290139 315911
rect 250085 299489 250119 299523
rect 267013 309009 267047 309043
rect 327457 318733 327491 318767
rect 292865 309145 292899 309179
rect 298477 317373 298511 317407
rect 290105 307785 290139 307819
rect 327457 309145 327491 309179
rect 342545 318733 342579 318767
rect 342545 309145 342579 309179
rect 345213 318733 345247 318767
rect 345213 309145 345247 309179
rect 434269 309077 434303 309111
rect 298477 307785 298511 307819
rect 347973 309009 348007 309043
rect 267013 299489 267047 299523
rect 305469 307717 305503 307751
rect 234905 298129 234939 298163
rect 262597 299421 262631 299455
rect 235089 298061 235123 298095
rect 240425 298061 240459 298095
rect 240425 288405 240459 288439
rect 241897 298061 241931 298095
rect 262597 289901 262631 289935
rect 287345 299421 287379 299455
rect 298477 299421 298511 299455
rect 287345 289833 287379 289867
rect 291485 298061 291519 298095
rect 241897 288405 241931 288439
rect 288725 289697 288759 289731
rect 235089 280177 235123 280211
rect 262505 288337 262539 288371
rect 229385 280109 229419 280143
rect 254225 280109 254259 280143
rect 229385 273105 229419 273139
rect 235089 278681 235123 278715
rect 229385 270453 229419 270487
rect 229385 263449 229419 263483
rect 239321 274057 239355 274091
rect 251465 273853 251499 273887
rect 239321 267733 239355 267767
rect 244289 270453 244323 270487
rect 235089 260865 235123 260899
rect 244289 260865 244323 260899
rect 245945 270453 245979 270487
rect 245945 260865 245979 260899
rect 316325 307717 316359 307751
rect 342453 307717 342487 307751
rect 305469 298129 305503 298163
rect 310805 298129 310839 298163
rect 316325 298129 316359 298163
rect 324605 299421 324639 299455
rect 310805 296701 310839 296735
rect 347973 299557 348007 299591
rect 434269 299489 434303 299523
rect 342453 298129 342487 298163
rect 327273 298061 327307 298095
rect 324605 289901 324639 289935
rect 325985 294661 326019 294695
rect 298477 289833 298511 289867
rect 325985 289833 326019 289867
rect 291485 288405 291519 288439
rect 316233 288473 316267 288507
rect 327273 288405 327307 288439
rect 345213 289765 345247 289799
rect 316233 287045 316267 287079
rect 288725 282829 288759 282863
rect 345213 280245 345247 280279
rect 434269 289765 434303 289799
rect 434269 280177 434303 280211
rect 262505 278817 262539 278851
rect 287345 280109 287379 280143
rect 254225 270521 254259 270555
rect 262505 278681 262539 278715
rect 251465 260865 251499 260899
rect 255605 270385 255639 270419
rect 290105 280109 290139 280143
rect 290105 272969 290139 273003
rect 298477 280109 298511 280143
rect 342545 280109 342579 280143
rect 324513 278681 324547 278715
rect 310713 273377 310747 273411
rect 298477 270589 298511 270623
rect 309425 273173 309459 273207
rect 287345 270521 287379 270555
rect 307953 270453 307987 270487
rect 288725 270385 288759 270419
rect 288725 263517 288759 263551
rect 262505 263449 262539 263483
rect 255605 260865 255639 260899
rect 229385 260797 229419 260831
rect 254225 260797 254259 260831
rect 229385 253793 229419 253827
rect 235089 259369 235123 259403
rect 251465 259369 251499 259403
rect 244289 251141 244323 251175
rect 235089 241485 235123 241519
rect 239137 249849 239171 249883
rect 244289 241485 244323 241519
rect 245945 251141 245979 251175
rect 262597 260797 262631 260831
rect 254225 251209 254259 251243
rect 255605 260729 255639 260763
rect 255605 251209 255639 251243
rect 262597 251209 262631 251243
rect 287345 260797 287379 260831
rect 290105 260797 290139 260831
rect 290105 252841 290139 252875
rect 291485 260797 291519 260831
rect 291485 251277 291519 251311
rect 298477 260797 298511 260831
rect 310713 267801 310747 267835
rect 309425 267733 309459 267767
rect 342545 270521 342579 270555
rect 363153 280109 363187 280143
rect 363153 270521 363187 270555
rect 324513 263449 324547 263483
rect 345213 270453 345247 270487
rect 345213 260933 345247 260967
rect 347973 270453 348007 270487
rect 347973 260933 348007 260967
rect 434269 270453 434303 270487
rect 434269 260865 434303 260899
rect 307953 258077 307987 258111
rect 324605 260797 324639 260831
rect 298477 251277 298511 251311
rect 310805 256649 310839 256683
rect 287345 251209 287379 251243
rect 251465 251073 251499 251107
rect 291485 251141 291519 251175
rect 245945 241485 245979 241519
rect 251465 241485 251499 241519
rect 291485 241485 291519 241519
rect 298477 251141 298511 251175
rect 298477 241485 298511 241519
rect 305193 251141 305227 251175
rect 307953 251141 307987 251175
rect 307953 244205 307987 244239
rect 305193 241485 305227 241519
rect 239137 240125 239171 240159
rect 251465 240125 251499 240159
rect 234905 240057 234939 240091
rect 288725 240057 288759 240091
rect 234905 230469 234939 230503
rect 251465 239989 251499 240023
rect 324605 251209 324639 251243
rect 342545 260797 342579 260831
rect 342545 251209 342579 251243
rect 363153 260797 363187 260831
rect 435281 260797 435315 260831
rect 435281 251277 435315 251311
rect 363153 251209 363187 251243
rect 327273 251141 327307 251175
rect 327273 242641 327307 242675
rect 345213 251141 345247 251175
rect 345213 241485 345247 241519
rect 347973 251141 348007 251175
rect 347973 241485 348007 241519
rect 434269 251141 434303 251175
rect 434269 241485 434303 241519
rect 435097 251141 435131 251175
rect 435097 241485 435131 241519
rect 310805 239989 310839 240023
rect 288725 231829 288759 231863
rect 251465 230469 251499 230503
rect 435097 224961 435131 224995
rect 435097 222173 435131 222207
rect 229293 220745 229327 220779
rect 229293 215237 229327 215271
rect 235089 220745 235123 220779
rect 291393 220745 291427 220779
rect 267013 215305 267047 215339
rect 267013 212517 267047 212551
rect 288725 215305 288759 215339
rect 288725 212517 288759 212551
rect 235089 211157 235123 211191
rect 239137 211089 239171 211123
rect 239137 202793 239171 202827
rect 267013 211089 267047 211123
rect 288817 205649 288851 205683
rect 434269 220745 434303 220779
rect 310897 219385 310931 219419
rect 308045 217413 308079 217447
rect 434269 215237 434303 215271
rect 310897 214557 310931 214591
rect 308045 212517 308079 212551
rect 343741 211089 343775 211123
rect 291393 202929 291427 202963
rect 305285 205649 305319 205683
rect 288817 202861 288851 202895
rect 305285 202861 305319 202895
rect 267013 202793 267047 202827
rect 343741 202793 343775 202827
rect 234813 201433 234847 201467
rect 240425 201433 240459 201467
rect 238861 198441 238895 198475
rect 238861 198033 238895 198067
rect 305285 201433 305319 201467
rect 240425 193137 240459 193171
rect 267013 200073 267047 200107
rect 234813 192253 234847 192287
rect 255605 191777 255639 191811
rect 255605 186269 255639 186303
rect 262597 191777 262631 191811
rect 298477 196061 298511 196095
rect 288725 195993 288759 196027
rect 288725 193205 288759 193239
rect 345029 201433 345063 201467
rect 310805 200073 310839 200107
rect 305285 195925 305319 195959
rect 308045 195993 308079 196027
rect 298477 193205 298511 193239
rect 308045 193205 308079 193239
rect 267013 190485 267047 190519
rect 288817 186337 288851 186371
rect 434453 195993 434487 196027
rect 434453 193205 434487 193239
rect 345029 192729 345063 192763
rect 316233 191845 316267 191879
rect 316233 190485 316267 190519
rect 310805 185589 310839 185623
rect 288817 183549 288851 183583
rect 262597 183481 262631 183515
rect 239137 182121 239171 182155
rect 255605 182121 255639 182155
rect 241805 178789 241839 178823
rect 241805 173893 241839 173927
rect 239137 173825 239171 173859
rect 327365 180761 327399 180795
rect 255605 172533 255639 172567
rect 310805 179333 310839 179367
rect 251373 171037 251407 171071
rect 241897 162809 241931 162843
rect 234997 161381 235031 161415
rect 234905 161313 234939 161347
rect 238861 159681 238895 159715
rect 238861 159341 238895 159375
rect 234997 151793 235031 151827
rect 239045 154649 239079 154683
rect 240425 154581 240459 154615
rect 240425 153289 240459 153323
rect 327365 171105 327399 171139
rect 310805 169745 310839 169779
rect 313565 171037 313599 171071
rect 287345 164169 287379 164203
rect 251373 161449 251407 161483
rect 261309 162809 261343 162843
rect 241897 153221 241931 153255
rect 261309 153221 261343 153255
rect 262505 162809 262539 162843
rect 305285 162809 305319 162843
rect 287345 154581 287379 154615
rect 288725 161381 288759 161415
rect 288725 153833 288759 153867
rect 262505 153221 262539 153255
rect 313565 161449 313599 161483
rect 324605 164169 324639 164203
rect 305285 153221 305319 153255
rect 308045 161381 308079 161415
rect 239045 151793 239079 151827
rect 240333 153153 240367 153187
rect 305285 153085 305319 153119
rect 240333 143565 240367 143599
rect 288817 149005 288851 149039
rect 251557 143497 251591 143531
rect 234905 140845 234939 140879
rect 239137 142069 239171 142103
rect 234813 140709 234847 140743
rect 234813 134589 234847 134623
rect 233433 132481 233467 132515
rect 239137 132481 239171 132515
rect 240333 142069 240367 142103
rect 287253 143497 287287 143531
rect 240333 132481 240367 132515
rect 241897 135201 241931 135235
rect 251557 135201 251591 135235
rect 262689 139349 262723 139383
rect 233433 131121 233467 131155
rect 235089 128333 235123 128367
rect 233433 125477 233467 125511
rect 241897 125613 241931 125647
rect 251465 133841 251499 133875
rect 444113 164169 444147 164203
rect 324605 154581 324639 154615
rect 343925 162809 343959 162843
rect 308045 151793 308079 151827
rect 327365 153493 327399 153527
rect 313657 150569 313691 150603
rect 313657 150433 313691 150467
rect 305285 142137 305319 142171
rect 309517 149005 309551 149039
rect 288817 139485 288851 139519
rect 343925 153221 343959 153255
rect 345213 162809 345247 162843
rect 327365 147577 327399 147611
rect 343833 148325 343867 148359
rect 309517 139417 309551 139451
rect 316325 142069 316359 142103
rect 287253 137785 287287 137819
rect 262689 129761 262723 129795
rect 267105 135201 267139 135235
rect 310805 133841 310839 133875
rect 267105 128265 267139 128299
rect 305377 132413 305411 132447
rect 251465 124185 251499 124219
rect 254225 125545 254259 125579
rect 235089 122825 235123 122859
rect 241897 124117 241931 124151
rect 233433 121465 233467 121499
rect 240333 122757 240367 122791
rect 234905 120037 234939 120071
rect 229293 115889 229327 115923
rect 229293 106301 229327 106335
rect 291577 124185 291611 124219
rect 261217 124117 261251 124151
rect 434453 159137 434487 159171
rect 444113 157301 444147 157335
rect 434453 154581 434487 154615
rect 444113 154513 444147 154547
rect 444113 144993 444147 145027
rect 345213 144925 345247 144959
rect 434453 143497 434487 143531
rect 434453 137921 434487 137955
rect 444113 143497 444147 143531
rect 343833 135269 343867 135303
rect 316325 132481 316359 132515
rect 327365 135201 327399 135235
rect 327365 128265 327399 128299
rect 444113 128265 444147 128299
rect 310805 124185 310839 124219
rect 328469 125545 328503 125579
rect 305377 122825 305411 122859
rect 291577 121465 291611 121499
rect 261217 118609 261251 118643
rect 262689 120037 262723 120071
rect 254225 115957 254259 115991
rect 241897 114529 241931 114563
rect 245945 115889 245979 115923
rect 245945 106301 245979 106335
rect 255605 114461 255639 114495
rect 240333 104873 240367 104907
rect 255605 104873 255639 104907
rect 234813 100725 234847 100759
rect 234905 100725 234939 100759
rect 241805 104805 241839 104839
rect 229293 96577 229327 96611
rect 251465 104805 251499 104839
rect 347973 125545 348007 125579
rect 328469 118609 328503 118643
rect 345213 124117 345247 124151
rect 298477 115889 298511 115923
rect 287345 114461 287379 114495
rect 287345 104873 287379 104907
rect 288725 114461 288759 114495
rect 298477 108817 298511 108851
rect 309333 115209 309367 115243
rect 288725 104873 288759 104907
rect 305285 106233 305319 106267
rect 262689 102153 262723 102187
rect 280537 104805 280571 104839
rect 267013 102085 267047 102119
rect 262505 99433 262539 99467
rect 251465 95285 251499 95319
rect 255697 98685 255731 98719
rect 241805 95217 241839 95251
rect 244473 94605 244507 94639
rect 234813 92021 234847 92055
rect 240517 93789 240551 93823
rect 229293 86989 229327 87023
rect 244473 85561 244507 85595
rect 248705 94605 248739 94639
rect 255697 93857 255731 93891
rect 248705 85561 248739 85595
rect 255697 93721 255731 93755
rect 240517 84201 240551 84235
rect 262505 86921 262539 86955
rect 255697 84201 255731 84235
rect 234813 84133 234847 84167
rect 444205 125545 444239 125579
rect 444205 118609 444239 118643
rect 347973 116025 348007 116059
rect 345213 114529 345247 114563
rect 342545 114461 342579 114495
rect 309333 102425 309367 102459
rect 313657 113101 313691 113135
rect 324697 106301 324731 106335
rect 342545 104941 342579 104975
rect 347973 106233 348007 106267
rect 324697 104873 324731 104907
rect 313657 102425 313691 102459
rect 327365 104805 327399 104839
rect 305285 102153 305319 102187
rect 280537 95217 280571 95251
rect 288633 99433 288667 99467
rect 327365 95217 327399 95251
rect 342545 104805 342579 104839
rect 345213 104805 345247 104839
rect 345213 98685 345247 98719
rect 444113 106233 444147 106267
rect 347973 96713 348007 96747
rect 434361 104805 434395 104839
rect 342545 95217 342579 95251
rect 444113 99297 444147 99331
rect 434361 95217 434395 95251
rect 345213 93789 345247 93823
rect 288633 86105 288667 86139
rect 309425 89777 309459 89811
rect 309425 85561 309459 85595
rect 327365 86853 327399 86887
rect 267013 82841 267047 82875
rect 307953 84133 307987 84167
rect 291485 79305 291519 79339
rect 267105 77945 267139 77979
rect 234813 74545 234847 74579
rect 240517 75837 240551 75871
rect 229293 74477 229327 74511
rect 248797 75837 248831 75871
rect 240517 66317 240551 66351
rect 244289 67541 244323 67575
rect 229293 64957 229327 64991
rect 234813 64821 234847 64855
rect 240333 64821 240367 64855
rect 234813 55233 234847 55267
rect 239045 57885 239079 57919
rect 248797 66249 248831 66283
rect 262781 75837 262815 75871
rect 267105 67609 267139 67643
rect 288725 73797 288759 73831
rect 262781 66249 262815 66283
rect 255605 66181 255639 66215
rect 255605 64685 255639 64719
rect 244289 57953 244323 57987
rect 267013 61081 267047 61115
rect 240333 55233 240367 55267
rect 245945 57885 245979 57919
rect 239045 51017 239079 51051
rect 307953 74545 307987 74579
rect 313657 84133 313691 84167
rect 327365 77265 327399 77299
rect 343741 85493 343775 85527
rect 343741 75973 343775 76007
rect 434361 91749 434395 91783
rect 434361 87125 434395 87159
rect 362969 86921 363003 86955
rect 444113 86921 444147 86955
rect 362969 77265 363003 77299
rect 435189 85493 435223 85527
rect 345213 75905 345247 75939
rect 362969 77129 363003 77163
rect 313657 74545 313691 74579
rect 343741 75837 343775 75871
rect 291485 66249 291519 66283
rect 305285 74409 305319 74443
rect 327365 67609 327399 67643
rect 305285 64889 305319 64923
rect 308045 66249 308079 66283
rect 327365 66249 327399 66283
rect 343741 66249 343775 66283
rect 347973 74477 348007 74511
rect 308045 64889 308079 64923
rect 324605 66181 324639 66215
rect 288725 57953 288759 57987
rect 267013 56593 267047 56627
rect 245945 48297 245979 48331
rect 254133 56525 254167 56559
rect 254133 46937 254167 46971
rect 255605 55165 255639 55199
rect 290013 55097 290047 55131
rect 261217 53125 261251 53159
rect 261217 48297 261251 48331
rect 267105 48229 267139 48263
rect 255605 45645 255639 45679
rect 262873 46869 262907 46903
rect 234813 45509 234847 45543
rect 229293 41429 229327 41463
rect 229293 38709 229327 38743
rect 234813 35921 234847 35955
rect 241805 44081 241839 44115
rect 241805 28985 241839 29019
rect 245945 38573 245979 38607
rect 345213 66181 345247 66215
rect 324605 53057 324639 53091
rect 336933 57885 336967 57919
rect 299857 51153 299891 51187
rect 299857 48297 299891 48331
rect 444113 77265 444147 77299
rect 435189 75905 435223 75939
rect 362969 70261 363003 70295
rect 434269 75837 434303 75871
rect 434269 66317 434303 66351
rect 347973 64889 348007 64923
rect 435189 66181 435223 66215
rect 345213 56593 345247 56627
rect 363153 57885 363187 57919
rect 347881 55165 347915 55199
rect 336933 48297 336967 48331
rect 342545 51153 342579 51187
rect 342545 46937 342579 46971
rect 346593 51153 346627 51187
rect 290013 45577 290047 45611
rect 345213 46869 345247 46903
rect 267105 38641 267139 38675
rect 280537 44489 280571 44523
rect 262873 37281 262907 37315
rect 267013 37213 267047 37247
rect 245945 28985 245979 29019
rect 261217 31773 261251 31807
rect 261217 27625 261251 27659
rect 280537 28849 280571 28883
rect 290013 35853 290047 35887
rect 267013 27625 267047 27659
rect 251373 27557 251407 27591
rect 234813 26197 234847 26231
rect 229201 17901 229235 17935
rect 231317 12529 231351 12563
rect 234721 12461 234755 12495
rect 234721 11169 234755 11203
rect 231317 9673 231351 9707
rect 234905 26197 234939 26231
rect 234905 16609 234939 16643
rect 238953 26197 238987 26231
rect 234813 8925 234847 8959
rect 229201 8313 229235 8347
rect 305377 35853 305411 35887
rect 290013 26265 290047 26299
rect 292773 30685 292807 30719
rect 292773 26265 292807 26299
rect 328561 31841 328595 31875
rect 305377 24837 305411 24871
rect 324605 28917 324639 28951
rect 262597 24157 262631 24191
rect 251373 17969 251407 18003
rect 252753 22729 252787 22763
rect 238953 8313 238987 8347
rect 240241 17901 240275 17935
rect 240241 8313 240275 8347
rect 241621 17901 241655 17935
rect 252753 9673 252787 9707
rect 254133 22729 254167 22763
rect 262597 19329 262631 19363
rect 308137 19465 308171 19499
rect 299857 16677 299891 16711
rect 299857 15181 299891 15215
rect 435189 51017 435223 51051
rect 363153 48297 363187 48331
rect 347881 45645 347915 45679
rect 435281 48229 435315 48263
rect 346593 45577 346627 45611
rect 435281 38641 435315 38675
rect 444113 48229 444147 48263
rect 444113 38641 444147 38675
rect 345213 28985 345247 29019
rect 363153 38573 363187 38607
rect 434453 35037 434487 35071
rect 434453 29053 434487 29087
rect 444113 31841 444147 31875
rect 363153 28985 363187 29019
rect 444113 28985 444147 29019
rect 328561 27625 328595 27659
rect 435281 28917 435315 28951
rect 342453 27557 342487 27591
rect 324605 19329 324639 19363
rect 328469 22729 328503 22763
rect 308137 12937 308171 12971
rect 327273 19261 327307 19295
rect 290105 12461 290139 12495
rect 290105 12189 290139 12223
rect 254133 9673 254167 9707
rect 328469 12325 328503 12359
rect 327273 9673 327307 9707
rect 342453 9673 342487 9707
rect 345213 27557 345247 27591
rect 434637 27557 434671 27591
rect 346409 26197 346443 26231
rect 346409 16609 346443 16643
rect 363245 19261 363279 19295
rect 345213 9673 345247 9707
rect 435281 19329 435315 19363
rect 434637 17969 434671 18003
rect 363245 9673 363279 9707
rect 241621 8313 241655 8347
rect 251189 8245 251223 8279
rect 251189 7973 251223 8007
rect 254593 8245 254627 8279
rect 254593 7973 254627 8007
rect 227637 7565 227671 7599
rect 227637 6885 227671 6919
rect 224233 4913 224267 4947
rect 2789 4845 2823 4879
rect 2789 4709 2823 4743
rect 12449 4845 12483 4879
rect 12449 4709 12483 4743
rect 19349 4845 19383 4879
rect 19349 4709 19383 4743
rect 31769 4845 31803 4879
rect 31769 4709 31803 4743
rect 41429 4845 41463 4879
rect 41429 4709 41463 4743
rect 51089 4845 51123 4879
rect 51089 4709 51123 4743
rect 60749 4845 60783 4879
rect 60749 4709 60783 4743
rect 128369 4845 128403 4879
rect 128369 4709 128403 4743
rect 138029 4845 138063 4879
rect 138029 4709 138063 4743
rect 147689 4845 147723 4879
rect 147689 4709 147723 4743
rect 157349 4845 157383 4879
rect 157349 4709 157383 4743
rect 167009 4845 167043 4879
rect 167009 4709 167043 4743
rect 173909 4845 173943 4879
rect 173909 4709 173943 4743
rect 186329 4845 186363 4879
rect 186329 4709 186363 4743
rect 195989 4845 196023 4879
rect 195989 4709 196023 4743
rect 205649 4845 205683 4879
rect 205649 4573 205683 4607
rect 215217 4845 215251 4879
rect 215217 4573 215251 4607
rect 224141 4777 224175 4811
rect 224233 4777 224267 4811
rect 305101 4709 305135 4743
rect 306849 4709 306883 4743
rect 306941 4709 306975 4743
rect 304825 4573 304859 4607
rect 307125 4437 307159 4471
rect 306941 4369 306975 4403
rect 224141 4233 224175 4267
rect 284677 4097 284711 4131
rect 349905 4097 349939 4131
rect 284677 3893 284711 3927
rect 321569 3961 321603 3995
rect 263609 3485 263643 3519
rect 290933 3485 290967 3519
rect 263517 3417 263551 3451
rect 270509 3417 270543 3451
rect 270601 3417 270635 3451
rect 280077 3417 280111 3451
rect 289737 3417 289771 3451
rect 280077 3213 280111 3247
rect 280169 3281 280203 3315
rect 82921 3145 82955 3179
rect 280169 3077 280203 3111
rect 292405 3417 292439 3451
rect 292589 3417 292623 3451
rect 302249 3417 302283 3451
rect 290933 3349 290967 3383
rect 289737 3077 289771 3111
rect 335277 3961 335311 3995
rect 330585 3757 330619 3791
rect 326445 3689 326479 3723
rect 321569 3349 321603 3383
rect 326353 3485 326387 3519
rect 326353 3349 326387 3383
rect 330585 3485 330619 3519
rect 331229 3417 331263 3451
rect 331413 3417 331447 3451
rect 82921 2941 82955 2975
rect 102793 2941 102827 2975
rect 302249 2941 302283 2975
rect 326353 3213 326387 3247
rect 326445 3213 326479 3247
rect 326353 2941 326387 2975
rect 326537 3009 326571 3043
rect 326537 2873 326571 2907
rect 326629 2873 326663 2907
rect 326353 2805 326387 2839
rect 344569 3893 344603 3927
rect 394065 4029 394099 4063
rect 349905 3825 349939 3859
rect 388361 3893 388395 3927
rect 393697 3893 393731 3927
rect 393973 3893 394007 3927
rect 344569 3553 344603 3587
rect 387165 3485 387199 3519
rect 387165 3349 387199 3383
rect 394065 3621 394099 3655
rect 394341 3757 394375 3791
rect 394525 3757 394559 3791
rect 394433 3689 394467 3723
rect 394433 3485 394467 3519
rect 442273 3553 442307 3587
rect 394525 3417 394559 3451
rect 400321 3417 400355 3451
rect 394433 3349 394467 3383
rect 388361 3213 388395 3247
rect 442181 3417 442215 3451
rect 404921 3349 404955 3383
rect 422401 3349 422435 3383
rect 404921 3145 404955 3179
rect 422309 3213 422343 3247
rect 400321 2941 400355 2975
rect 422309 2941 422343 2975
rect 427185 3349 427219 3383
rect 427093 3213 427127 3247
rect 427185 3213 427219 3247
rect 432521 3213 432555 3247
rect 427093 3009 427127 3043
rect 422401 2873 422435 2907
rect 432613 3213 432647 3247
rect 432613 3009 432647 3043
rect 441997 3213 442031 3247
rect 441997 2941 442031 2975
rect 432521 2873 432555 2907
rect 442273 3213 442307 3247
rect 446689 3485 446723 3519
rect 446689 2941 446723 2975
rect 456165 3485 456199 3519
rect 442181 2873 442215 2907
rect 446321 2873 446355 2907
rect 456165 2873 456199 2907
rect 335277 2805 335311 2839
rect 102793 2737 102827 2771
rect 446321 2737 446355 2771
<< metal1 >>
rect 328362 700952 328368 701004
rect 328420 700992 328426 701004
rect 478506 700992 478512 701004
rect 328420 700964 478512 700992
rect 328420 700952 328426 700964
rect 478506 700952 478512 700964
rect 478564 700952 478570 701004
rect 170306 700884 170312 700936
rect 170364 700924 170370 700936
rect 351914 700924 351920 700936
rect 170364 700896 351920 700924
rect 170364 700884 170370 700896
rect 351914 700884 351920 700896
rect 351972 700884 351978 700936
rect 154114 700816 154120 700868
rect 154172 700856 154178 700868
rect 356054 700856 356060 700868
rect 154172 700828 356060 700856
rect 154172 700816 154178 700828
rect 356054 700816 356060 700828
rect 356112 700816 356118 700868
rect 320082 700748 320088 700800
rect 320140 700788 320146 700800
rect 527174 700788 527180 700800
rect 320140 700760 527180 700788
rect 320140 700748 320146 700760
rect 527174 700748 527180 700760
rect 527232 700748 527238 700800
rect 137830 700680 137836 700732
rect 137888 700720 137894 700732
rect 353294 700720 353300 700732
rect 137888 700692 353300 700720
rect 137888 700680 137894 700692
rect 353294 700680 353300 700692
rect 353352 700680 353358 700732
rect 321462 700612 321468 700664
rect 321520 700652 321526 700664
rect 543458 700652 543464 700664
rect 321520 700624 543464 700652
rect 321520 700612 321526 700624
rect 543458 700612 543464 700624
rect 543516 700612 543522 700664
rect 105446 700544 105452 700596
rect 105504 700584 105510 700596
rect 357434 700584 357440 700596
rect 105504 700556 357440 700584
rect 105504 700544 105510 700556
rect 357434 700544 357440 700556
rect 357492 700544 357498 700596
rect 89162 700476 89168 700528
rect 89220 700516 89226 700528
rect 361574 700516 361580 700528
rect 89220 700488 361580 700516
rect 89220 700476 89226 700488
rect 361574 700476 361580 700488
rect 361632 700476 361638 700528
rect 72970 700408 72976 700460
rect 73028 700448 73034 700460
rect 358814 700448 358820 700460
rect 73028 700420 358820 700448
rect 73028 700408 73034 700420
rect 358814 700408 358820 700420
rect 358872 700408 358878 700460
rect 40494 700340 40500 700392
rect 40552 700380 40558 700392
rect 362954 700380 362960 700392
rect 40552 700352 362960 700380
rect 40552 700340 40558 700352
rect 362954 700340 362960 700352
rect 363012 700340 363018 700392
rect 24302 700272 24308 700324
rect 24360 700312 24366 700324
rect 367094 700312 367100 700324
rect 24360 700284 367100 700312
rect 24360 700272 24366 700284
rect 367094 700272 367100 700284
rect 367152 700272 367158 700324
rect 202782 700204 202788 700256
rect 202840 700244 202846 700256
rect 347866 700244 347872 700256
rect 202840 700216 347872 700244
rect 202840 700204 202846 700216
rect 347866 700204 347872 700216
rect 347924 700204 347930 700256
rect 348418 700204 348424 700256
rect 348476 700244 348482 700256
rect 364978 700244 364984 700256
rect 348476 700216 364984 700244
rect 348476 700204 348482 700216
rect 364978 700204 364984 700216
rect 365036 700204 365042 700256
rect 325602 700136 325608 700188
rect 325660 700176 325666 700188
rect 462314 700176 462320 700188
rect 325660 700148 462320 700176
rect 325660 700136 325666 700148
rect 462314 700136 462320 700148
rect 462372 700136 462378 700188
rect 218974 700068 218980 700120
rect 219032 700108 219038 700120
rect 349154 700108 349160 700120
rect 219032 700080 349160 700108
rect 219032 700068 219038 700080
rect 349154 700068 349160 700080
rect 349212 700068 349218 700120
rect 235166 700000 235172 700052
rect 235224 700040 235230 700052
rect 346394 700040 346400 700052
rect 235224 700012 346400 700040
rect 235224 700000 235230 700012
rect 346394 700000 346400 700012
rect 346452 700000 346458 700052
rect 333882 699932 333888 699984
rect 333940 699972 333946 699984
rect 413646 699972 413652 699984
rect 333940 699944 413652 699972
rect 333940 699932 333946 699944
rect 413646 699932 413652 699944
rect 413704 699932 413710 699984
rect 267642 699864 267648 699916
rect 267700 699904 267706 699916
rect 342254 699904 342260 699916
rect 267700 699876 342260 699904
rect 267700 699864 267706 699876
rect 342254 699864 342260 699876
rect 342312 699864 342318 699916
rect 331122 699796 331128 699848
rect 331180 699836 331186 699848
rect 397454 699836 397460 699848
rect 331180 699808 397460 699836
rect 331180 699796 331186 699808
rect 397454 699796 397460 699808
rect 397512 699796 397518 699848
rect 283834 699728 283840 699780
rect 283892 699768 283898 699780
rect 343634 699768 343640 699780
rect 283892 699740 343640 699768
rect 283892 699728 283898 699740
rect 343634 699728 343640 699740
rect 343692 699728 343698 699780
rect 300118 699660 300124 699712
rect 300176 699700 300182 699712
rect 300762 699700 300768 699712
rect 300176 699672 300768 699700
rect 300176 699660 300182 699672
rect 300762 699660 300768 699672
rect 300820 699660 300826 699712
rect 332502 699660 332508 699712
rect 332560 699700 332566 699712
rect 336734 699700 336740 699712
rect 332560 699672 336740 699700
rect 332560 699660 332566 699672
rect 336734 699660 336740 699672
rect 336792 699660 336798 699712
rect 339402 699660 339408 699712
rect 339460 699700 339466 699712
rect 348786 699700 348792 699712
rect 339460 699672 348792 699700
rect 339460 699660 339466 699672
rect 348786 699660 348792 699672
rect 348844 699660 348850 699712
rect 314562 696940 314568 696992
rect 314620 696980 314626 696992
rect 580166 696980 580172 696992
rect 314620 696952 580172 696980
rect 314620 696940 314626 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 429378 688576 429384 688628
rect 429436 688616 429442 688628
rect 429838 688616 429844 688628
rect 429436 688588 429844 688616
rect 429436 688576 429442 688588
rect 429838 688576 429844 688588
rect 429896 688576 429902 688628
rect 559098 688576 559104 688628
rect 559156 688616 559162 688628
rect 559650 688616 559656 688628
rect 559156 688588 559656 688616
rect 559156 688576 559162 688588
rect 559650 688576 559656 688588
rect 559708 688576 559714 688628
rect 429212 685936 429976 685964
rect 315942 685856 315948 685908
rect 316000 685896 316006 685908
rect 429212 685896 429240 685936
rect 316000 685868 429240 685896
rect 429948 685896 429976 685936
rect 552584 685936 559788 685964
rect 552584 685896 552612 685936
rect 429948 685868 552612 685896
rect 559760 685896 559788 685936
rect 580166 685896 580172 685908
rect 559760 685868 580172 685896
rect 316000 685856 316006 685868
rect 580166 685856 580172 685868
rect 580224 685856 580230 685908
rect 429286 684428 429292 684480
rect 429344 684468 429350 684480
rect 429565 684471 429623 684477
rect 429565 684468 429577 684471
rect 429344 684440 429577 684468
rect 429344 684428 429350 684440
rect 429565 684437 429577 684440
rect 429611 684437 429623 684471
rect 429565 684431 429623 684437
rect 559006 684428 559012 684480
rect 559064 684468 559070 684480
rect 559285 684471 559343 684477
rect 559285 684468 559297 684471
rect 559064 684440 559297 684468
rect 559064 684428 559070 684440
rect 559285 684437 559297 684440
rect 559331 684437 559343 684471
rect 559285 684431 559343 684437
rect 3510 681708 3516 681760
rect 3568 681748 3574 681760
rect 368474 681748 368480 681760
rect 3568 681720 368480 681748
rect 3568 681708 3574 681720
rect 368474 681708 368480 681720
rect 368532 681708 368538 681760
rect 494054 676172 494060 676184
rect 494015 676144 494060 676172
rect 494054 676132 494060 676144
rect 494112 676132 494118 676184
rect 311802 673480 311808 673532
rect 311860 673520 311866 673532
rect 580166 673520 580172 673532
rect 311860 673492 580172 673520
rect 311860 673480 311866 673492
rect 580166 673480 580172 673492
rect 580224 673480 580230 673532
rect 3418 667904 3424 667956
rect 3476 667944 3482 667956
rect 372614 667944 372620 667956
rect 3476 667916 372620 667944
rect 3476 667904 3482 667916
rect 372614 667904 372620 667916
rect 372672 667904 372678 667956
rect 429565 666587 429623 666593
rect 429565 666553 429577 666587
rect 429611 666584 429623 666587
rect 429654 666584 429660 666596
rect 429611 666556 429660 666584
rect 429611 666553 429623 666556
rect 429565 666547 429623 666553
rect 429654 666544 429660 666556
rect 429712 666544 429718 666596
rect 494057 666587 494115 666593
rect 494057 666553 494069 666587
rect 494103 666584 494115 666587
rect 494146 666584 494152 666596
rect 494103 666556 494152 666584
rect 494103 666553 494115 666556
rect 494057 666547 494115 666553
rect 494146 666544 494152 666556
rect 494204 666544 494210 666596
rect 559285 666587 559343 666593
rect 559285 666553 559297 666587
rect 559331 666584 559343 666587
rect 559374 666584 559380 666596
rect 559331 666556 559380 666584
rect 559331 666553 559343 666556
rect 559285 666547 559343 666553
rect 559374 666544 559380 666556
rect 559432 666544 559438 666596
rect 494054 654100 494060 654152
rect 494112 654140 494118 654152
rect 494238 654140 494244 654152
rect 494112 654112 494244 654140
rect 494112 654100 494118 654112
rect 494238 654100 494244 654112
rect 494296 654100 494302 654152
rect 3050 652740 3056 652792
rect 3108 652780 3114 652792
rect 371234 652780 371240 652792
rect 3108 652752 371240 652780
rect 3108 652740 3114 652752
rect 371234 652740 371240 652752
rect 371292 652740 371298 652792
rect 309042 650020 309048 650072
rect 309100 650060 309106 650072
rect 580166 650060 580172 650072
rect 309100 650032 580172 650060
rect 309100 650020 309106 650032
rect 580166 650020 580172 650032
rect 580224 650020 580230 650072
rect 429378 647232 429384 647284
rect 429436 647272 429442 647284
rect 429470 647272 429476 647284
rect 429436 647244 429476 647272
rect 429436 647232 429442 647244
rect 429470 647232 429476 647244
rect 429528 647232 429534 647284
rect 559098 647232 559104 647284
rect 559156 647272 559162 647284
rect 559190 647272 559196 647284
rect 559156 647244 559196 647272
rect 559156 647232 559162 647244
rect 559190 647232 559196 647244
rect 559248 647232 559254 647284
rect 429378 640364 429384 640416
rect 429436 640404 429442 640416
rect 429470 640404 429476 640416
rect 429436 640376 429476 640404
rect 429436 640364 429442 640376
rect 429470 640364 429476 640376
rect 429528 640364 429534 640416
rect 559098 640364 559104 640416
rect 559156 640404 559162 640416
rect 559190 640404 559196 640416
rect 559156 640376 559196 640404
rect 559156 640364 559162 640376
rect 559190 640364 559196 640376
rect 559248 640364 559254 640416
rect 310422 638936 310428 638988
rect 310480 638976 310486 638988
rect 580166 638976 580172 638988
rect 310480 638948 580172 638976
rect 310480 638936 310486 638948
rect 580166 638936 580172 638948
rect 580224 638936 580230 638988
rect 494054 634788 494060 634840
rect 494112 634828 494118 634840
rect 494238 634828 494244 634840
rect 494112 634800 494244 634828
rect 494112 634788 494118 634800
rect 494238 634788 494244 634800
rect 494296 634788 494302 634840
rect 429286 630640 429292 630692
rect 429344 630680 429350 630692
rect 429470 630680 429476 630692
rect 429344 630652 429476 630680
rect 429344 630640 429350 630652
rect 429470 630640 429476 630652
rect 429528 630640 429534 630692
rect 559006 630640 559012 630692
rect 559064 630680 559070 630692
rect 559190 630680 559196 630692
rect 559064 630652 559196 630680
rect 559064 630640 559070 630652
rect 559190 630640 559196 630652
rect 559248 630640 559254 630692
rect 306282 626560 306288 626612
rect 306340 626600 306346 626612
rect 580166 626600 580172 626612
rect 306340 626572 580172 626600
rect 306340 626560 306346 626572
rect 580166 626560 580172 626572
rect 580224 626560 580230 626612
rect 3418 623772 3424 623824
rect 3476 623812 3482 623824
rect 375374 623812 375380 623824
rect 3476 623784 375380 623812
rect 3476 623772 3482 623784
rect 375374 623772 375380 623784
rect 375432 623772 375438 623824
rect 494054 615476 494060 615528
rect 494112 615516 494118 615528
rect 494238 615516 494244 615528
rect 494112 615488 494244 615516
rect 494112 615476 494118 615488
rect 494238 615476 494244 615488
rect 494296 615476 494302 615528
rect 429286 611328 429292 611380
rect 429344 611368 429350 611380
rect 429470 611368 429476 611380
rect 429344 611340 429476 611368
rect 429344 611328 429350 611340
rect 429470 611328 429476 611340
rect 429528 611328 429534 611380
rect 559006 611328 559012 611380
rect 559064 611368 559070 611380
rect 559190 611368 559196 611380
rect 559064 611340 559196 611368
rect 559064 611328 559070 611340
rect 559190 611328 559196 611340
rect 559248 611328 559254 611380
rect 3418 609968 3424 610020
rect 3476 610008 3482 610020
rect 378134 610008 378140 610020
rect 3476 609980 378140 610008
rect 3476 609968 3482 609980
rect 378134 609968 378140 609980
rect 378192 609968 378198 610020
rect 429378 608580 429384 608592
rect 429339 608552 429384 608580
rect 429378 608540 429384 608552
rect 429436 608540 429442 608592
rect 559098 608580 559104 608592
rect 559059 608552 559104 608580
rect 559098 608540 559104 608552
rect 559156 608540 559162 608592
rect 302142 603100 302148 603152
rect 302200 603140 302206 603152
rect 580166 603140 580172 603152
rect 302200 603112 580172 603140
rect 302200 603100 302206 603112
rect 580166 603100 580172 603112
rect 580224 603100 580230 603152
rect 429381 601715 429439 601721
rect 429381 601681 429393 601715
rect 429427 601712 429439 601715
rect 429562 601712 429568 601724
rect 429427 601684 429568 601712
rect 429427 601681 429439 601684
rect 429381 601675 429439 601681
rect 429562 601672 429568 601684
rect 429620 601672 429626 601724
rect 559101 601715 559159 601721
rect 559101 601681 559113 601715
rect 559147 601712 559159 601715
rect 559282 601712 559288 601724
rect 559147 601684 559288 601712
rect 559147 601681 559159 601684
rect 559101 601675 559159 601681
rect 559282 601672 559288 601684
rect 559340 601672 559346 601724
rect 429562 598924 429568 598936
rect 429523 598896 429568 598924
rect 429562 598884 429568 598896
rect 429620 598884 429626 598936
rect 559282 598924 559288 598936
rect 559243 598896 559288 598924
rect 559282 598884 559288 598896
rect 559340 598884 559346 598936
rect 494054 596164 494060 596216
rect 494112 596204 494118 596216
rect 494238 596204 494244 596216
rect 494112 596176 494244 596204
rect 494112 596164 494118 596176
rect 494238 596164 494244 596176
rect 494296 596164 494302 596216
rect 3234 594804 3240 594856
rect 3292 594844 3298 594856
rect 376754 594844 376760 594856
rect 3292 594816 376760 594844
rect 3292 594804 3298 594816
rect 376754 594804 376760 594816
rect 376812 594804 376818 594856
rect 304902 592016 304908 592068
rect 304960 592056 304966 592068
rect 580166 592056 580172 592068
rect 304960 592028 580172 592056
rect 304960 592016 304966 592028
rect 580166 592016 580172 592028
rect 580224 592016 580230 592068
rect 429565 589339 429623 589345
rect 429565 589305 429577 589339
rect 429611 589336 429623 589339
rect 429654 589336 429660 589348
rect 429611 589308 429660 589336
rect 429611 589305 429623 589308
rect 429565 589299 429623 589305
rect 429654 589296 429660 589308
rect 429712 589296 429718 589348
rect 559285 589339 559343 589345
rect 559285 589305 559297 589339
rect 559331 589336 559343 589339
rect 559374 589336 559380 589348
rect 559331 589308 559380 589336
rect 559331 589305 559343 589308
rect 559285 589299 559343 589305
rect 559374 589296 559380 589308
rect 559432 589296 559438 589348
rect 425072 579720 429884 579748
rect 300670 579640 300676 579692
rect 300728 579680 300734 579692
rect 425072 579680 425100 579720
rect 300728 579652 425100 579680
rect 429856 579680 429884 579720
rect 493980 579720 494284 579748
rect 493980 579680 494008 579720
rect 429856 579652 494008 579680
rect 494256 579680 494284 579720
rect 555436 579720 559420 579748
rect 555436 579680 555464 579720
rect 494256 579652 555464 579680
rect 559392 579680 559420 579720
rect 580166 579680 580172 579692
rect 559392 579652 580172 579680
rect 300728 579640 300734 579652
rect 580166 579640 580172 579652
rect 580224 579640 580230 579692
rect 429473 579615 429531 579621
rect 429473 579581 429485 579615
rect 429519 579612 429531 579615
rect 429562 579612 429568 579624
rect 429519 579584 429568 579612
rect 429519 579581 429531 579584
rect 429473 579575 429531 579581
rect 429562 579572 429568 579584
rect 429620 579572 429626 579624
rect 494054 579612 494060 579624
rect 494015 579584 494060 579612
rect 494054 579572 494060 579584
rect 494112 579572 494118 579624
rect 559282 579612 559288 579624
rect 559243 579584 559288 579612
rect 559282 579572 559288 579584
rect 559340 579572 559346 579624
rect 429470 569956 429476 569968
rect 429431 569928 429476 569956
rect 429470 569916 429476 569928
rect 429528 569916 429534 569968
rect 494057 569959 494115 569965
rect 494057 569925 494069 569959
rect 494103 569956 494115 569959
rect 494238 569956 494244 569968
rect 494103 569928 494244 569956
rect 494103 569925 494115 569928
rect 494057 569919 494115 569925
rect 494238 569916 494244 569928
rect 494296 569916 494302 569968
rect 559285 569959 559343 569965
rect 559285 569925 559297 569959
rect 559331 569956 559343 569959
rect 559374 569956 559380 569968
rect 559331 569928 559380 569956
rect 559331 569925 559343 569928
rect 559285 569919 559343 569925
rect 559374 569916 559380 569928
rect 559432 569916 559438 569968
rect 3418 567196 3424 567248
rect 3476 567236 3482 567248
rect 380894 567236 380900 567248
rect 3476 567208 380900 567236
rect 3476 567196 3482 567208
rect 380894 567196 380900 567208
rect 380952 567196 380958 567248
rect 307754 565088 307760 565140
rect 307812 565128 307818 565140
rect 309042 565128 309048 565140
rect 307812 565100 309048 565128
rect 307812 565088 307818 565100
rect 309042 565088 309048 565100
rect 309100 565088 309106 565140
rect 309134 565088 309140 565140
rect 309192 565128 309198 565140
rect 310422 565128 310428 565140
rect 309192 565100 310428 565128
rect 309192 565088 309198 565100
rect 310422 565088 310428 565100
rect 310480 565088 310486 565140
rect 310514 565088 310520 565140
rect 310572 565128 310578 565140
rect 311802 565128 311808 565140
rect 310572 565100 311808 565128
rect 310572 565088 310578 565100
rect 311802 565088 311808 565100
rect 311860 565088 311866 565140
rect 313274 565088 313280 565140
rect 313332 565128 313338 565140
rect 314562 565128 314568 565140
rect 313332 565100 314568 565128
rect 313332 565088 313338 565100
rect 314562 565088 314568 565100
rect 314620 565088 314626 565140
rect 314654 565088 314660 565140
rect 314712 565128 314718 565140
rect 315942 565128 315948 565140
rect 314712 565100 315948 565128
rect 314712 565088 314718 565100
rect 315942 565088 315948 565100
rect 316000 565088 316006 565140
rect 327074 565088 327080 565140
rect 327132 565128 327138 565140
rect 328362 565128 328368 565140
rect 327132 565100 328368 565128
rect 327132 565088 327138 565100
rect 328362 565088 328368 565100
rect 328420 565088 328426 565140
rect 329834 565088 329840 565140
rect 329892 565128 329898 565140
rect 331122 565128 331128 565140
rect 329892 565100 331128 565128
rect 329892 565088 329898 565100
rect 331122 565088 331128 565100
rect 331180 565088 331186 565140
rect 332594 565088 332600 565140
rect 332652 565128 332658 565140
rect 333882 565128 333888 565140
rect 332652 565100 333888 565128
rect 332652 565088 332658 565100
rect 333882 565088 333888 565100
rect 333940 565088 333946 565140
rect 333974 563932 333980 563984
rect 334032 563972 334038 563984
rect 348418 563972 348424 563984
rect 334032 563944 348424 563972
rect 334032 563932 334038 563944
rect 348418 563932 348424 563944
rect 348476 563932 348482 563984
rect 300762 563864 300768 563916
rect 300820 563904 300826 563916
rect 340690 563904 340696 563916
rect 300820 563876 340696 563904
rect 300820 563864 300826 563876
rect 340690 563864 340696 563876
rect 340748 563864 340754 563916
rect 328454 563796 328460 563848
rect 328512 563836 328518 563848
rect 429470 563836 429476 563848
rect 328512 563808 429476 563836
rect 328512 563796 328518 563808
rect 429470 563796 429476 563808
rect 429528 563796 429534 563848
rect 323302 563728 323308 563780
rect 323360 563768 323366 563780
rect 494238 563768 494244 563780
rect 323360 563740 494244 563768
rect 323360 563728 323366 563740
rect 494238 563728 494244 563740
rect 494296 563728 494302 563780
rect 317506 563660 317512 563712
rect 317564 563700 317570 563712
rect 559374 563700 559380 563712
rect 317564 563672 559380 563700
rect 317564 563660 317570 563672
rect 559374 563660 559380 563672
rect 559432 563660 559438 563712
rect 303985 563091 304043 563097
rect 303985 563057 303997 563091
rect 304031 563088 304043 563091
rect 304031 563060 305040 563088
rect 304031 563057 304043 563060
rect 303985 563051 304043 563057
rect 289814 562980 289820 563032
rect 289872 563020 289878 563032
rect 305012 563020 305040 563060
rect 306929 563023 306987 563029
rect 306929 563020 306941 563023
rect 289872 562992 304948 563020
rect 305012 562992 306941 563020
rect 289872 562980 289878 562992
rect 298278 562912 298284 562964
rect 298336 562952 298342 562964
rect 303985 562955 304043 562961
rect 303985 562952 303997 562955
rect 298336 562924 303997 562952
rect 298336 562912 298342 562924
rect 303985 562921 303997 562924
rect 304031 562921 304043 562955
rect 304920 562952 304948 562992
rect 306929 562989 306941 562992
rect 306975 562989 306987 563023
rect 412082 563020 412088 563032
rect 306929 562983 306987 562989
rect 307036 562992 412088 563020
rect 307036 562952 307064 562992
rect 412082 562980 412088 562992
rect 412140 562980 412146 563032
rect 304920 562924 307064 562952
rect 307113 562955 307171 562961
rect 303985 562915 304043 562921
rect 307113 562921 307125 562955
rect 307159 562952 307171 562955
rect 310425 562955 310483 562961
rect 310425 562952 310437 562955
rect 307159 562924 310437 562952
rect 307159 562921 307171 562924
rect 307113 562915 307171 562921
rect 310425 562921 310437 562924
rect 310471 562921 310483 562955
rect 310425 562915 310483 562921
rect 310514 562912 310520 562964
rect 310572 562952 310578 562964
rect 311710 562952 311716 562964
rect 310572 562924 311716 562952
rect 310572 562912 310578 562924
rect 311710 562912 311716 562924
rect 311768 562912 311774 562964
rect 311805 562955 311863 562961
rect 311805 562921 311817 562955
rect 311851 562952 311863 562955
rect 450446 562952 450452 562964
rect 311851 562924 450452 562952
rect 311851 562921 311863 562924
rect 311805 562915 311863 562921
rect 450446 562912 450452 562924
rect 450504 562912 450510 562964
rect 255774 562844 255780 562896
rect 255832 562884 255838 562896
rect 286962 562884 286968 562896
rect 255832 562856 286968 562884
rect 255832 562844 255838 562856
rect 286962 562844 286968 562856
rect 287020 562844 287026 562896
rect 292482 562844 292488 562896
rect 292540 562884 292546 562896
rect 450354 562884 450360 562896
rect 292540 562856 450360 562884
rect 292540 562844 292546 562856
rect 450354 562844 450360 562856
rect 450412 562844 450418 562896
rect 284754 562776 284760 562828
rect 284812 562816 284818 562828
rect 451090 562816 451096 562828
rect 284812 562788 451096 562816
rect 284812 562776 284818 562788
rect 451090 562776 451096 562788
rect 451148 562776 451154 562828
rect 280890 562708 280896 562760
rect 280948 562748 280954 562760
rect 450722 562748 450728 562760
rect 280948 562720 450728 562748
rect 280948 562708 280954 562720
rect 450722 562708 450728 562720
rect 450780 562708 450786 562760
rect 278958 562640 278964 562692
rect 279016 562680 279022 562692
rect 450998 562680 451004 562692
rect 279016 562652 451004 562680
rect 279016 562640 279022 562652
rect 450998 562640 451004 562652
rect 451056 562640 451062 562692
rect 261570 562572 261576 562624
rect 261628 562612 261634 562624
rect 278774 562612 278780 562624
rect 261628 562584 278780 562612
rect 261628 562572 261634 562584
rect 278774 562572 278780 562584
rect 278832 562572 278838 562624
rect 286686 562572 286692 562624
rect 286744 562612 286750 562624
rect 462958 562612 462964 562624
rect 286744 562584 462964 562612
rect 286744 562572 286750 562584
rect 462958 562572 462964 562584
rect 463016 562572 463022 562624
rect 273162 562504 273168 562556
rect 273220 562544 273226 562556
rect 450630 562544 450636 562556
rect 273220 562516 450636 562544
rect 273220 562504 273226 562516
rect 450630 562504 450636 562516
rect 450688 562504 450694 562556
rect 259638 562436 259644 562488
rect 259696 562476 259702 562488
rect 580902 562476 580908 562488
rect 259696 562448 580908 562476
rect 259696 562436 259702 562448
rect 580902 562436 580908 562448
rect 580960 562436 580966 562488
rect 6546 562368 6552 562420
rect 6604 562408 6610 562420
rect 388898 562408 388904 562420
rect 6604 562380 388904 562408
rect 6604 562368 6610 562380
rect 388898 562368 388904 562380
rect 388956 562368 388962 562420
rect 3050 562300 3056 562352
rect 3108 562340 3114 562352
rect 386966 562340 386972 562352
rect 3108 562312 386972 562340
rect 3108 562300 3114 562312
rect 386966 562300 386972 562312
rect 387024 562300 387030 562352
rect 6638 562232 6644 562284
rect 6696 562272 6702 562284
rect 390830 562272 390836 562284
rect 6696 562244 390836 562272
rect 6696 562232 6702 562244
rect 390830 562232 390836 562244
rect 390888 562232 390894 562284
rect 3142 562164 3148 562216
rect 3200 562204 3206 562216
rect 392762 562204 392768 562216
rect 3200 562176 392768 562204
rect 3200 562164 3206 562176
rect 392762 562164 392768 562176
rect 392820 562164 392826 562216
rect 5442 562096 5448 562148
rect 5500 562136 5506 562148
rect 394694 562136 394700 562148
rect 5500 562108 394700 562136
rect 5500 562096 5506 562108
rect 394694 562096 394700 562108
rect 394752 562096 394758 562148
rect 395341 562139 395399 562145
rect 395341 562105 395353 562139
rect 395387 562136 395399 562139
rect 417878 562136 417884 562148
rect 395387 562108 417884 562136
rect 395387 562105 395399 562108
rect 395341 562099 395399 562105
rect 417878 562096 417884 562108
rect 417936 562096 417942 562148
rect 6454 562028 6460 562080
rect 6512 562068 6518 562080
rect 396626 562068 396632 562080
rect 6512 562040 396632 562068
rect 6512 562028 6518 562040
rect 396626 562028 396632 562040
rect 396684 562028 396690 562080
rect 3234 561960 3240 562012
rect 3292 562000 3298 562012
rect 398558 562000 398564 562012
rect 3292 561972 398564 562000
rect 3292 561960 3298 561972
rect 398558 561960 398564 561972
rect 398616 561960 398622 562012
rect 5350 561892 5356 561944
rect 5408 561932 5414 561944
rect 400490 561932 400496 561944
rect 5408 561904 400496 561932
rect 5408 561892 5414 561904
rect 400490 561892 400496 561904
rect 400548 561892 400554 561944
rect 6362 561824 6368 561876
rect 6420 561864 6426 561876
rect 402422 561864 402428 561876
rect 6420 561836 402428 561864
rect 6420 561824 6426 561836
rect 402422 561824 402428 561836
rect 402480 561824 402486 561876
rect 3326 561756 3332 561808
rect 3384 561796 3390 561808
rect 408218 561796 408224 561808
rect 3384 561768 408224 561796
rect 3384 561756 3390 561768
rect 408218 561756 408224 561768
rect 408276 561756 408282 561808
rect 6270 561688 6276 561740
rect 6328 561728 6334 561740
rect 414014 561728 414020 561740
rect 6328 561700 414020 561728
rect 6328 561688 6334 561700
rect 414014 561688 414020 561700
rect 414072 561688 414078 561740
rect 390646 561008 390652 561060
rect 390704 561048 390710 561060
rect 395341 561051 395399 561057
rect 395341 561048 395353 561051
rect 390704 561020 395353 561048
rect 390704 561008 390710 561020
rect 395341 561017 395353 561020
rect 395387 561017 395399 561051
rect 395341 561011 395399 561017
rect 4062 560940 4068 560992
rect 4120 560980 4126 560992
rect 289814 560980 289820 560992
rect 4120 560952 289820 560980
rect 4120 560940 4126 560952
rect 289814 560940 289820 560952
rect 289872 560940 289878 560992
rect 296346 560940 296352 560992
rect 296404 560980 296410 560992
rect 450814 560980 450820 560992
rect 296404 560952 450820 560980
rect 296404 560940 296410 560952
rect 450814 560940 450820 560952
rect 450872 560940 450878 560992
rect 290550 560872 290556 560924
rect 290608 560912 290614 560924
rect 400217 560915 400275 560921
rect 400217 560912 400229 560915
rect 290608 560884 400229 560912
rect 290608 560872 290614 560884
rect 400217 560881 400229 560884
rect 400263 560881 400275 560915
rect 400217 560875 400275 560881
rect 400401 560915 400459 560921
rect 400401 560881 400413 560915
rect 400447 560912 400459 560915
rect 451182 560912 451188 560924
rect 400447 560884 451188 560912
rect 400447 560881 400459 560884
rect 400401 560875 400459 560881
rect 451182 560872 451188 560884
rect 451240 560872 451246 560924
rect 282822 560804 282828 560856
rect 282880 560844 282886 560856
rect 400309 560847 400367 560853
rect 400309 560844 400321 560847
rect 282880 560816 400321 560844
rect 282880 560804 282886 560816
rect 400309 560813 400321 560816
rect 400355 560813 400367 560847
rect 400309 560807 400367 560813
rect 400493 560847 400551 560853
rect 400493 560813 400505 560847
rect 400539 560844 400551 560847
rect 450262 560844 450268 560856
rect 400539 560816 450268 560844
rect 400539 560813 400551 560816
rect 400493 560807 400551 560813
rect 450262 560804 450268 560816
rect 450320 560804 450326 560856
rect 277026 560736 277032 560788
rect 277084 560776 277090 560788
rect 400214 560776 400220 560788
rect 277084 560748 400220 560776
rect 277084 560736 277090 560748
rect 400214 560736 400220 560748
rect 400272 560736 400278 560788
rect 400582 560736 400588 560788
rect 400640 560776 400646 560788
rect 449618 560776 449624 560788
rect 400640 560748 449624 560776
rect 400640 560736 400646 560748
rect 449618 560736 449624 560748
rect 449676 560736 449682 560788
rect 271230 560668 271236 560720
rect 271288 560708 271294 560720
rect 400309 560711 400367 560717
rect 400309 560708 400321 560711
rect 271288 560680 400321 560708
rect 271288 560668 271294 560680
rect 400309 560677 400321 560680
rect 400355 560677 400367 560711
rect 400309 560671 400367 560677
rect 400493 560711 400551 560717
rect 400493 560677 400505 560711
rect 400539 560708 400551 560711
rect 450538 560708 450544 560720
rect 400539 560680 450544 560708
rect 400539 560677 400551 560680
rect 400493 560671 400551 560677
rect 450538 560668 450544 560680
rect 450596 560668 450602 560720
rect 286962 560600 286968 560652
rect 287020 560640 287026 560652
rect 287793 560643 287851 560649
rect 287793 560640 287805 560643
rect 287020 560612 287805 560640
rect 287020 560600 287026 560612
rect 287793 560609 287805 560612
rect 287839 560609 287851 560643
rect 287793 560603 287851 560609
rect 294414 560600 294420 560652
rect 294472 560640 294478 560652
rect 400217 560643 400275 560649
rect 400217 560640 400229 560643
rect 294472 560612 400229 560640
rect 294472 560600 294478 560612
rect 400217 560609 400229 560612
rect 400263 560609 400275 560643
rect 400217 560603 400275 560609
rect 400401 560643 400459 560649
rect 400401 560609 400413 560643
rect 400447 560640 400459 560643
rect 548518 560640 548524 560652
rect 400447 560612 548524 560640
rect 400447 560609 400459 560612
rect 400401 560603 400459 560609
rect 548518 560600 548524 560612
rect 548576 560600 548582 560652
rect 5258 560532 5264 560584
rect 5316 560572 5322 560584
rect 372157 560575 372215 560581
rect 372157 560572 372169 560575
rect 5316 560544 372169 560572
rect 5316 560532 5322 560544
rect 372157 560541 372169 560544
rect 372203 560541 372215 560575
rect 372157 560535 372215 560541
rect 372341 560575 372399 560581
rect 372341 560541 372353 560575
rect 372387 560572 372399 560575
rect 400309 560575 400367 560581
rect 400309 560572 400321 560575
rect 372387 560544 400321 560572
rect 372387 560541 372399 560544
rect 372341 560535 372399 560541
rect 400309 560541 400321 560544
rect 400355 560541 400367 560575
rect 400309 560535 400367 560541
rect 400493 560575 400551 560581
rect 400493 560541 400505 560575
rect 400539 560572 400551 560575
rect 410150 560572 410156 560584
rect 400539 560544 410156 560572
rect 400539 560541 400551 560544
rect 400493 560535 400551 560541
rect 410150 560532 410156 560544
rect 410208 560532 410214 560584
rect 411346 560532 411352 560584
rect 411404 560572 411410 560584
rect 424318 560572 424324 560584
rect 411404 560544 424324 560572
rect 411404 560532 411410 560544
rect 424318 560532 424324 560544
rect 424376 560532 424382 560584
rect 5166 560464 5172 560516
rect 5224 560504 5230 560516
rect 372249 560507 372307 560513
rect 372249 560504 372261 560507
rect 5224 560476 372261 560504
rect 5224 560464 5230 560476
rect 372249 560473 372261 560476
rect 372295 560473 372307 560507
rect 372249 560467 372307 560473
rect 372433 560507 372491 560513
rect 372433 560473 372445 560507
rect 372479 560504 372491 560507
rect 400217 560507 400275 560513
rect 400217 560504 400229 560507
rect 372479 560476 400229 560504
rect 372479 560473 372491 560476
rect 372433 560467 372491 560473
rect 400217 560473 400229 560476
rect 400263 560473 400275 560507
rect 400217 560467 400275 560473
rect 400401 560507 400459 560513
rect 400401 560473 400413 560507
rect 400447 560504 400459 560507
rect 421742 560504 421748 560516
rect 400447 560476 421748 560504
rect 400447 560473 400459 560476
rect 400401 560467 400459 560473
rect 421742 560464 421748 560476
rect 421800 560464 421806 560516
rect 4982 560396 4988 560448
rect 5040 560436 5046 560448
rect 372341 560439 372399 560445
rect 372341 560436 372353 560439
rect 5040 560408 372353 560436
rect 5040 560396 5046 560408
rect 372341 560405 372353 560408
rect 372387 560405 372399 560439
rect 372341 560399 372399 560405
rect 372525 560439 372583 560445
rect 372525 560405 372537 560439
rect 372571 560436 372583 560439
rect 400309 560439 400367 560445
rect 400309 560436 400321 560439
rect 372571 560408 400321 560436
rect 372571 560405 372583 560408
rect 372525 560399 372583 560405
rect 400309 560405 400321 560408
rect 400355 560405 400367 560439
rect 400309 560399 400367 560405
rect 400493 560439 400551 560445
rect 400493 560405 400505 560439
rect 400539 560436 400551 560439
rect 427538 560436 427544 560448
rect 400539 560408 427544 560436
rect 400539 560405 400551 560408
rect 400493 560399 400551 560405
rect 427538 560396 427544 560408
rect 427596 560396 427602 560448
rect 4798 560328 4804 560380
rect 4856 560368 4862 560380
rect 400214 560368 400220 560380
rect 4856 560340 400220 560368
rect 4856 560328 4862 560340
rect 400214 560328 400220 560340
rect 400272 560328 400278 560380
rect 400582 560328 400588 560380
rect 400640 560368 400646 560380
rect 433334 560368 433340 560380
rect 400640 560340 433340 560368
rect 400640 560328 400646 560340
rect 433334 560328 433340 560340
rect 433392 560328 433398 560380
rect 6178 560260 6184 560312
rect 6236 560300 6242 560312
rect 372341 560303 372399 560309
rect 372341 560300 372353 560303
rect 6236 560272 372353 560300
rect 6236 560260 6242 560272
rect 372341 560269 372353 560272
rect 372387 560269 372399 560303
rect 372341 560263 372399 560269
rect 372525 560303 372583 560309
rect 372525 560269 372537 560303
rect 372571 560300 372583 560303
rect 400309 560303 400367 560309
rect 400309 560300 400321 560303
rect 372571 560272 400321 560300
rect 372571 560269 372583 560272
rect 372525 560263 372583 560269
rect 400309 560269 400321 560272
rect 400355 560269 400367 560303
rect 400309 560263 400367 560269
rect 400493 560303 400551 560309
rect 400493 560269 400505 560303
rect 400539 560300 400551 560303
rect 439130 560300 439136 560312
rect 400539 560272 439136 560300
rect 400539 560269 400551 560272
rect 400493 560263 400551 560269
rect 439130 560260 439136 560272
rect 439188 560260 439194 560312
rect 287793 560235 287851 560241
rect 287793 560201 287805 560235
rect 287839 560232 287851 560235
rect 372157 560235 372215 560241
rect 372157 560232 372169 560235
rect 287839 560204 372169 560232
rect 287839 560201 287851 560204
rect 287793 560195 287851 560201
rect 372157 560201 372169 560204
rect 372203 560201 372215 560235
rect 372157 560195 372215 560201
rect 372249 560235 372307 560241
rect 372249 560201 372261 560235
rect 372295 560232 372307 560235
rect 400214 560232 400220 560244
rect 372295 560204 400220 560232
rect 372295 560201 372307 560204
rect 372249 560195 372307 560201
rect 400214 560192 400220 560204
rect 400272 560192 400278 560244
rect 400582 560192 400588 560244
rect 400640 560232 400646 560244
rect 579798 560232 579804 560244
rect 400640 560204 579804 560232
rect 400640 560192 400646 560204
rect 579798 560192 579804 560204
rect 579856 560192 579862 560244
rect 278774 560124 278780 560176
rect 278832 560164 278838 560176
rect 400309 560167 400367 560173
rect 400309 560164 400321 560167
rect 278832 560136 400321 560164
rect 278832 560124 278838 560136
rect 400309 560133 400321 560136
rect 400355 560133 400367 560167
rect 400309 560127 400367 560133
rect 400493 560167 400551 560173
rect 400493 560133 400505 560167
rect 400539 560164 400551 560167
rect 580074 560164 580080 560176
rect 400539 560136 580080 560164
rect 400539 560133 400551 560136
rect 400493 560127 400551 560133
rect 580074 560124 580080 560136
rect 580132 560124 580138 560176
rect 275094 560056 275100 560108
rect 275152 560096 275158 560108
rect 400214 560096 400220 560108
rect 275152 560068 400220 560096
rect 275152 560056 275158 560068
rect 400214 560056 400220 560068
rect 400272 560056 400278 560108
rect 400582 560056 400588 560108
rect 400640 560096 400646 560108
rect 579890 560096 579896 560108
rect 400640 560068 579896 560096
rect 400640 560056 400646 560068
rect 579890 560056 579896 560068
rect 579948 560056 579954 560108
rect 269666 559988 269672 560040
rect 269724 560028 269730 560040
rect 400309 560031 400367 560037
rect 400309 560028 400321 560031
rect 269724 560000 400321 560028
rect 269724 559988 269730 560000
rect 400309 559997 400321 560000
rect 400355 559997 400367 560031
rect 400309 559991 400367 559997
rect 400493 560031 400551 560037
rect 400493 559997 400505 560031
rect 400539 560028 400551 560031
rect 579982 560028 579988 560040
rect 400539 560000 579988 560028
rect 400539 559997 400551 560000
rect 400493 559991 400551 559997
rect 579982 559988 579988 560000
rect 580040 559988 580046 560040
rect 267642 559920 267648 559972
rect 267700 559960 267706 559972
rect 372157 559963 372215 559969
rect 372157 559960 372169 559963
rect 267700 559932 372169 559960
rect 267700 559920 267706 559932
rect 372157 559929 372169 559932
rect 372203 559929 372215 559963
rect 372157 559923 372215 559929
rect 372709 559963 372767 559969
rect 372709 559929 372721 559963
rect 372755 559960 372767 559963
rect 400214 559960 400220 559972
rect 372755 559932 400220 559960
rect 372755 559929 372767 559932
rect 372709 559923 372767 559929
rect 400214 559920 400220 559932
rect 400272 559920 400278 559972
rect 400582 559920 400588 559972
rect 400640 559960 400646 559972
rect 577590 559960 577596 559972
rect 400640 559932 577596 559960
rect 400640 559920 400646 559932
rect 577590 559920 577596 559932
rect 577648 559920 577654 559972
rect 265802 559852 265808 559904
rect 265860 559892 265866 559904
rect 372246 559892 372252 559904
rect 265860 559864 372252 559892
rect 265860 559852 265866 559864
rect 372246 559852 372252 559864
rect 372304 559852 372310 559904
rect 389082 559852 389088 559904
rect 389140 559892 389146 559904
rect 390557 559895 390615 559901
rect 390557 559892 390569 559895
rect 389140 559864 390569 559892
rect 389140 559852 389146 559864
rect 390557 559861 390569 559864
rect 390603 559861 390615 559895
rect 390557 559855 390615 559861
rect 390741 559895 390799 559901
rect 390741 559861 390753 559895
rect 390787 559892 390799 559895
rect 400306 559892 400312 559904
rect 390787 559864 400312 559892
rect 390787 559861 390799 559864
rect 390741 559855 390799 559861
rect 400306 559852 400312 559864
rect 400364 559852 400370 559904
rect 400674 559852 400680 559904
rect 400732 559892 400738 559904
rect 409874 559892 409880 559904
rect 400732 559864 409880 559892
rect 400732 559852 400738 559864
rect 409874 559852 409880 559864
rect 409932 559852 409938 559904
rect 419350 559852 419356 559904
rect 419408 559892 419414 559904
rect 419537 559895 419595 559901
rect 419537 559892 419549 559895
rect 419408 559864 419549 559892
rect 419408 559852 419414 559864
rect 419537 559861 419549 559864
rect 419583 559861 419595 559895
rect 419537 559855 419595 559861
rect 419629 559895 419687 559901
rect 419629 559861 419641 559895
rect 419675 559892 419687 559895
rect 577498 559892 577504 559904
rect 419675 559864 577504 559892
rect 419675 559861 419687 559864
rect 419629 559855 419687 559861
rect 577498 559852 577504 559864
rect 577556 559852 577562 559904
rect 263594 559784 263600 559836
rect 263652 559824 263658 559836
rect 372157 559827 372215 559833
rect 372157 559824 372169 559827
rect 263652 559796 372169 559824
rect 263652 559784 263658 559796
rect 372157 559793 372169 559796
rect 372203 559793 372215 559827
rect 372157 559787 372215 559793
rect 372525 559827 372583 559833
rect 372525 559793 372537 559827
rect 372571 559824 372583 559827
rect 390649 559827 390707 559833
rect 390649 559824 390661 559827
rect 372571 559796 390661 559824
rect 372571 559793 372583 559796
rect 372525 559787 372583 559793
rect 390649 559793 390661 559796
rect 390695 559793 390707 559827
rect 390649 559787 390707 559793
rect 390833 559827 390891 559833
rect 390833 559793 390845 559827
rect 390879 559824 390891 559827
rect 400217 559827 400275 559833
rect 400217 559824 400229 559827
rect 390879 559796 400229 559824
rect 390879 559793 390891 559796
rect 390833 559787 390891 559793
rect 400217 559793 400229 559796
rect 400263 559793 400275 559827
rect 400217 559787 400275 559793
rect 400401 559827 400459 559833
rect 400401 559793 400413 559827
rect 400447 559824 400459 559827
rect 580166 559824 580172 559836
rect 400447 559796 580172 559824
rect 400447 559793 400459 559796
rect 400401 559787 400459 559793
rect 580166 559784 580172 559796
rect 580224 559784 580230 559836
rect 3878 559716 3884 559768
rect 3936 559756 3942 559768
rect 372249 559759 372307 559765
rect 372249 559756 372261 559759
rect 3936 559728 372261 559756
rect 3936 559716 3942 559728
rect 372249 559725 372261 559728
rect 372295 559725 372307 559759
rect 372249 559719 372307 559725
rect 372433 559759 372491 559765
rect 372433 559725 372445 559759
rect 372479 559756 372491 559759
rect 390554 559756 390560 559768
rect 372479 559728 390560 559756
rect 372479 559725 372491 559728
rect 372433 559719 372491 559725
rect 390554 559716 390560 559728
rect 390612 559716 390618 559768
rect 258074 559648 258080 559700
rect 258132 559688 258138 559700
rect 390649 559691 390707 559697
rect 390649 559688 390661 559691
rect 258132 559660 390661 559688
rect 258132 559648 258138 559660
rect 390649 559657 390661 559660
rect 390695 559657 390707 559691
rect 390649 559651 390707 559657
rect 390833 559691 390891 559697
rect 390833 559657 390845 559691
rect 390879 559688 390891 559691
rect 580718 559688 580724 559700
rect 390879 559660 580724 559688
rect 390879 559657 390891 559660
rect 390833 559651 390891 559657
rect 580718 559648 580724 559660
rect 580776 559648 580782 559700
rect 248782 559620 248788 559632
rect 240152 559592 248788 559620
rect 234617 559555 234675 559561
rect 234617 559521 234629 559555
rect 234663 559552 234675 559555
rect 234663 559524 239444 559552
rect 234663 559521 234675 559524
rect 234617 559515 234675 559521
rect 229741 559487 229799 559493
rect 229741 559453 229753 559487
rect 229787 559484 229799 559487
rect 236733 559487 236791 559493
rect 236733 559484 236745 559487
rect 229787 559456 236745 559484
rect 229787 559453 229799 559456
rect 229741 559447 229799 559453
rect 236733 559453 236745 559456
rect 236779 559453 236791 559487
rect 236733 559447 236791 559453
rect 5534 559376 5540 559428
rect 5592 559416 5598 559428
rect 234617 559419 234675 559425
rect 234617 559416 234629 559419
rect 5592 559388 234629 559416
rect 5592 559376 5598 559388
rect 234617 559385 234629 559388
rect 234663 559385 234675 559419
rect 234617 559379 234675 559385
rect 236825 559419 236883 559425
rect 236825 559385 236837 559419
rect 236871 559416 236883 559419
rect 239416 559416 239444 559524
rect 240152 559496 240180 559592
rect 248782 559580 248788 559592
rect 248840 559580 248846 559632
rect 252186 559580 252192 559632
rect 252244 559620 252250 559632
rect 390557 559623 390615 559629
rect 390557 559620 390569 559623
rect 252244 559592 390569 559620
rect 252244 559580 252250 559592
rect 390557 559589 390569 559592
rect 390603 559589 390615 559623
rect 390557 559583 390615 559589
rect 390741 559623 390799 559629
rect 390741 559589 390753 559623
rect 390787 559620 390799 559623
rect 580626 559620 580632 559632
rect 390787 559592 580632 559620
rect 390787 559589 390799 559592
rect 390741 559583 390799 559589
rect 580626 559580 580632 559592
rect 580684 559580 580690 559632
rect 246482 559512 246488 559564
rect 246540 559552 246546 559564
rect 372249 559555 372307 559561
rect 372249 559552 372261 559555
rect 246540 559524 372261 559552
rect 246540 559512 246546 559524
rect 372249 559521 372261 559524
rect 372295 559521 372307 559555
rect 372249 559515 372307 559521
rect 372341 559555 372399 559561
rect 372341 559521 372353 559555
rect 372387 559552 372399 559555
rect 580442 559552 580448 559564
rect 372387 559524 580448 559552
rect 372387 559521 372399 559524
rect 372341 559515 372399 559521
rect 580442 559512 580448 559524
rect 580500 559512 580506 559564
rect 240134 559444 240140 559496
rect 240192 559444 240198 559496
rect 240594 559444 240600 559496
rect 240652 559484 240658 559496
rect 580258 559484 580264 559496
rect 240652 559456 580264 559484
rect 240652 559444 240658 559456
rect 580258 559444 580264 559456
rect 580316 559444 580322 559496
rect 384850 559416 384856 559428
rect 236871 559388 239352 559416
rect 239416 559388 384856 559416
rect 236871 559385 236883 559388
rect 236825 559379 236883 559385
rect 3694 559308 3700 559360
rect 3752 559348 3758 559360
rect 236641 559351 236699 559357
rect 236641 559348 236653 559351
rect 3752 559320 236653 559348
rect 3752 559308 3758 559320
rect 236641 559317 236653 559320
rect 236687 559317 236699 559351
rect 236641 559311 236699 559317
rect 236733 559351 236791 559357
rect 236733 559317 236745 559351
rect 236779 559317 236791 559351
rect 239324 559348 239352 559388
rect 384850 559376 384856 559388
rect 384908 559376 384914 559428
rect 385313 559419 385371 559425
rect 385313 559416 385325 559419
rect 384960 559388 385325 559416
rect 301685 559351 301743 559357
rect 301685 559348 301697 559351
rect 239324 559320 301697 559348
rect 236733 559311 236791 559317
rect 301685 559317 301697 559320
rect 301731 559317 301743 559351
rect 301685 559311 301743 559317
rect 301869 559351 301927 559357
rect 301869 559317 301881 559351
rect 301915 559348 301927 559351
rect 321005 559351 321063 559357
rect 321005 559348 321017 559351
rect 301915 559320 321017 559348
rect 301915 559317 301927 559320
rect 301869 559311 301927 559317
rect 321005 559317 321017 559320
rect 321051 559317 321063 559351
rect 321005 559311 321063 559317
rect 321189 559351 321247 559357
rect 321189 559317 321201 559351
rect 321235 559348 321247 559351
rect 340325 559351 340383 559357
rect 340325 559348 340337 559351
rect 321235 559320 340337 559348
rect 321235 559317 321247 559320
rect 321189 559311 321247 559317
rect 340325 559317 340337 559320
rect 340371 559317 340383 559351
rect 340325 559311 340383 559317
rect 340509 559351 340567 559357
rect 340509 559317 340521 559351
rect 340555 559348 340567 559351
rect 369765 559351 369823 559357
rect 369765 559348 369777 559351
rect 340555 559320 369777 559348
rect 340555 559317 340567 559320
rect 340509 559311 340567 559317
rect 369765 559317 369777 559320
rect 369811 559317 369823 559351
rect 369765 559311 369823 559317
rect 229741 559283 229799 559289
rect 229741 559280 229753 559283
rect 224880 559252 229753 559280
rect 19245 559215 19303 559221
rect 19245 559181 19257 559215
rect 19291 559212 19303 559215
rect 20441 559215 20499 559221
rect 20441 559212 20453 559215
rect 19291 559184 20453 559212
rect 19291 559181 19303 559184
rect 19245 559175 19303 559181
rect 20441 559181 20453 559184
rect 20487 559181 20499 559215
rect 20441 559175 20499 559181
rect 41509 559215 41567 559221
rect 41509 559181 41521 559215
rect 41555 559212 41567 559215
rect 48317 559215 48375 559221
rect 48317 559212 48329 559215
rect 41555 559184 48329 559212
rect 41555 559181 41567 559184
rect 41509 559175 41567 559181
rect 48317 559181 48329 559184
rect 48363 559181 48375 559215
rect 48317 559175 48375 559181
rect 60829 559215 60887 559221
rect 60829 559181 60841 559215
rect 60875 559212 60887 559215
rect 67637 559215 67695 559221
rect 67637 559212 67649 559215
rect 60875 559184 67649 559212
rect 60875 559181 60887 559184
rect 60829 559175 60887 559181
rect 67637 559181 67649 559184
rect 67683 559181 67695 559215
rect 67637 559175 67695 559181
rect 80149 559215 80207 559221
rect 80149 559181 80161 559215
rect 80195 559212 80207 559215
rect 86957 559215 87015 559221
rect 86957 559212 86969 559215
rect 80195 559184 86969 559212
rect 80195 559181 80207 559184
rect 80149 559175 80207 559181
rect 86957 559181 86969 559184
rect 87003 559181 87015 559215
rect 86957 559175 87015 559181
rect 99469 559215 99527 559221
rect 99469 559181 99481 559215
rect 99515 559212 99527 559215
rect 106277 559215 106335 559221
rect 106277 559212 106289 559215
rect 99515 559184 106289 559212
rect 99515 559181 99527 559184
rect 99469 559175 99527 559181
rect 106277 559181 106289 559184
rect 106323 559181 106335 559215
rect 106277 559175 106335 559181
rect 118789 559215 118847 559221
rect 118789 559181 118801 559215
rect 118835 559212 118847 559215
rect 125597 559215 125655 559221
rect 125597 559212 125609 559215
rect 118835 559184 125609 559212
rect 118835 559181 118847 559184
rect 118789 559175 118847 559181
rect 125597 559181 125609 559184
rect 125643 559181 125655 559215
rect 125597 559175 125655 559181
rect 138109 559215 138167 559221
rect 138109 559181 138121 559215
rect 138155 559212 138167 559215
rect 144917 559215 144975 559221
rect 144917 559212 144929 559215
rect 138155 559184 144929 559212
rect 138155 559181 138167 559184
rect 138109 559175 138167 559181
rect 144917 559181 144929 559184
rect 144963 559181 144975 559215
rect 144917 559175 144975 559181
rect 157429 559215 157487 559221
rect 157429 559181 157441 559215
rect 157475 559212 157487 559215
rect 164237 559215 164295 559221
rect 164237 559212 164249 559215
rect 157475 559184 164249 559212
rect 157475 559181 157487 559184
rect 157429 559175 157487 559181
rect 164237 559181 164249 559184
rect 164283 559181 164295 559215
rect 164237 559175 164295 559181
rect 176749 559215 176807 559221
rect 176749 559181 176761 559215
rect 176795 559212 176807 559215
rect 183557 559215 183615 559221
rect 183557 559212 183569 559215
rect 176795 559184 183569 559212
rect 176795 559181 176807 559184
rect 176749 559175 176807 559181
rect 183557 559181 183569 559184
rect 183603 559181 183615 559215
rect 183557 559175 183615 559181
rect 196069 559215 196127 559221
rect 196069 559181 196081 559215
rect 196115 559212 196127 559215
rect 202877 559215 202935 559221
rect 202877 559212 202889 559215
rect 196115 559184 202889 559212
rect 196115 559181 196127 559184
rect 196069 559175 196127 559181
rect 202877 559181 202889 559184
rect 202923 559181 202935 559215
rect 224880 559212 224908 559252
rect 229741 559249 229753 559252
rect 229787 559249 229799 559283
rect 236748 559280 236776 559311
rect 369854 559308 369860 559360
rect 369912 559308 369918 559360
rect 370041 559351 370099 559357
rect 370041 559317 370053 559351
rect 370087 559348 370099 559351
rect 384960 559348 384988 559388
rect 385313 559385 385325 559388
rect 385359 559385 385371 559419
rect 385313 559379 385371 559385
rect 396350 559376 396356 559428
rect 396408 559376 396414 559428
rect 396445 559419 396503 559425
rect 396445 559385 396457 559419
rect 396491 559416 396503 559419
rect 408313 559419 408371 559425
rect 408313 559416 408325 559419
rect 396491 559388 408325 559416
rect 396491 559385 396503 559388
rect 396445 559379 396503 559385
rect 408313 559385 408325 559388
rect 408359 559385 408371 559419
rect 408313 559379 408371 559385
rect 408497 559419 408555 559425
rect 408497 559385 408509 559419
rect 408543 559385 408555 559419
rect 415857 559419 415915 559425
rect 415857 559416 415869 559419
rect 408497 559379 408555 559385
rect 415688 559388 415869 559416
rect 370087 559320 384988 559348
rect 370087 559317 370099 559320
rect 370041 559311 370099 559317
rect 385126 559308 385132 559360
rect 385184 559308 385190 559360
rect 385497 559351 385555 559357
rect 385497 559317 385509 559351
rect 385543 559348 385555 559351
rect 396074 559348 396080 559360
rect 385543 559320 396080 559348
rect 385543 559317 385555 559320
rect 385497 559311 385555 559317
rect 396074 559308 396080 559320
rect 396132 559308 396138 559360
rect 396261 559351 396319 559357
rect 396261 559317 396273 559351
rect 396307 559317 396319 559351
rect 396368 559348 396396 559376
rect 408405 559351 408463 559357
rect 408405 559348 408417 559351
rect 396368 559320 408417 559348
rect 396261 559311 396319 559317
rect 408405 559317 408417 559320
rect 408451 559317 408463 559351
rect 408405 559311 408463 559317
rect 369872 559280 369900 559308
rect 236748 559252 369900 559280
rect 385144 559280 385172 559308
rect 396276 559280 396304 559311
rect 385144 559252 396304 559280
rect 408512 559280 408540 559379
rect 408589 559351 408647 559357
rect 408589 559317 408601 559351
rect 408635 559348 408647 559351
rect 415688 559348 415716 559388
rect 415857 559385 415869 559388
rect 415903 559385 415915 559419
rect 434990 559416 434996 559428
rect 415857 559379 415915 559385
rect 415964 559388 434996 559416
rect 408635 559320 415716 559348
rect 408635 559317 408647 559320
rect 408589 559311 408647 559317
rect 415964 559280 415992 559388
rect 434990 559376 434996 559388
rect 435048 559376 435054 559428
rect 416041 559351 416099 559357
rect 416041 559317 416053 559351
rect 416087 559348 416099 559351
rect 431126 559348 431132 559360
rect 416087 559320 431132 559348
rect 416087 559317 416099 559320
rect 416041 559311 416099 559317
rect 431126 559308 431132 559320
rect 431184 559308 431190 559360
rect 408512 559252 415992 559280
rect 229741 559243 229799 559249
rect 202877 559175 202935 559181
rect 215312 559184 224908 559212
rect 3510 559104 3516 559156
rect 3568 559144 3574 559156
rect 9677 559147 9735 559153
rect 9677 559144 9689 559147
rect 3568 559116 9689 559144
rect 3568 559104 3574 559116
rect 9677 559113 9689 559116
rect 9723 559113 9735 559147
rect 9677 559107 9735 559113
rect 38565 559147 38623 559153
rect 38565 559113 38577 559147
rect 38611 559144 38623 559147
rect 41325 559147 41383 559153
rect 41325 559144 41337 559147
rect 38611 559116 41337 559144
rect 38611 559113 38623 559116
rect 38565 559107 38623 559113
rect 41325 559113 41337 559116
rect 41371 559113 41383 559147
rect 41325 559107 41383 559113
rect 57885 559147 57943 559153
rect 57885 559113 57897 559147
rect 57931 559144 57943 559147
rect 60645 559147 60703 559153
rect 60645 559144 60657 559147
rect 57931 559116 60657 559144
rect 57931 559113 57943 559116
rect 57885 559107 57943 559113
rect 60645 559113 60657 559116
rect 60691 559113 60703 559147
rect 60645 559107 60703 559113
rect 77205 559147 77263 559153
rect 77205 559113 77217 559147
rect 77251 559144 77263 559147
rect 79965 559147 80023 559153
rect 79965 559144 79977 559147
rect 77251 559116 79977 559144
rect 77251 559113 77263 559116
rect 77205 559107 77263 559113
rect 79965 559113 79977 559116
rect 80011 559113 80023 559147
rect 79965 559107 80023 559113
rect 96525 559147 96583 559153
rect 96525 559113 96537 559147
rect 96571 559144 96583 559147
rect 99285 559147 99343 559153
rect 99285 559144 99297 559147
rect 96571 559116 99297 559144
rect 96571 559113 96583 559116
rect 96525 559107 96583 559113
rect 99285 559113 99297 559116
rect 99331 559113 99343 559147
rect 99285 559107 99343 559113
rect 115845 559147 115903 559153
rect 115845 559113 115857 559147
rect 115891 559144 115903 559147
rect 118605 559147 118663 559153
rect 118605 559144 118617 559147
rect 115891 559116 118617 559144
rect 115891 559113 115903 559116
rect 115845 559107 115903 559113
rect 118605 559113 118617 559116
rect 118651 559113 118663 559147
rect 118605 559107 118663 559113
rect 135165 559147 135223 559153
rect 135165 559113 135177 559147
rect 135211 559144 135223 559147
rect 137925 559147 137983 559153
rect 137925 559144 137937 559147
rect 135211 559116 137937 559144
rect 135211 559113 135223 559116
rect 135165 559107 135223 559113
rect 137925 559113 137937 559116
rect 137971 559113 137983 559147
rect 137925 559107 137983 559113
rect 154485 559147 154543 559153
rect 154485 559113 154497 559147
rect 154531 559144 154543 559147
rect 157245 559147 157303 559153
rect 157245 559144 157257 559147
rect 154531 559116 157257 559144
rect 154531 559113 154543 559116
rect 154485 559107 154543 559113
rect 157245 559113 157257 559116
rect 157291 559113 157303 559147
rect 157245 559107 157303 559113
rect 173805 559147 173863 559153
rect 173805 559113 173817 559147
rect 173851 559144 173863 559147
rect 176565 559147 176623 559153
rect 176565 559144 176577 559147
rect 173851 559116 176577 559144
rect 173851 559113 173863 559116
rect 173805 559107 173863 559113
rect 176565 559113 176577 559116
rect 176611 559113 176623 559147
rect 176565 559107 176623 559113
rect 193125 559147 193183 559153
rect 193125 559113 193137 559147
rect 193171 559144 193183 559147
rect 195885 559147 195943 559153
rect 195885 559144 195897 559147
rect 193171 559116 195897 559144
rect 193171 559113 193183 559116
rect 193125 559107 193183 559113
rect 195885 559113 195897 559116
rect 195931 559113 195943 559147
rect 195885 559107 195943 559113
rect 212445 559147 212503 559153
rect 212445 559113 212457 559147
rect 212491 559144 212503 559147
rect 215312 559144 215340 559184
rect 212491 559116 215340 559144
rect 212491 559113 212503 559116
rect 212445 559107 212503 559113
rect 20441 559079 20499 559085
rect 20441 559045 20453 559079
rect 20487 559076 20499 559079
rect 28997 559079 29055 559085
rect 28997 559076 29009 559079
rect 20487 559048 29009 559076
rect 20487 559045 20499 559048
rect 20441 559039 20499 559045
rect 28997 559045 29009 559048
rect 29043 559045 29055 559079
rect 28997 559039 29055 559045
rect 9677 559011 9735 559017
rect 9677 558977 9689 559011
rect 9723 559008 9735 559011
rect 19245 559011 19303 559017
rect 19245 559008 19257 559011
rect 9723 558980 19257 559008
rect 9723 558977 9735 558980
rect 9677 558971 9735 558977
rect 19245 558977 19257 558980
rect 19291 558977 19303 559011
rect 19245 558971 19303 558977
rect 48317 559011 48375 559017
rect 48317 558977 48329 559011
rect 48363 559008 48375 559011
rect 57885 559011 57943 559017
rect 57885 559008 57897 559011
rect 48363 558980 57897 559008
rect 48363 558977 48375 558980
rect 48317 558971 48375 558977
rect 57885 558977 57897 558980
rect 57931 558977 57943 559011
rect 57885 558971 57943 558977
rect 67637 559011 67695 559017
rect 67637 558977 67649 559011
rect 67683 559008 67695 559011
rect 77205 559011 77263 559017
rect 77205 559008 77217 559011
rect 67683 558980 77217 559008
rect 67683 558977 67695 558980
rect 67637 558971 67695 558977
rect 77205 558977 77217 558980
rect 77251 558977 77263 559011
rect 77205 558971 77263 558977
rect 86957 559011 87015 559017
rect 86957 558977 86969 559011
rect 87003 559008 87015 559011
rect 96525 559011 96583 559017
rect 96525 559008 96537 559011
rect 87003 558980 96537 559008
rect 87003 558977 87015 558980
rect 86957 558971 87015 558977
rect 96525 558977 96537 558980
rect 96571 558977 96583 559011
rect 96525 558971 96583 558977
rect 106277 559011 106335 559017
rect 106277 558977 106289 559011
rect 106323 559008 106335 559011
rect 115845 559011 115903 559017
rect 115845 559008 115857 559011
rect 106323 558980 115857 559008
rect 106323 558977 106335 558980
rect 106277 558971 106335 558977
rect 115845 558977 115857 558980
rect 115891 558977 115903 559011
rect 115845 558971 115903 558977
rect 125597 559011 125655 559017
rect 125597 558977 125609 559011
rect 125643 559008 125655 559011
rect 135165 559011 135223 559017
rect 135165 559008 135177 559011
rect 125643 558980 135177 559008
rect 125643 558977 125655 558980
rect 125597 558971 125655 558977
rect 135165 558977 135177 558980
rect 135211 558977 135223 559011
rect 135165 558971 135223 558977
rect 144917 559011 144975 559017
rect 144917 558977 144929 559011
rect 144963 559008 144975 559011
rect 154485 559011 154543 559017
rect 154485 559008 154497 559011
rect 144963 558980 154497 559008
rect 144963 558977 144975 558980
rect 144917 558971 144975 558977
rect 154485 558977 154497 558980
rect 154531 558977 154543 559011
rect 154485 558971 154543 558977
rect 164237 559011 164295 559017
rect 164237 558977 164249 559011
rect 164283 559008 164295 559011
rect 173805 559011 173863 559017
rect 173805 559008 173817 559011
rect 164283 558980 173817 559008
rect 164283 558977 164295 558980
rect 164237 558971 164295 558977
rect 173805 558977 173817 558980
rect 173851 558977 173863 559011
rect 173805 558971 173863 558977
rect 183557 559011 183615 559017
rect 183557 558977 183569 559011
rect 183603 559008 183615 559011
rect 193125 559011 193183 559017
rect 193125 559008 193137 559011
rect 183603 558980 193137 559008
rect 183603 558977 183615 558980
rect 183557 558971 183615 558977
rect 193125 558977 193137 558980
rect 193171 558977 193183 559011
rect 193125 558971 193183 558977
rect 202877 559011 202935 559017
rect 202877 558977 202889 559011
rect 202923 559008 202935 559011
rect 212445 559011 212503 559017
rect 212445 559008 212457 559011
rect 202923 558980 212457 559008
rect 202923 558977 202935 558980
rect 202877 558971 202935 558977
rect 212445 558977 212457 558980
rect 212491 558977 212503 559011
rect 212445 558971 212503 558977
rect 28997 558943 29055 558949
rect 28997 558909 29009 558943
rect 29043 558940 29055 558943
rect 38565 558943 38623 558949
rect 38565 558940 38577 558943
rect 29043 558912 38577 558940
rect 29043 558909 29055 558912
rect 28997 558903 29055 558909
rect 38565 558909 38577 558912
rect 38611 558909 38623 558943
rect 38565 558903 38623 558909
rect 450814 557472 450820 557524
rect 450872 557512 450878 557524
rect 579706 557512 579712 557524
rect 450872 557484 579712 557512
rect 450872 557472 450878 557484
rect 579706 557472 579712 557484
rect 579764 557472 579770 557524
rect 450262 557268 450268 557320
rect 450320 557308 450326 557320
rect 450906 557308 450912 557320
rect 450320 557280 450912 557308
rect 450320 557268 450326 557280
rect 450906 557268 450912 557280
rect 450964 557268 450970 557320
rect 450354 557132 450360 557184
rect 450412 557172 450418 557184
rect 451090 557172 451096 557184
rect 450412 557144 451096 557172
rect 450412 557132 450418 557144
rect 451090 557132 451096 557144
rect 451148 557132 451154 557184
rect 2774 553052 2780 553104
rect 2832 553092 2838 553104
rect 5534 553092 5540 553104
rect 2832 553064 5540 553092
rect 2832 553052 2838 553064
rect 5534 553052 5540 553064
rect 5592 553052 5598 553104
rect 579798 552644 579804 552696
rect 579856 552684 579862 552696
rect 580810 552684 580816 552696
rect 579856 552656 580816 552684
rect 579856 552644 579862 552656
rect 580810 552644 580816 552656
rect 580868 552644 580874 552696
rect 450446 546388 450452 546440
rect 450504 546428 450510 546440
rect 579798 546428 579804 546440
rect 450504 546400 579804 546428
rect 450504 546388 450510 546400
rect 579798 546388 579804 546400
rect 579856 546388 579862 546440
rect 548518 534012 548524 534064
rect 548576 534052 548582 534064
rect 579798 534052 579804 534064
rect 548576 534024 579804 534052
rect 548576 534012 548582 534024
rect 579798 534012 579804 534024
rect 579856 534012 579862 534064
rect 451182 510552 451188 510604
rect 451240 510592 451246 510604
rect 579798 510592 579804 510604
rect 451240 510564 579804 510592
rect 451240 510552 451246 510564
rect 579798 510552 579804 510564
rect 579856 510552 579862 510604
rect 451090 499468 451096 499520
rect 451148 499508 451154 499520
rect 579798 499508 579804 499520
rect 451148 499480 579804 499508
rect 451148 499468 451154 499480
rect 579798 499468 579804 499480
rect 579856 499468 579862 499520
rect 3050 495524 3056 495576
rect 3108 495564 3114 495576
rect 6638 495564 6644 495576
rect 3108 495536 6644 495564
rect 3108 495524 3114 495536
rect 6638 495524 6644 495536
rect 6696 495524 6702 495576
rect 3050 481108 3056 481160
rect 3108 481148 3114 481160
rect 6546 481148 6552 481160
rect 3108 481120 6552 481148
rect 3108 481108 3114 481120
rect 6546 481108 6552 481120
rect 6604 481108 6610 481160
rect 450998 463632 451004 463684
rect 451056 463672 451062 463684
rect 579798 463672 579804 463684
rect 451056 463644 579804 463672
rect 451056 463632 451062 463644
rect 579798 463632 579804 463644
rect 579856 463632 579862 463684
rect 462958 452548 462964 452600
rect 463016 452588 463022 452600
rect 579798 452588 579804 452600
rect 463016 452560 579804 452588
rect 463016 452548 463022 452560
rect 579798 452548 579804 452560
rect 579856 452548 579862 452600
rect 450906 440172 450912 440224
rect 450964 440212 450970 440224
rect 579798 440212 579804 440224
rect 450964 440184 579804 440212
rect 450964 440172 450970 440184
rect 579798 440172 579804 440184
rect 579856 440172 579862 440224
rect 3142 438676 3148 438728
rect 3200 438716 3206 438728
rect 6454 438716 6460 438728
rect 3200 438688 6460 438716
rect 3200 438676 3206 438688
rect 6454 438676 6460 438688
rect 6512 438676 6518 438728
rect 2774 424668 2780 424720
rect 2832 424708 2838 424720
rect 5442 424708 5448 424720
rect 2832 424680 5448 424708
rect 2832 424668 2838 424680
rect 5442 424668 5448 424680
rect 5500 424668 5506 424720
rect 450814 416712 450820 416764
rect 450872 416752 450878 416764
rect 579798 416752 579804 416764
rect 450872 416724 579804 416752
rect 450872 416712 450878 416724
rect 579798 416712 579804 416724
rect 579856 416712 579862 416764
rect 450722 405628 450728 405680
rect 450780 405668 450786 405680
rect 579798 405668 579804 405680
rect 450780 405640 579804 405668
rect 450780 405628 450786 405640
rect 579798 405628 579804 405640
rect 579856 405628 579862 405680
rect 449710 393252 449716 393304
rect 449768 393292 449774 393304
rect 579798 393292 579804 393304
rect 449768 393264 579804 393292
rect 449768 393252 449774 393264
rect 579798 393252 579804 393264
rect 579856 393252 579862 393304
rect 3142 380604 3148 380656
rect 3200 380644 3206 380656
rect 6362 380644 6368 380656
rect 3200 380616 6368 380644
rect 3200 380604 3206 380616
rect 6362 380604 6368 380616
rect 6420 380604 6426 380656
rect 450630 369792 450636 369844
rect 450688 369832 450694 369844
rect 579798 369832 579804 369844
rect 450688 369804 579804 369832
rect 450688 369792 450694 369804
rect 579798 369792 579804 369804
rect 579856 369792 579862 369844
rect 2774 366936 2780 366988
rect 2832 366976 2838 366988
rect 5350 366976 5356 366988
rect 2832 366948 5356 366976
rect 2832 366936 2838 366948
rect 5350 366936 5356 366948
rect 5408 366936 5414 366988
rect 450538 346332 450544 346384
rect 450596 346372 450602 346384
rect 579890 346372 579896 346384
rect 450596 346344 579896 346372
rect 450596 346332 450602 346344
rect 579890 346332 579896 346344
rect 579948 346332 579954 346384
rect 363046 340076 363052 340128
rect 363104 340116 363110 340128
rect 363874 340116 363880 340128
rect 363104 340088 363880 340116
rect 363104 340076 363110 340088
rect 363874 340076 363880 340088
rect 363932 340076 363938 340128
rect 345198 339056 345204 339108
rect 345256 339096 345262 339108
rect 345750 339096 345756 339108
rect 345256 339068 345756 339096
rect 345256 339056 345262 339068
rect 345750 339056 345756 339068
rect 345808 339056 345814 339108
rect 270586 338376 270592 338428
rect 270644 338416 270650 338428
rect 271230 338416 271236 338428
rect 270644 338388 271236 338416
rect 270644 338376 270650 338388
rect 271230 338376 271236 338388
rect 271288 338376 271294 338428
rect 433429 338215 433487 338221
rect 433429 338212 433441 338215
rect 432340 338184 433441 338212
rect 239122 338104 239128 338156
rect 239180 338144 239186 338156
rect 239858 338144 239864 338156
rect 239180 338116 239864 338144
rect 239180 338104 239186 338116
rect 239858 338104 239864 338116
rect 239916 338104 239922 338156
rect 425609 338147 425667 338153
rect 425609 338113 425621 338147
rect 425655 338144 425667 338147
rect 425655 338116 427124 338144
rect 425655 338113 425667 338116
rect 425609 338107 425667 338113
rect 79318 338036 79324 338088
rect 79376 338076 79382 338088
rect 258258 338076 258264 338088
rect 79376 338048 258264 338076
rect 79376 338036 79382 338048
rect 258258 338036 258264 338048
rect 258316 338036 258322 338088
rect 292482 338036 292488 338088
rect 292540 338076 292546 338088
rect 302145 338079 302203 338085
rect 302145 338076 302157 338079
rect 292540 338048 302157 338076
rect 292540 338036 292546 338048
rect 302145 338045 302157 338048
rect 302191 338045 302203 338079
rect 302145 338039 302203 338045
rect 303433 338079 303491 338085
rect 303433 338045 303445 338079
rect 303479 338076 303491 338079
rect 341794 338076 341800 338088
rect 303479 338048 341800 338076
rect 303479 338045 303491 338048
rect 303433 338039 303491 338045
rect 341794 338036 341800 338048
rect 341852 338036 341858 338088
rect 347961 338079 348019 338085
rect 347961 338045 347973 338079
rect 348007 338076 348019 338079
rect 348234 338076 348240 338088
rect 348007 338048 348240 338076
rect 348007 338045 348019 338048
rect 347961 338039 348019 338045
rect 348234 338036 348240 338048
rect 348292 338036 348298 338088
rect 349798 338036 349804 338088
rect 349856 338076 349862 338088
rect 353021 338079 353079 338085
rect 349856 338048 352972 338076
rect 349856 338036 349862 338048
rect 71038 337968 71044 338020
rect 71096 338008 71102 338020
rect 250162 338008 250168 338020
rect 71096 337980 250168 338008
rect 71096 337968 71102 337980
rect 250162 337968 250168 337980
rect 250220 337968 250226 338020
rect 259457 338011 259515 338017
rect 259457 337977 259469 338011
rect 259503 338008 259515 338011
rect 263594 338008 263600 338020
rect 259503 337980 263600 338008
rect 259503 337977 259515 337980
rect 259457 337971 259515 337977
rect 263594 337968 263600 337980
rect 263652 337968 263658 338020
rect 294049 338011 294107 338017
rect 294049 337977 294061 338011
rect 294095 338008 294107 338011
rect 335906 338008 335912 338020
rect 294095 337980 335912 338008
rect 294095 337977 294107 337980
rect 294049 337971 294107 337977
rect 335906 337968 335912 337980
rect 335964 337968 335970 338020
rect 336553 338011 336611 338017
rect 336553 337977 336565 338011
rect 336599 338008 336611 338011
rect 344462 338008 344468 338020
rect 336599 337980 344468 338008
rect 336599 337977 336611 337980
rect 336553 337971 336611 337977
rect 344462 337968 344468 337980
rect 344520 337968 344526 338020
rect 349062 337968 349068 338020
rect 349120 338008 349126 338020
rect 352837 338011 352895 338017
rect 352837 338008 352849 338011
rect 349120 337980 352849 338008
rect 349120 337968 349126 337980
rect 352837 337977 352849 337980
rect 352883 337977 352895 338011
rect 352944 338008 352972 338048
rect 353021 338045 353033 338079
rect 353067 338076 353079 338079
rect 357434 338076 357440 338088
rect 353067 338048 357440 338076
rect 353067 338045 353079 338048
rect 353021 338039 353079 338045
rect 357434 338036 357440 338048
rect 357492 338036 357498 338088
rect 363046 338036 363052 338088
rect 363104 338076 363110 338088
rect 363138 338076 363144 338088
rect 363104 338048 363144 338076
rect 363104 338036 363110 338048
rect 363138 338036 363144 338048
rect 363196 338036 363202 338088
rect 377674 338036 377680 338088
rect 377732 338076 377738 338088
rect 377732 338048 383424 338076
rect 377732 338036 377738 338048
rect 360194 338008 360200 338020
rect 352944 337980 360200 338008
rect 352837 337971 352895 337977
rect 360194 337968 360200 337980
rect 360252 337968 360258 338020
rect 376294 337968 376300 338020
rect 376352 338008 376358 338020
rect 381817 338011 381875 338017
rect 381817 338008 381829 338011
rect 376352 337980 381829 338008
rect 376352 337968 376358 337980
rect 381817 337977 381829 337980
rect 381863 337977 381875 338011
rect 381817 337971 381875 337977
rect 66898 337900 66904 337952
rect 66956 337940 66962 337952
rect 245654 337940 245660 337952
rect 66956 337912 245660 337940
rect 66956 337900 66962 337912
rect 245654 337900 245660 337912
rect 245712 337900 245718 337952
rect 251818 337900 251824 337952
rect 251876 337940 251882 337952
rect 256878 337940 256884 337952
rect 251876 337912 256884 337940
rect 251876 337900 251882 337912
rect 256878 337900 256884 337912
rect 256936 337900 256942 337952
rect 259546 337900 259552 337952
rect 259604 337940 259610 337952
rect 266354 337940 266360 337952
rect 259604 337912 266360 337940
rect 259604 337900 259610 337912
rect 266354 337900 266360 337912
rect 266412 337900 266418 337952
rect 297361 337943 297419 337949
rect 297361 337909 297373 337943
rect 297407 337940 297419 337943
rect 334526 337940 334532 337952
rect 297407 337912 334532 337940
rect 297407 337909 297419 337912
rect 297361 337903 297419 337909
rect 334526 337900 334532 337912
rect 334584 337900 334590 337952
rect 334710 337900 334716 337952
rect 334768 337940 334774 337952
rect 345382 337940 345388 337952
rect 334768 337912 345388 337940
rect 334768 337900 334774 337912
rect 345382 337900 345388 337912
rect 345440 337900 345446 337952
rect 345750 337900 345756 337952
rect 345808 337940 345814 337952
rect 351638 337940 351644 337952
rect 345808 337912 351644 337940
rect 345808 337900 345814 337912
rect 351638 337900 351644 337912
rect 351696 337900 351702 337952
rect 351822 337900 351828 337952
rect 351880 337940 351886 337952
rect 355137 337943 355195 337949
rect 355137 337940 355149 337943
rect 351880 337912 355149 337940
rect 351880 337900 351886 337912
rect 355137 337909 355149 337912
rect 355183 337909 355195 337943
rect 361022 337940 361028 337952
rect 355137 337903 355195 337909
rect 355244 337912 361028 337940
rect 61378 337832 61384 337884
rect 61436 337872 61442 337884
rect 246114 337872 246120 337884
rect 61436 337844 246120 337872
rect 61436 337832 61442 337844
rect 246114 337832 246120 337844
rect 246172 337832 246178 337884
rect 250438 337832 250444 337884
rect 250496 337872 250502 337884
rect 254210 337872 254216 337884
rect 250496 337844 254216 337872
rect 250496 337832 250502 337844
rect 254210 337832 254216 337844
rect 254268 337832 254274 337884
rect 259365 337875 259423 337881
rect 259365 337872 259377 337875
rect 254320 337844 259377 337872
rect 57238 337764 57244 337816
rect 57296 337804 57302 337816
rect 242986 337804 242992 337816
rect 57296 337776 242992 337804
rect 57296 337764 57302 337776
rect 242986 337764 242992 337776
rect 243044 337764 243050 337816
rect 253845 337807 253903 337813
rect 253845 337773 253857 337807
rect 253891 337804 253903 337807
rect 254320 337804 254348 337844
rect 259365 337841 259377 337844
rect 259411 337841 259423 337875
rect 259365 337835 259423 337841
rect 302145 337875 302203 337881
rect 302145 337841 302157 337875
rect 302191 337872 302203 337875
rect 339954 337872 339960 337884
rect 302191 337844 339960 337872
rect 302191 337841 302203 337844
rect 302145 337835 302203 337841
rect 339954 337832 339960 337844
rect 340012 337832 340018 337884
rect 341705 337875 341763 337881
rect 341705 337841 341717 337875
rect 341751 337872 341763 337875
rect 349430 337872 349436 337884
rect 341751 337844 349436 337872
rect 341751 337841 341763 337844
rect 341705 337835 341763 337841
rect 349430 337832 349436 337844
rect 349488 337832 349494 337884
rect 352006 337832 352012 337884
rect 352064 337872 352070 337884
rect 352742 337872 352748 337884
rect 352064 337844 352748 337872
rect 352064 337832 352070 337844
rect 352742 337832 352748 337844
rect 352800 337832 352806 337884
rect 352837 337875 352895 337881
rect 352837 337841 352849 337875
rect 352883 337872 352895 337875
rect 355244 337872 355272 337912
rect 361022 337900 361028 337912
rect 361080 337900 361086 337952
rect 379422 337900 379428 337952
rect 379480 337940 379486 337952
rect 383396 337940 383424 338048
rect 384850 338036 384856 338088
rect 384908 338076 384914 338088
rect 390557 338079 390615 338085
rect 390557 338076 390569 338079
rect 384908 338048 390569 338076
rect 384908 338036 384914 338048
rect 390557 338045 390569 338048
rect 390603 338045 390615 338079
rect 390557 338039 390615 338045
rect 418522 338036 418528 338088
rect 418580 338076 418586 338088
rect 426989 338079 427047 338085
rect 426989 338076 427001 338079
rect 418580 338048 427001 338076
rect 418580 338036 418586 338048
rect 426989 338045 427001 338048
rect 427035 338045 427047 338079
rect 427096 338076 427124 338116
rect 431034 338104 431040 338156
rect 431092 338144 431098 338156
rect 431092 338116 431356 338144
rect 431092 338104 431098 338116
rect 431218 338076 431224 338088
rect 427096 338048 431224 338076
rect 426989 338039 427047 338045
rect 431218 338036 431224 338048
rect 431276 338036 431282 338088
rect 431328 338076 431356 338116
rect 432340 338076 432368 338184
rect 433429 338181 433441 338184
rect 433475 338181 433487 338215
rect 433429 338175 433487 338181
rect 434070 338144 434076 338156
rect 432432 338116 434076 338144
rect 432432 338085 432460 338116
rect 434070 338104 434076 338116
rect 434128 338104 434134 338156
rect 431328 338048 432368 338076
rect 432417 338079 432475 338085
rect 432417 338045 432429 338079
rect 432463 338045 432475 338079
rect 432417 338039 432475 338045
rect 432509 338079 432567 338085
rect 432509 338045 432521 338079
rect 432555 338076 432567 338079
rect 502978 338076 502984 338088
rect 432555 338048 502984 338076
rect 432555 338045 432567 338048
rect 432509 338039 432567 338045
rect 502978 338036 502984 338048
rect 503036 338036 503042 338088
rect 383565 338011 383623 338017
rect 383565 337977 383577 338011
rect 383611 338008 383623 338011
rect 383611 337980 388484 338008
rect 383611 337977 383623 337980
rect 383565 337971 383623 337977
rect 388456 337940 388484 337980
rect 390278 337968 390284 338020
rect 390336 338008 390342 338020
rect 396905 338011 396963 338017
rect 396905 338008 396917 338011
rect 390336 337980 396917 338008
rect 390336 337968 390342 337980
rect 396905 337977 396917 337980
rect 396951 337977 396963 338011
rect 396905 337971 396963 337977
rect 396994 337968 397000 338020
rect 397052 338008 397058 338020
rect 406378 338008 406384 338020
rect 397052 337980 406384 338008
rect 397052 337968 397058 337980
rect 406378 337968 406384 337980
rect 406436 337968 406442 338020
rect 421190 337968 421196 338020
rect 421248 338008 421254 338020
rect 500218 338008 500224 338020
rect 421248 337980 500224 338008
rect 421248 337968 421254 337980
rect 500218 337968 500224 337980
rect 500276 337968 500282 338020
rect 393958 337940 393964 337952
rect 379480 337912 383240 337940
rect 383396 337912 386092 337940
rect 388456 337912 393964 337940
rect 379480 337900 379486 337912
rect 352883 337844 355272 337872
rect 352883 337841 352895 337844
rect 352837 337835 352895 337841
rect 355318 337832 355324 337884
rect 355376 337872 355382 337884
rect 359274 337872 359280 337884
rect 355376 337844 359280 337872
rect 355376 337832 355382 337844
rect 359274 337832 359280 337844
rect 359332 337832 359338 337884
rect 370038 337832 370044 337884
rect 370096 337872 370102 337884
rect 371050 337872 371056 337884
rect 370096 337844 371056 337872
rect 370096 337832 370102 337844
rect 371050 337832 371056 337844
rect 371108 337832 371114 337884
rect 380802 337832 380808 337884
rect 380860 337832 380866 337884
rect 383212 337872 383240 337912
rect 385957 337875 386015 337881
rect 385957 337872 385969 337875
rect 383212 337844 385969 337872
rect 385957 337841 385969 337844
rect 386003 337841 386015 337875
rect 386064 337872 386092 337912
rect 393958 337900 393964 337912
rect 394016 337900 394022 337952
rect 399478 337940 399484 337952
rect 395908 337912 399484 337940
rect 388438 337872 388444 337884
rect 386064 337844 388444 337872
rect 385957 337835 386015 337841
rect 388438 337832 388444 337844
rect 388496 337832 388502 337884
rect 388533 337875 388591 337881
rect 388533 337841 388545 337875
rect 388579 337872 388591 337875
rect 395338 337872 395344 337884
rect 388579 337844 395344 337872
rect 388579 337841 388591 337844
rect 388533 337835 388591 337841
rect 395338 337832 395344 337844
rect 395396 337832 395402 337884
rect 253891 337776 254348 337804
rect 253891 337773 253903 337776
rect 253845 337767 253903 337773
rect 254578 337764 254584 337816
rect 254636 337804 254642 337816
rect 259457 337807 259515 337813
rect 259457 337804 259469 337807
rect 254636 337776 259469 337804
rect 254636 337764 254642 337776
rect 259457 337773 259469 337776
rect 259503 337773 259515 337807
rect 260926 337804 260932 337816
rect 259457 337767 259515 337773
rect 259564 337776 260932 337804
rect 42058 337696 42064 337748
rect 42116 337736 42122 337748
rect 229833 337739 229891 337745
rect 229833 337736 229845 337739
rect 42116 337708 229845 337736
rect 42116 337696 42122 337708
rect 229833 337705 229845 337708
rect 229879 337705 229891 337739
rect 229833 337699 229891 337705
rect 229925 337739 229983 337745
rect 229925 337705 229937 337739
rect 229971 337736 229983 337739
rect 233970 337736 233976 337748
rect 229971 337708 233976 337736
rect 229971 337705 229983 337708
rect 229925 337699 229983 337705
rect 233970 337696 233976 337708
rect 234028 337696 234034 337748
rect 259365 337739 259423 337745
rect 259365 337705 259377 337739
rect 259411 337736 259423 337739
rect 259564 337736 259592 337776
rect 260926 337764 260932 337776
rect 260984 337764 260990 337816
rect 285582 337764 285588 337816
rect 285640 337804 285646 337816
rect 337286 337804 337292 337816
rect 285640 337776 337292 337804
rect 285640 337764 285646 337776
rect 337286 337764 337292 337776
rect 337344 337764 337350 337816
rect 337933 337807 337991 337813
rect 337933 337773 337945 337807
rect 337979 337804 337991 337807
rect 344002 337804 344008 337816
rect 337979 337776 344008 337804
rect 337979 337773 337991 337776
rect 337933 337767 337991 337773
rect 344002 337764 344008 337776
rect 344060 337764 344066 337816
rect 344922 337764 344928 337816
rect 344980 337804 344986 337816
rect 359734 337804 359740 337816
rect 344980 337776 359740 337804
rect 344980 337764 344986 337776
rect 359734 337764 359740 337776
rect 359792 337764 359798 337816
rect 374546 337764 374552 337816
rect 374604 337804 374610 337816
rect 376018 337804 376024 337816
rect 374604 337776 376024 337804
rect 374604 337764 374610 337776
rect 376018 337764 376024 337776
rect 376076 337764 376082 337816
rect 380820 337804 380848 337832
rect 380820 337776 382320 337804
rect 259411 337708 259592 337736
rect 259411 337705 259423 337708
rect 259365 337699 259423 337705
rect 276750 337696 276756 337748
rect 276808 337736 276814 337748
rect 329650 337736 329656 337748
rect 276808 337708 329656 337736
rect 276808 337696 276814 337708
rect 329650 337696 329656 337708
rect 329708 337696 329714 337748
rect 331122 337696 331128 337748
rect 331180 337736 331186 337748
rect 340049 337739 340107 337745
rect 340049 337736 340061 337739
rect 331180 337708 340061 337736
rect 331180 337696 331186 337708
rect 340049 337705 340061 337708
rect 340095 337705 340107 337739
rect 345661 337739 345719 337745
rect 345661 337736 345673 337739
rect 340049 337699 340107 337705
rect 340156 337708 345673 337736
rect 39298 337628 39304 337680
rect 39356 337668 39362 337680
rect 243446 337668 243452 337680
rect 39356 337640 243452 337668
rect 39356 337628 39362 337640
rect 243446 337628 243452 337640
rect 243504 337628 243510 337680
rect 254854 337628 254860 337680
rect 254912 337668 254918 337680
rect 259454 337668 259460 337680
rect 254912 337640 259460 337668
rect 254912 337628 254918 337640
rect 259454 337628 259460 337640
rect 259512 337628 259518 337680
rect 287701 337671 287759 337677
rect 287701 337637 287713 337671
rect 287747 337668 287759 337671
rect 326249 337671 326307 337677
rect 326249 337668 326261 337671
rect 287747 337640 326261 337668
rect 287747 337637 287759 337640
rect 287701 337631 287759 337637
rect 326249 337637 326261 337640
rect 326295 337637 326307 337671
rect 333698 337668 333704 337680
rect 326249 337631 326307 337637
rect 326356 337640 333704 337668
rect 35158 337560 35164 337612
rect 35216 337600 35222 337612
rect 240778 337600 240784 337612
rect 35216 337572 240784 337600
rect 35216 337560 35222 337572
rect 240778 337560 240784 337572
rect 240836 337560 240842 337612
rect 258810 337560 258816 337612
rect 258868 337600 258874 337612
rect 259549 337603 259607 337609
rect 259549 337600 259561 337603
rect 258868 337572 259561 337600
rect 258868 337560 258874 337572
rect 259549 337569 259561 337572
rect 259595 337569 259607 337603
rect 259549 337563 259607 337569
rect 259733 337603 259791 337609
rect 259733 337569 259745 337603
rect 259779 337600 259791 337603
rect 275738 337600 275744 337612
rect 259779 337572 275744 337600
rect 259779 337569 259791 337572
rect 259733 337563 259791 337569
rect 275738 337560 275744 337572
rect 275796 337560 275802 337612
rect 276658 337560 276664 337612
rect 276716 337600 276722 337612
rect 326356 337600 326384 337640
rect 333698 337628 333704 337640
rect 333756 337628 333762 337680
rect 276716 337572 326384 337600
rect 326433 337603 326491 337609
rect 276716 337560 276722 337572
rect 326433 337569 326445 337603
rect 326479 337600 326491 337603
rect 330386 337600 330392 337612
rect 326479 337572 330392 337600
rect 326479 337569 326491 337572
rect 326433 337563 326491 337569
rect 330386 337560 330392 337572
rect 330444 337560 330450 337612
rect 330478 337560 330484 337612
rect 330536 337600 330542 337612
rect 340156 337600 340184 337708
rect 345661 337705 345673 337708
rect 345707 337705 345719 337739
rect 345661 337699 345719 337705
rect 352558 337696 352564 337748
rect 352616 337736 352622 337748
rect 353386 337736 353392 337748
rect 352616 337708 353392 337736
rect 352616 337696 352622 337708
rect 353386 337696 353392 337708
rect 353444 337696 353450 337748
rect 353481 337739 353539 337745
rect 353481 337705 353493 337739
rect 353527 337736 353539 337739
rect 356609 337739 356667 337745
rect 356609 337736 356621 337739
rect 353527 337708 356621 337736
rect 353527 337705 353539 337708
rect 353481 337699 353539 337705
rect 356609 337705 356621 337708
rect 356655 337705 356667 337739
rect 356609 337699 356667 337705
rect 356698 337696 356704 337748
rect 356756 337736 356762 337748
rect 360562 337736 360568 337748
rect 356756 337708 360568 337736
rect 356756 337696 356762 337708
rect 360562 337696 360568 337708
rect 360620 337696 360626 337748
rect 372246 337696 372252 337748
rect 372304 337736 372310 337748
rect 373258 337736 373264 337748
rect 372304 337708 373264 337736
rect 372304 337696 372310 337708
rect 373258 337696 373264 337708
rect 373316 337696 373322 337748
rect 374086 337696 374092 337748
rect 374144 337736 374150 337748
rect 375282 337736 375288 337748
rect 374144 337708 375288 337736
rect 374144 337696 374150 337708
rect 375282 337696 375288 337708
rect 375340 337696 375346 337748
rect 377214 337696 377220 337748
rect 377272 337736 377278 337748
rect 377950 337736 377956 337748
rect 377272 337708 377956 337736
rect 377272 337696 377278 337708
rect 377950 337696 377956 337708
rect 378008 337696 378014 337748
rect 379882 337696 379888 337748
rect 379940 337736 379946 337748
rect 380802 337736 380808 337748
rect 379940 337708 380808 337736
rect 379940 337696 379946 337708
rect 380802 337696 380808 337708
rect 380860 337696 380866 337748
rect 381262 337696 381268 337748
rect 381320 337736 381326 337748
rect 382182 337736 382188 337748
rect 381320 337708 382188 337736
rect 381320 337696 381326 337708
rect 382182 337696 382188 337708
rect 382240 337696 382246 337748
rect 382292 337736 382320 337776
rect 382642 337764 382648 337816
rect 382700 337804 382706 337816
rect 383565 337807 383623 337813
rect 383565 337804 383577 337807
rect 382700 337776 383577 337804
rect 382700 337764 382706 337776
rect 383565 337773 383577 337776
rect 383611 337773 383623 337807
rect 383565 337767 383623 337773
rect 393866 337764 393872 337816
rect 393924 337804 393930 337816
rect 394418 337804 394424 337816
rect 393924 337776 394424 337804
rect 393924 337764 393930 337776
rect 394418 337764 394424 337776
rect 394476 337764 394482 337816
rect 383841 337739 383899 337745
rect 383841 337736 383853 337739
rect 382292 337708 383853 337736
rect 383841 337705 383853 337708
rect 383887 337705 383899 337739
rect 383841 337699 383899 337705
rect 383930 337696 383936 337748
rect 383988 337736 383994 337748
rect 384942 337736 384948 337748
rect 383988 337708 384948 337736
rect 383988 337696 383994 337708
rect 384942 337696 384948 337708
rect 385000 337696 385006 337748
rect 389358 337696 389364 337748
rect 389416 337736 389422 337748
rect 390462 337736 390468 337748
rect 389416 337708 390468 337736
rect 389416 337696 389422 337708
rect 390462 337696 390468 337708
rect 390520 337696 390526 337748
rect 390557 337739 390615 337745
rect 390557 337705 390569 337739
rect 390603 337736 390615 337739
rect 395908 337736 395936 337912
rect 399478 337900 399484 337912
rect 399536 337900 399542 337952
rect 406746 337900 406752 337952
rect 406804 337940 406810 337952
rect 406804 337912 415072 337940
rect 406804 337900 406810 337912
rect 398282 337832 398288 337884
rect 398340 337872 398346 337884
rect 409138 337872 409144 337884
rect 398340 337844 409144 337872
rect 398340 337832 398346 337844
rect 409138 337832 409144 337844
rect 409196 337832 409202 337884
rect 415044 337872 415072 337912
rect 415854 337900 415860 337952
rect 415912 337940 415918 337952
rect 427081 337943 427139 337949
rect 427081 337940 427093 337943
rect 415912 337912 427093 337940
rect 415912 337900 415918 337912
rect 427081 337909 427093 337912
rect 427127 337909 427139 337943
rect 427081 337903 427139 337909
rect 427170 337900 427176 337952
rect 427228 337940 427234 337952
rect 428458 337940 428464 337952
rect 427228 337912 428464 337940
rect 427228 337900 427234 337912
rect 428458 337900 428464 337912
rect 428516 337900 428522 337952
rect 429102 337900 429108 337952
rect 429160 337940 429166 337952
rect 432417 337943 432475 337949
rect 432417 337940 432429 337943
rect 429160 337912 432429 337940
rect 429160 337900 429166 337912
rect 432417 337909 432429 337912
rect 432463 337909 432475 337943
rect 507118 337940 507124 337952
rect 432417 337903 432475 337909
rect 432616 337912 507124 337940
rect 417418 337872 417424 337884
rect 415044 337844 417424 337872
rect 417418 337832 417424 337844
rect 417476 337832 417482 337884
rect 423858 337832 423864 337884
rect 423916 337872 423922 337884
rect 432509 337875 432567 337881
rect 432509 337872 432521 337875
rect 423916 337844 432521 337872
rect 423916 337832 423922 337844
rect 432509 337841 432521 337844
rect 432555 337841 432567 337875
rect 432509 337835 432567 337841
rect 399110 337804 399116 337816
rect 390603 337708 395936 337736
rect 396000 337776 399116 337804
rect 390603 337705 390615 337708
rect 390557 337699 390615 337705
rect 340782 337628 340788 337680
rect 340840 337668 340846 337680
rect 358354 337668 358360 337680
rect 340840 337640 358360 337668
rect 340840 337628 340846 337640
rect 358354 337628 358360 337640
rect 358412 337628 358418 337680
rect 372706 337628 372712 337680
rect 372764 337668 372770 337680
rect 373902 337668 373908 337680
rect 372764 337640 373908 337668
rect 372764 337628 372770 337640
rect 373902 337628 373908 337640
rect 373960 337628 373966 337680
rect 375834 337628 375840 337680
rect 375892 337668 375898 337680
rect 377398 337668 377404 337680
rect 375892 337640 377404 337668
rect 375892 337628 375898 337640
rect 377398 337628 377404 337640
rect 377456 337628 377462 337680
rect 378594 337628 378600 337680
rect 378652 337668 378658 337680
rect 380158 337668 380164 337680
rect 378652 337640 380164 337668
rect 378652 337628 378658 337640
rect 380158 337628 380164 337640
rect 380216 337628 380222 337680
rect 380342 337628 380348 337680
rect 380400 337668 380406 337680
rect 396000 337668 396028 337776
rect 399110 337764 399116 337776
rect 399168 337764 399174 337816
rect 403710 337764 403716 337816
rect 403768 337804 403774 337816
rect 411898 337804 411904 337816
rect 403768 337776 411904 337804
rect 403768 337764 403774 337776
rect 411898 337764 411904 337776
rect 411956 337764 411962 337816
rect 420178 337804 420184 337816
rect 413940 337776 420184 337804
rect 396534 337696 396540 337748
rect 396592 337736 396598 337748
rect 397270 337736 397276 337748
rect 396592 337708 397276 337736
rect 396592 337696 396598 337708
rect 397270 337696 397276 337708
rect 397328 337696 397334 337748
rect 397822 337696 397828 337748
rect 397880 337736 397886 337748
rect 398558 337736 398564 337748
rect 397880 337708 398564 337736
rect 397880 337696 397886 337708
rect 398558 337696 398564 337708
rect 398616 337696 398622 337748
rect 399202 337696 399208 337748
rect 399260 337736 399266 337748
rect 400030 337736 400036 337748
rect 399260 337708 400036 337736
rect 399260 337696 399266 337708
rect 400030 337696 400036 337708
rect 400088 337696 400094 337748
rect 400582 337696 400588 337748
rect 400640 337736 400646 337748
rect 401410 337736 401416 337748
rect 400640 337708 401416 337736
rect 400640 337696 400646 337708
rect 401410 337696 401416 337708
rect 401468 337696 401474 337748
rect 401870 337696 401876 337748
rect 401928 337736 401934 337748
rect 402790 337736 402796 337748
rect 401928 337708 402796 337736
rect 401928 337696 401934 337708
rect 402790 337696 402796 337708
rect 402848 337696 402854 337748
rect 403250 337696 403256 337748
rect 403308 337736 403314 337748
rect 404170 337736 404176 337748
rect 403308 337708 404176 337736
rect 403308 337696 403314 337708
rect 404170 337696 404176 337708
rect 404228 337696 404234 337748
rect 404630 337696 404636 337748
rect 404688 337736 404694 337748
rect 405550 337736 405556 337748
rect 404688 337708 405556 337736
rect 404688 337696 404694 337708
rect 405550 337696 405556 337708
rect 405608 337696 405614 337748
rect 405918 337696 405924 337748
rect 405976 337736 405982 337748
rect 406930 337736 406936 337748
rect 405976 337708 406936 337736
rect 405976 337696 405982 337708
rect 406930 337696 406936 337708
rect 406988 337696 406994 337748
rect 407298 337696 407304 337748
rect 407356 337736 407362 337748
rect 408310 337736 408316 337748
rect 407356 337708 408316 337736
rect 407356 337696 407362 337708
rect 408310 337696 408316 337708
rect 408368 337696 408374 337748
rect 409046 337696 409052 337748
rect 409104 337736 409110 337748
rect 413940 337736 413968 337776
rect 420178 337764 420184 337776
rect 420236 337764 420242 337816
rect 422570 337764 422576 337816
rect 422628 337804 422634 337816
rect 422628 337776 426572 337804
rect 422628 337764 422634 337776
rect 409104 337708 413968 337736
rect 409104 337696 409110 337708
rect 414014 337696 414020 337748
rect 414072 337736 414078 337748
rect 415302 337736 415308 337748
rect 414072 337708 415308 337736
rect 414072 337696 414078 337708
rect 415302 337696 415308 337708
rect 415360 337696 415366 337748
rect 423030 337696 423036 337748
rect 423088 337736 423094 337748
rect 423582 337736 423588 337748
rect 423088 337708 423588 337736
rect 423088 337696 423094 337708
rect 423582 337696 423588 337708
rect 423640 337696 423646 337748
rect 424318 337696 424324 337748
rect 424376 337736 424382 337748
rect 424962 337736 424968 337748
rect 424376 337708 424968 337736
rect 424376 337696 424382 337708
rect 424962 337696 424968 337708
rect 425020 337696 425026 337748
rect 425609 337739 425667 337745
rect 425609 337736 425621 337739
rect 425164 337708 425621 337736
rect 380400 337640 396028 337668
rect 380400 337628 380406 337640
rect 396074 337628 396080 337680
rect 396132 337668 396138 337680
rect 397362 337668 397368 337680
rect 396132 337640 397368 337668
rect 396132 337628 396138 337640
rect 397362 337628 397368 337640
rect 397420 337628 397426 337680
rect 397454 337628 397460 337680
rect 397512 337668 397518 337680
rect 398650 337668 398656 337680
rect 397512 337640 398656 337668
rect 397512 337628 397518 337640
rect 398650 337628 398656 337640
rect 398708 337628 398714 337680
rect 401042 337628 401048 337680
rect 401100 337668 401106 337680
rect 410518 337668 410524 337680
rect 401100 337640 410524 337668
rect 401100 337628 401106 337640
rect 410518 337628 410524 337640
rect 410576 337628 410582 337680
rect 412634 337628 412640 337680
rect 412692 337668 412698 337680
rect 413922 337668 413928 337680
rect 412692 337640 413928 337668
rect 412692 337628 412698 337640
rect 413922 337628 413928 337640
rect 413980 337628 413986 337680
rect 414474 337628 414480 337680
rect 414532 337668 414538 337680
rect 417053 337671 417111 337677
rect 417053 337668 417065 337671
rect 414532 337640 417065 337668
rect 414532 337628 414538 337640
rect 417053 337637 417065 337640
rect 417099 337637 417111 337671
rect 417053 337631 417111 337637
rect 417142 337628 417148 337680
rect 417200 337668 417206 337680
rect 425164 337668 425192 337708
rect 425609 337705 425621 337708
rect 425655 337705 425667 337739
rect 425609 337699 425667 337705
rect 425698 337696 425704 337748
rect 425756 337736 425762 337748
rect 426342 337736 426348 337748
rect 425756 337708 426348 337736
rect 425756 337696 425762 337708
rect 426342 337696 426348 337708
rect 426400 337696 426406 337748
rect 426544 337736 426572 337776
rect 426618 337764 426624 337816
rect 426676 337804 426682 337816
rect 432616 337804 432644 337912
rect 507118 337900 507124 337912
rect 507176 337900 507182 337952
rect 432693 337875 432751 337881
rect 432693 337841 432705 337875
rect 432739 337872 432751 337875
rect 437293 337875 437351 337881
rect 437293 337872 437305 337875
rect 432739 337844 437305 337872
rect 432739 337841 432751 337844
rect 432693 337835 432751 337841
rect 437293 337841 437305 337844
rect 437339 337841 437351 337875
rect 437293 337835 437351 337841
rect 437382 337832 437388 337884
rect 437440 337872 437446 337884
rect 442169 337875 442227 337881
rect 442169 337872 442181 337875
rect 437440 337844 442181 337872
rect 437440 337832 437446 337844
rect 442169 337841 442181 337844
rect 442215 337841 442227 337875
rect 442169 337835 442227 337841
rect 442261 337875 442319 337881
rect 442261 337841 442273 337875
rect 442307 337872 442319 337875
rect 514018 337872 514024 337884
rect 442307 337844 514024 337872
rect 442307 337841 442319 337844
rect 442261 337835 442319 337841
rect 514018 337832 514024 337844
rect 514076 337832 514082 337884
rect 426676 337776 432644 337804
rect 433337 337807 433395 337813
rect 426676 337764 426682 337776
rect 433337 337773 433349 337807
rect 433383 337804 433395 337807
rect 511258 337804 511264 337816
rect 433383 337776 511264 337804
rect 433383 337773 433395 337776
rect 433337 337767 433395 337773
rect 511258 337764 511264 337776
rect 511316 337764 511322 337816
rect 426986 337736 426992 337748
rect 426544 337708 426992 337736
rect 426986 337696 426992 337708
rect 427044 337696 427050 337748
rect 427078 337696 427084 337748
rect 427136 337736 427142 337748
rect 427722 337736 427728 337748
rect 427136 337708 427728 337736
rect 427136 337696 427142 337708
rect 427722 337696 427728 337708
rect 427780 337696 427786 337748
rect 427906 337696 427912 337748
rect 427964 337736 427970 337748
rect 429102 337736 429108 337748
rect 427964 337708 429108 337736
rect 427964 337696 427970 337708
rect 429102 337696 429108 337708
rect 429160 337696 429166 337748
rect 429286 337696 429292 337748
rect 429344 337736 429350 337748
rect 429344 337708 431908 337736
rect 429344 337696 429350 337708
rect 417200 337640 425192 337668
rect 417200 337628 417206 337640
rect 425238 337628 425244 337680
rect 425296 337668 425302 337680
rect 429838 337668 429844 337680
rect 425296 337640 429844 337668
rect 425296 337628 425302 337640
rect 429838 337628 429844 337640
rect 429896 337628 429902 337680
rect 431880 337668 431908 337708
rect 431954 337696 431960 337748
rect 432012 337736 432018 337748
rect 437017 337739 437075 337745
rect 437017 337736 437029 337739
rect 432012 337708 437029 337736
rect 432012 337696 432018 337708
rect 437017 337705 437029 337708
rect 437063 337705 437075 337739
rect 437017 337699 437075 337705
rect 438762 337696 438768 337748
rect 438820 337736 438826 337748
rect 442905 337739 442963 337745
rect 442905 337736 442917 337739
rect 438820 337708 442917 337736
rect 438820 337696 438826 337708
rect 442905 337705 442917 337708
rect 442951 337705 442963 337739
rect 442905 337699 442963 337705
rect 444098 337696 444104 337748
rect 444156 337736 444162 337748
rect 446953 337739 447011 337745
rect 446953 337736 446965 337739
rect 444156 337708 446965 337736
rect 444156 337696 444162 337708
rect 446953 337705 446965 337708
rect 446999 337705 447011 337739
rect 518158 337736 518164 337748
rect 446953 337699 447011 337705
rect 447152 337708 518164 337736
rect 433337 337671 433395 337677
rect 433337 337668 433349 337671
rect 431880 337640 433349 337668
rect 433337 337637 433349 337640
rect 433383 337637 433395 337671
rect 433337 337631 433395 337637
rect 433429 337671 433487 337677
rect 433429 337637 433441 337671
rect 433475 337668 433487 337671
rect 436370 337668 436376 337680
rect 433475 337640 436376 337668
rect 433475 337637 433487 337640
rect 433429 337631 433487 337637
rect 436370 337628 436376 337640
rect 436428 337628 436434 337680
rect 436462 337628 436468 337680
rect 436520 337668 436526 337680
rect 437382 337668 437388 337680
rect 436520 337640 437388 337668
rect 436520 337628 436526 337640
rect 437382 337628 437388 337640
rect 437440 337628 437446 337680
rect 441430 337628 441436 337680
rect 441488 337668 441494 337680
rect 444834 337668 444840 337680
rect 441488 337640 444840 337668
rect 441488 337628 441494 337640
rect 444834 337628 444840 337640
rect 444892 337628 444898 337680
rect 444929 337671 444987 337677
rect 444929 337637 444941 337671
rect 444975 337668 444987 337671
rect 445665 337671 445723 337677
rect 445665 337668 445677 337671
rect 444975 337640 445677 337668
rect 444975 337637 444987 337640
rect 444929 337631 444987 337637
rect 445665 337637 445677 337640
rect 445711 337637 445723 337671
rect 445665 337631 445723 337637
rect 445938 337628 445944 337680
rect 445996 337668 446002 337680
rect 447042 337668 447048 337680
rect 445996 337640 447048 337668
rect 445996 337628 446002 337640
rect 447042 337628 447048 337640
rect 447100 337628 447106 337680
rect 330536 337572 340184 337600
rect 340233 337603 340291 337609
rect 330536 337560 330542 337572
rect 340233 337569 340245 337603
rect 340279 337600 340291 337603
rect 356974 337600 356980 337612
rect 340279 337572 356980 337600
rect 340279 337569 340291 337572
rect 340233 337563 340291 337569
rect 356974 337560 356980 337572
rect 357032 337560 357038 337612
rect 358078 337560 358084 337612
rect 358136 337600 358142 337612
rect 363322 337600 363328 337612
rect 358136 337572 363328 337600
rect 358136 337560 358142 337572
rect 363322 337560 363328 337572
rect 363380 337560 363386 337612
rect 375374 337560 375380 337612
rect 375432 337600 375438 337612
rect 376662 337600 376668 337612
rect 375432 337572 376668 337600
rect 375432 337560 375438 337572
rect 376662 337560 376668 337572
rect 376720 337560 376726 337612
rect 379054 337560 379060 337612
rect 379112 337600 379118 337612
rect 381630 337600 381636 337612
rect 379112 337572 381636 337600
rect 379112 337560 379118 337572
rect 381630 337560 381636 337572
rect 381688 337560 381694 337612
rect 381740 337572 385172 337600
rect 28258 337492 28264 337544
rect 28316 337532 28322 337544
rect 229833 337535 229891 337541
rect 28316 337504 229784 337532
rect 28316 337492 28322 337504
rect 19978 337424 19984 337476
rect 20036 337464 20042 337476
rect 229649 337467 229707 337473
rect 229649 337464 229661 337467
rect 20036 337436 229661 337464
rect 20036 337424 20042 337436
rect 229649 337433 229661 337436
rect 229695 337433 229707 337467
rect 229756 337464 229784 337504
rect 229833 337501 229845 337535
rect 229879 337532 229891 337535
rect 237558 337532 237564 337544
rect 229879 337504 237564 337532
rect 229879 337501 229891 337504
rect 229833 337495 229891 337501
rect 237558 337492 237564 337504
rect 237616 337492 237622 337544
rect 258718 337492 258724 337544
rect 258776 337532 258782 337544
rect 273070 337532 273076 337544
rect 258776 337504 273076 337532
rect 258776 337492 258782 337504
rect 273070 337492 273076 337504
rect 273128 337492 273134 337544
rect 274542 337492 274548 337544
rect 274600 337532 274606 337544
rect 333238 337532 333244 337544
rect 274600 337504 333244 337532
rect 274600 337492 274606 337504
rect 333238 337492 333244 337504
rect 333296 337492 333302 337544
rect 334618 337492 334624 337544
rect 334676 337532 334682 337544
rect 345569 337535 345627 337541
rect 345569 337532 345581 337535
rect 334676 337504 345581 337532
rect 334676 337492 334682 337504
rect 345569 337501 345581 337504
rect 345615 337501 345627 337535
rect 345569 337495 345627 337501
rect 348418 337492 348424 337544
rect 348476 337532 348482 337544
rect 353021 337535 353079 337541
rect 353021 337532 353033 337535
rect 348476 337504 353033 337532
rect 348476 337492 348482 337504
rect 353021 337501 353033 337504
rect 353067 337501 353079 337535
rect 353021 337495 353079 337501
rect 353202 337492 353208 337544
rect 353260 337532 353266 337544
rect 353481 337535 353539 337541
rect 353481 337532 353493 337535
rect 353260 337504 353493 337532
rect 353260 337492 353266 337504
rect 353481 337501 353493 337504
rect 353527 337501 353539 337535
rect 353481 337495 353539 337501
rect 355137 337535 355195 337541
rect 355137 337501 355149 337535
rect 355183 337532 355195 337535
rect 362402 337532 362408 337544
rect 355183 337504 362408 337532
rect 355183 337501 355195 337504
rect 355137 337495 355195 337501
rect 362402 337492 362408 337504
rect 362460 337492 362466 337544
rect 371418 337492 371424 337544
rect 371476 337532 371482 337544
rect 374086 337532 374092 337544
rect 371476 337504 374092 337532
rect 371476 337492 371482 337504
rect 374086 337492 374092 337504
rect 374144 337492 374150 337544
rect 378134 337492 378140 337544
rect 378192 337532 378198 337544
rect 381740 337532 381768 337572
rect 378192 337504 381768 337532
rect 381817 337535 381875 337541
rect 378192 337492 378198 337504
rect 381817 337501 381829 337535
rect 381863 337532 381875 337535
rect 384298 337532 384304 337544
rect 381863 337504 384304 337532
rect 381863 337501 381875 337504
rect 381817 337495 381875 337501
rect 384298 337492 384304 337504
rect 384356 337492 384362 337544
rect 385144 337532 385172 337572
rect 386598 337560 386604 337612
rect 386656 337600 386662 337612
rect 387518 337600 387524 337612
rect 386656 337572 387524 337600
rect 386656 337560 386662 337572
rect 387518 337560 387524 337572
rect 387576 337560 387582 337612
rect 390646 337560 390652 337612
rect 390704 337600 390710 337612
rect 391658 337600 391664 337612
rect 390704 337572 391664 337600
rect 390704 337560 390710 337572
rect 391658 337560 391664 337572
rect 391716 337560 391722 337612
rect 392026 337560 392032 337612
rect 392084 337600 392090 337612
rect 393038 337600 393044 337612
rect 392084 337572 393044 337600
rect 392084 337560 392090 337572
rect 393038 337560 393044 337572
rect 393096 337560 393102 337612
rect 407758 337600 407764 337612
rect 393148 337572 407764 337600
rect 387058 337532 387064 337544
rect 385144 337504 387064 337532
rect 387058 337492 387064 337504
rect 387116 337492 387122 337544
rect 387978 337492 387984 337544
rect 388036 337532 388042 337544
rect 393148 337532 393176 337572
rect 407758 337560 407764 337572
rect 407816 337560 407822 337612
rect 408678 337560 408684 337612
rect 408736 337600 408742 337612
rect 435269 337603 435327 337609
rect 435269 337600 435281 337603
rect 408736 337572 435281 337600
rect 408736 337560 408742 337572
rect 435269 337569 435281 337572
rect 435315 337569 435327 337603
rect 435269 337563 435327 337569
rect 438210 337560 438216 337612
rect 438268 337600 438274 337612
rect 447152 337600 447180 337708
rect 518158 337696 518164 337708
rect 518216 337696 518222 337748
rect 447226 337628 447232 337680
rect 447284 337668 447290 337680
rect 448422 337668 448428 337680
rect 447284 337640 448428 337668
rect 447284 337628 447290 337640
rect 448422 337628 448428 337640
rect 448480 337628 448486 337680
rect 448606 337628 448612 337680
rect 448664 337668 448670 337680
rect 449802 337668 449808 337680
rect 448664 337640 449808 337668
rect 448664 337628 448670 337640
rect 449802 337628 449808 337640
rect 449860 337628 449866 337680
rect 529198 337668 529204 337680
rect 449912 337640 529204 337668
rect 438268 337572 447180 337600
rect 438268 337560 438274 337572
rect 447318 337560 447324 337612
rect 447376 337600 447382 337612
rect 449912 337600 449940 337640
rect 529198 337628 529204 337640
rect 529256 337628 529262 337680
rect 447376 337572 449940 337600
rect 449989 337603 450047 337609
rect 447376 337560 447382 337572
rect 449989 337569 450001 337603
rect 450035 337600 450047 337603
rect 527818 337600 527824 337612
rect 450035 337572 527824 337600
rect 450035 337569 450047 337572
rect 449989 337563 450047 337569
rect 527818 337560 527824 337572
rect 527876 337560 527882 337612
rect 388036 337504 393176 337532
rect 393225 337535 393283 337541
rect 388036 337492 388042 337504
rect 393225 337501 393237 337535
rect 393271 337532 393283 337535
rect 405090 337532 405096 337544
rect 393271 337504 405096 337532
rect 393271 337501 393283 337504
rect 393225 337495 393283 337501
rect 405090 337492 405096 337504
rect 405148 337492 405154 337544
rect 411806 337492 411812 337544
rect 411864 337532 411870 337544
rect 428277 337535 428335 337541
rect 411864 337504 428228 337532
rect 411864 337492 411870 337504
rect 237190 337464 237196 337476
rect 229756 337436 237196 337464
rect 229649 337427 229707 337433
rect 237190 337424 237196 337436
rect 237248 337424 237254 337476
rect 253845 337467 253903 337473
rect 253845 337464 253857 337467
rect 240428 337436 253857 337464
rect 13078 337356 13084 337408
rect 13136 337396 13142 337408
rect 233602 337396 233608 337408
rect 13136 337368 233608 337396
rect 13136 337356 13142 337368
rect 233602 337356 233608 337368
rect 233660 337356 233666 337408
rect 234154 337356 234160 337408
rect 234212 337396 234218 337408
rect 240318 337396 240324 337408
rect 234212 337368 240324 337396
rect 234212 337356 234218 337368
rect 240318 337356 240324 337368
rect 240376 337356 240382 337408
rect 89625 337331 89683 337337
rect 89625 337297 89637 337331
rect 89671 337328 89683 337331
rect 99377 337331 99435 337337
rect 99377 337328 99389 337331
rect 89671 337300 99389 337328
rect 89671 337297 89683 337300
rect 89625 337291 89683 337297
rect 99377 337297 99389 337300
rect 99423 337297 99435 337331
rect 99377 337291 99435 337297
rect 108945 337331 109003 337337
rect 108945 337297 108957 337331
rect 108991 337328 109003 337331
rect 118697 337331 118755 337337
rect 118697 337328 118709 337331
rect 108991 337300 118709 337328
rect 108991 337297 109003 337300
rect 108945 337291 109003 337297
rect 118697 337297 118709 337300
rect 118743 337297 118755 337331
rect 118697 337291 118755 337297
rect 128265 337331 128323 337337
rect 128265 337297 128277 337331
rect 128311 337328 128323 337331
rect 138014 337328 138020 337340
rect 128311 337300 138020 337328
rect 128311 337297 128323 337300
rect 128265 337291 128323 337297
rect 138014 337288 138020 337300
rect 138072 337288 138078 337340
rect 147582 337288 147588 337340
rect 147640 337328 147646 337340
rect 157334 337328 157340 337340
rect 147640 337300 157340 337328
rect 147640 337288 147646 337300
rect 157334 337288 157340 337300
rect 157392 337288 157398 337340
rect 166902 337288 166908 337340
rect 166960 337328 166966 337340
rect 176654 337328 176660 337340
rect 166960 337300 176660 337328
rect 166960 337288 166966 337300
rect 176654 337288 176660 337300
rect 176712 337288 176718 337340
rect 186222 337288 186228 337340
rect 186280 337328 186286 337340
rect 195974 337328 195980 337340
rect 186280 337300 195980 337328
rect 186280 337288 186286 337300
rect 195974 337288 195980 337300
rect 196032 337288 196038 337340
rect 205542 337288 205548 337340
rect 205600 337328 205606 337340
rect 215294 337328 215300 337340
rect 205600 337300 215300 337328
rect 205600 337288 205606 337300
rect 215294 337288 215300 337300
rect 215352 337288 215358 337340
rect 224862 337288 224868 337340
rect 224920 337328 224926 337340
rect 240428 337328 240456 337436
rect 253845 337433 253857 337436
rect 253891 337433 253903 337467
rect 253845 337427 253903 337433
rect 257338 337424 257344 337476
rect 257396 337464 257402 337476
rect 271690 337464 271696 337476
rect 257396 337436 271696 337464
rect 257396 337424 257402 337436
rect 271690 337424 271696 337436
rect 271748 337424 271754 337476
rect 271782 337424 271788 337476
rect 271840 337464 271846 337476
rect 331858 337464 331864 337476
rect 271840 337436 331864 337464
rect 271840 337424 271846 337436
rect 331858 337424 331864 337436
rect 331916 337424 331922 337476
rect 333882 337424 333888 337476
rect 333940 337464 333946 337476
rect 355686 337464 355692 337476
rect 333940 337436 355692 337464
rect 333940 337424 333946 337436
rect 355686 337424 355692 337436
rect 355744 337424 355750 337476
rect 356609 337467 356667 337473
rect 356609 337433 356621 337467
rect 356655 337464 356667 337467
rect 362862 337464 362868 337476
rect 356655 337436 362868 337464
rect 356655 337433 356667 337436
rect 356609 337427 356667 337433
rect 362862 337424 362868 337436
rect 362920 337424 362926 337476
rect 373166 337424 373172 337476
rect 373224 337464 373230 337476
rect 373224 337436 376524 337464
rect 373224 337424 373230 337436
rect 252830 337396 252836 337408
rect 224920 337300 240456 337328
rect 246132 337368 252836 337396
rect 224920 337288 224926 337300
rect 77938 337220 77944 337272
rect 77996 337260 78002 337272
rect 246132 337260 246160 337368
rect 252830 337356 252836 337368
rect 252888 337356 252894 337408
rect 268654 337396 268660 337408
rect 261036 337368 268660 337396
rect 255958 337288 255964 337340
rect 256016 337328 256022 337340
rect 261036 337328 261064 337368
rect 268654 337356 268660 337368
rect 268712 337356 268718 337408
rect 269022 337356 269028 337408
rect 269080 337396 269086 337408
rect 326157 337399 326215 337405
rect 326157 337396 326169 337399
rect 269080 337368 326169 337396
rect 269080 337356 269086 337368
rect 326157 337365 326169 337368
rect 326203 337365 326215 337399
rect 326157 337359 326215 337365
rect 326249 337399 326307 337405
rect 326249 337365 326261 337399
rect 326295 337396 326307 337399
rect 334526 337396 334532 337408
rect 326295 337368 334532 337396
rect 326295 337365 326307 337368
rect 326249 337359 326307 337365
rect 334526 337356 334532 337368
rect 334584 337356 334590 337408
rect 334802 337356 334808 337408
rect 334860 337396 334866 337408
rect 336366 337396 336372 337408
rect 334860 337368 336372 337396
rect 334860 337356 334866 337368
rect 336366 337356 336372 337368
rect 336424 337356 336430 337408
rect 340049 337399 340107 337405
rect 340049 337365 340061 337399
rect 340095 337396 340107 337399
rect 345477 337399 345535 337405
rect 345477 337396 345489 337399
rect 340095 337368 345489 337396
rect 340095 337365 340107 337368
rect 340049 337359 340107 337365
rect 345477 337365 345489 337368
rect 345523 337365 345535 337399
rect 345477 337359 345535 337365
rect 345661 337399 345719 337405
rect 345661 337365 345673 337399
rect 345707 337396 345719 337399
rect 352190 337396 352196 337408
rect 345707 337368 352196 337396
rect 345707 337365 345719 337368
rect 345661 337359 345719 337365
rect 352190 337356 352196 337368
rect 352248 337356 352254 337408
rect 355962 337356 355968 337408
rect 356020 337396 356026 337408
rect 363782 337396 363788 337408
rect 356020 337368 363788 337396
rect 356020 337356 356026 337368
rect 363782 337356 363788 337368
rect 363840 337356 363846 337408
rect 376496 337396 376524 337436
rect 376754 337424 376760 337476
rect 376812 337464 376818 337476
rect 378042 337464 378048 337476
rect 376812 337436 378048 337464
rect 376812 337424 376818 337436
rect 378042 337424 378048 337436
rect 378100 337424 378106 337476
rect 381722 337424 381728 337476
rect 381780 337464 381786 337476
rect 381780 337436 394648 337464
rect 381780 337424 381786 337436
rect 379606 337396 379612 337408
rect 376496 337368 379612 337396
rect 379606 337356 379612 337368
rect 379664 337356 379670 337408
rect 383010 337356 383016 337408
rect 383068 337396 383074 337408
rect 394513 337399 394571 337405
rect 394513 337396 394525 337399
rect 383068 337368 394525 337396
rect 383068 337356 383074 337368
rect 394513 337365 394525 337368
rect 394559 337365 394571 337399
rect 394513 337359 394571 337365
rect 256016 337300 261064 337328
rect 256016 337288 256022 337300
rect 279970 337288 279976 337340
rect 280028 337328 280034 337340
rect 287701 337331 287759 337337
rect 287701 337328 287713 337331
rect 280028 337300 287713 337328
rect 280028 337288 280034 337300
rect 287701 337297 287713 337300
rect 287747 337297 287759 337331
rect 287701 337291 287759 337297
rect 288066 337288 288072 337340
rect 288124 337328 288130 337340
rect 297361 337331 297419 337337
rect 297361 337328 297373 337331
rect 288124 337300 297373 337328
rect 288124 337288 288130 337300
rect 297361 337297 297373 337300
rect 297407 337297 297419 337331
rect 297361 337291 297419 337297
rect 303522 337288 303528 337340
rect 303580 337328 303586 337340
rect 337933 337331 337991 337337
rect 337933 337328 337945 337331
rect 303580 337300 337945 337328
rect 303580 337288 303586 337300
rect 337933 337297 337945 337300
rect 337979 337297 337991 337331
rect 337933 337291 337991 337297
rect 338022 337288 338028 337340
rect 338080 337328 338086 337340
rect 340233 337331 340291 337337
rect 340233 337328 340245 337331
rect 338080 337300 340245 337328
rect 338080 337288 338086 337300
rect 340233 337297 340245 337300
rect 340279 337297 340291 337331
rect 340233 337291 340291 337297
rect 341797 337331 341855 337337
rect 341797 337297 341809 337331
rect 341843 337328 341855 337331
rect 347130 337328 347136 337340
rect 341843 337300 347136 337328
rect 341843 337297 341855 337300
rect 341797 337291 341855 337297
rect 347130 337288 347136 337300
rect 347188 337288 347194 337340
rect 351178 337288 351184 337340
rect 351236 337328 351242 337340
rect 361482 337328 361488 337340
rect 351236 337300 361488 337328
rect 351236 337288 351242 337300
rect 361482 337288 361488 337300
rect 361540 337288 361546 337340
rect 375006 337288 375012 337340
rect 375064 337328 375070 337340
rect 381538 337328 381544 337340
rect 375064 337300 381544 337328
rect 375064 337288 375070 337300
rect 381538 337288 381544 337300
rect 381596 337288 381602 337340
rect 385310 337288 385316 337340
rect 385368 337328 385374 337340
rect 393225 337331 393283 337337
rect 393225 337328 393237 337331
rect 385368 337300 393237 337328
rect 385368 337288 385374 337300
rect 393225 337297 393237 337300
rect 393271 337297 393283 337331
rect 394620 337328 394648 337436
rect 394694 337424 394700 337476
rect 394752 337464 394758 337476
rect 395798 337464 395804 337476
rect 394752 337436 395804 337464
rect 394752 337424 394758 337436
rect 395798 337424 395804 337436
rect 395856 337424 395862 337476
rect 396905 337467 396963 337473
rect 396905 337433 396917 337467
rect 396951 337464 396963 337467
rect 402238 337464 402244 337476
rect 396951 337436 402244 337464
rect 396951 337433 396963 337436
rect 396905 337427 396963 337433
rect 402238 337424 402244 337436
rect 402296 337424 402302 337476
rect 415394 337424 415400 337476
rect 415452 337464 415458 337476
rect 416590 337464 416596 337476
rect 415452 337436 416596 337464
rect 415452 337424 415458 337436
rect 416590 337424 416596 337436
rect 416648 337424 416654 337476
rect 417053 337467 417111 337473
rect 417053 337433 417065 337467
rect 417099 337464 417111 337467
rect 428093 337467 428151 337473
rect 428093 337464 428105 337467
rect 417099 337436 428105 337464
rect 417099 337433 417111 337436
rect 417053 337427 417111 337433
rect 428093 337433 428105 337436
rect 428139 337433 428151 337467
rect 428200 337464 428228 337504
rect 428277 337501 428289 337535
rect 428323 337532 428335 337535
rect 433978 337532 433984 337544
rect 428323 337504 433984 337532
rect 428323 337501 428335 337504
rect 428277 337495 428335 337501
rect 433978 337492 433984 337504
rect 434036 337492 434042 337544
rect 442169 337535 442227 337541
rect 442169 337501 442181 337535
rect 442215 337532 442227 337535
rect 442905 337535 442963 337541
rect 442215 337504 442396 337532
rect 442215 337501 442227 337504
rect 442169 337495 442227 337501
rect 432693 337467 432751 337473
rect 432693 337464 432705 337467
rect 428200 337436 432705 337464
rect 428093 337427 428151 337433
rect 432693 337433 432705 337436
rect 432739 337433 432751 337467
rect 432693 337427 432751 337433
rect 433334 337424 433340 337476
rect 433392 337464 433398 337476
rect 435082 337464 435088 337476
rect 433392 337436 435088 337464
rect 433392 337424 433398 337436
rect 435082 337424 435088 337436
rect 435140 337424 435146 337476
rect 437017 337467 437075 337473
rect 437017 337433 437029 337467
rect 437063 337464 437075 337467
rect 442261 337467 442319 337473
rect 442261 337464 442273 337467
rect 437063 337436 442273 337464
rect 437063 337433 437075 337436
rect 437017 337427 437075 337433
rect 442261 337433 442273 337436
rect 442307 337433 442319 337467
rect 442368 337464 442396 337504
rect 442905 337501 442917 337535
rect 442951 337532 442963 337535
rect 444745 337535 444803 337541
rect 444745 337532 444757 337535
rect 442951 337504 444757 337532
rect 442951 337501 442963 337504
rect 442905 337495 442963 337501
rect 444745 337501 444757 337504
rect 444791 337501 444803 337535
rect 444745 337495 444803 337501
rect 444834 337492 444840 337544
rect 444892 337532 444898 337544
rect 525058 337532 525064 337544
rect 444892 337504 525064 337532
rect 444892 337492 444898 337504
rect 525058 337492 525064 337504
rect 525116 337492 525122 337544
rect 520918 337464 520924 337476
rect 442368 337436 520924 337464
rect 442261 337427 442319 337433
rect 520918 337424 520924 337436
rect 520976 337424 520982 337476
rect 394789 337399 394847 337405
rect 394789 337365 394801 337399
rect 394835 337396 394847 337399
rect 404998 337396 405004 337408
rect 394835 337368 405004 337396
rect 394835 337365 394847 337368
rect 394789 337359 394847 337365
rect 404998 337356 405004 337368
rect 405056 337356 405062 337408
rect 411346 337356 411352 337408
rect 411404 337396 411410 337408
rect 428277 337399 428335 337405
rect 428277 337396 428289 337399
rect 411404 337368 428289 337396
rect 411404 337356 411410 337368
rect 428277 337365 428289 337368
rect 428323 337365 428335 337399
rect 428277 337359 428335 337365
rect 428366 337356 428372 337408
rect 428424 337396 428430 337408
rect 429102 337396 429108 337408
rect 428424 337368 429108 337396
rect 428424 337356 428430 337368
rect 429102 337356 429108 337368
rect 429160 337356 429166 337408
rect 429746 337356 429752 337408
rect 429804 337396 429810 337408
rect 430482 337396 430488 337408
rect 429804 337368 430488 337396
rect 429804 337356 429810 337368
rect 430482 337356 430488 337368
rect 430540 337356 430546 337408
rect 431126 337356 431132 337408
rect 431184 337396 431190 337408
rect 431862 337396 431868 337408
rect 431184 337368 431868 337396
rect 431184 337356 431190 337368
rect 431862 337356 431868 337368
rect 431920 337356 431926 337408
rect 432414 337356 432420 337408
rect 432472 337396 432478 337408
rect 433242 337396 433248 337408
rect 432472 337368 433248 337396
rect 432472 337356 432478 337368
rect 433242 337356 433248 337368
rect 433300 337356 433306 337408
rect 433794 337356 433800 337408
rect 433852 337396 433858 337408
rect 434622 337396 434628 337408
rect 433852 337368 434628 337396
rect 433852 337356 433858 337368
rect 434622 337356 434628 337368
rect 434680 337356 434686 337408
rect 436002 337356 436008 337408
rect 436060 337396 436066 337408
rect 436830 337396 436836 337408
rect 436060 337368 436836 337396
rect 436060 337356 436066 337368
rect 436830 337356 436836 337368
rect 436888 337356 436894 337408
rect 437842 337356 437848 337408
rect 437900 337396 437906 337408
rect 438762 337396 438768 337408
rect 437900 337368 438768 337396
rect 437900 337356 437906 337368
rect 438762 337356 438768 337368
rect 438820 337356 438826 337408
rect 439130 337356 439136 337408
rect 439188 337396 439194 337408
rect 440050 337396 440056 337408
rect 439188 337368 440056 337396
rect 439188 337356 439194 337368
rect 440050 337356 440056 337368
rect 440108 337356 440114 337408
rect 440510 337356 440516 337408
rect 440568 337396 440574 337408
rect 441522 337396 441528 337408
rect 440568 337368 441528 337396
rect 440568 337356 440574 337368
rect 441522 337356 441528 337368
rect 441580 337356 441586 337408
rect 441890 337356 441896 337408
rect 441948 337396 441954 337408
rect 442810 337396 442816 337408
rect 441948 337368 442816 337396
rect 441948 337356 441954 337368
rect 442810 337356 442816 337368
rect 442868 337356 442874 337408
rect 443178 337356 443184 337408
rect 443236 337396 443242 337408
rect 444282 337396 444288 337408
rect 443236 337368 444288 337396
rect 443236 337356 443242 337368
rect 444282 337356 444288 337368
rect 444340 337356 444346 337408
rect 444558 337356 444564 337408
rect 444616 337396 444622 337408
rect 445570 337396 445576 337408
rect 444616 337368 445576 337396
rect 444616 337356 444622 337368
rect 445570 337356 445576 337368
rect 445628 337356 445634 337408
rect 445665 337399 445723 337405
rect 445665 337365 445677 337399
rect 445711 337396 445723 337399
rect 523678 337396 523684 337408
rect 445711 337368 523684 337396
rect 445711 337365 445723 337368
rect 445665 337359 445723 337365
rect 523678 337356 523684 337368
rect 523736 337356 523742 337408
rect 401870 337328 401876 337340
rect 394620 337300 401876 337328
rect 393225 337291 393283 337297
rect 401870 337288 401876 337300
rect 401928 337288 401934 337340
rect 426989 337331 427047 337337
rect 426989 337297 427001 337331
rect 427035 337328 427047 337331
rect 496078 337328 496084 337340
rect 427035 337300 496084 337328
rect 427035 337297 427047 337300
rect 426989 337291 427047 337297
rect 496078 337288 496084 337300
rect 496136 337288 496142 337340
rect 77996 337232 246160 337260
rect 77996 337220 78002 337232
rect 246298 337220 246304 337272
rect 246356 337260 246362 337272
rect 247034 337260 247040 337272
rect 246356 337232 247040 337260
rect 246356 337220 246362 337232
rect 247034 337220 247040 337232
rect 247092 337220 247098 337272
rect 247770 337220 247776 337272
rect 247828 337260 247834 337272
rect 248782 337260 248788 337272
rect 247828 337232 248788 337260
rect 247828 337220 247834 337232
rect 248782 337220 248788 337232
rect 248840 337220 248846 337272
rect 249058 337220 249064 337272
rect 249116 337260 249122 337272
rect 251542 337260 251548 337272
rect 249116 337232 251548 337260
rect 249116 337220 249122 337232
rect 251542 337220 251548 337232
rect 251600 337220 251606 337272
rect 253198 337220 253204 337272
rect 253256 337260 253262 337272
rect 259638 337260 259644 337272
rect 253256 337232 259644 337260
rect 253256 337220 253262 337232
rect 259638 337220 259644 337232
rect 259696 337220 259702 337272
rect 267001 337263 267059 337269
rect 267001 337229 267013 337263
rect 267047 337260 267059 337263
rect 299385 337263 299443 337269
rect 299385 337260 299397 337263
rect 267047 337232 299397 337260
rect 267047 337229 267059 337232
rect 267001 337223 267059 337229
rect 299385 337229 299397 337232
rect 299431 337229 299443 337263
rect 299385 337223 299443 337229
rect 299477 337263 299535 337269
rect 299477 337229 299489 337263
rect 299523 337260 299535 337263
rect 305822 337260 305828 337272
rect 299523 337232 305828 337260
rect 299523 337229 299535 337232
rect 299477 337223 299535 337229
rect 305822 337220 305828 337232
rect 305880 337220 305886 337272
rect 350718 337260 350724 337272
rect 326264 337232 350724 337260
rect 97258 337152 97264 337204
rect 97316 337192 97322 337204
rect 264974 337192 264980 337204
rect 97316 337164 264980 337192
rect 97316 337152 97322 337164
rect 264974 337152 264980 337164
rect 265032 337152 265038 337204
rect 297910 337152 297916 337204
rect 297968 337192 297974 337204
rect 303433 337195 303491 337201
rect 303433 337192 303445 337195
rect 297968 337164 303445 337192
rect 297968 337152 297974 337164
rect 303433 337161 303445 337164
rect 303479 337161 303491 337195
rect 303433 337155 303491 337161
rect 312722 337152 312728 337204
rect 312780 337192 312786 337204
rect 326157 337195 326215 337201
rect 326157 337192 326169 337195
rect 312780 337164 326169 337192
rect 312780 337152 312786 337164
rect 326157 337161 326169 337164
rect 326203 337161 326215 337195
rect 326157 337155 326215 337161
rect 84838 337084 84844 337136
rect 84896 337124 84902 337136
rect 89625 337127 89683 337133
rect 89625 337124 89637 337127
rect 84896 337096 89637 337124
rect 84896 337084 84902 337096
rect 89625 337093 89637 337096
rect 89671 337093 89683 337127
rect 89625 337087 89683 337093
rect 100662 337084 100668 337136
rect 100720 337124 100726 337136
rect 267642 337124 267648 337136
rect 100720 337096 267648 337124
rect 100720 337084 100726 337096
rect 267642 337084 267648 337096
rect 267700 337084 267706 337136
rect 321462 337084 321468 337136
rect 321520 337124 321526 337136
rect 326264 337124 326292 337232
rect 350718 337220 350724 337232
rect 350776 337220 350782 337272
rect 385957 337263 386015 337269
rect 385957 337229 385969 337263
rect 386003 337260 386015 337263
rect 392578 337260 392584 337272
rect 386003 337232 392584 337260
rect 386003 337229 386015 337232
rect 385957 337223 386015 337229
rect 392578 337220 392584 337232
rect 392636 337220 392642 337272
rect 408034 337220 408040 337272
rect 408092 337260 408098 337272
rect 417421 337263 417479 337269
rect 417421 337260 417433 337263
rect 408092 337232 417433 337260
rect 408092 337220 408098 337232
rect 417421 337229 417433 337232
rect 417467 337229 417479 337263
rect 417421 337223 417479 337229
rect 419902 337220 419908 337272
rect 419960 337260 419966 337272
rect 421558 337260 421564 337272
rect 419960 337232 421564 337260
rect 419960 337220 419966 337232
rect 421558 337220 421564 337232
rect 421616 337220 421622 337272
rect 427081 337263 427139 337269
rect 427081 337229 427093 337263
rect 427127 337260 427139 337263
rect 492674 337260 492680 337272
rect 427127 337232 492680 337260
rect 427127 337229 427139 337232
rect 427081 337223 427139 337229
rect 492674 337220 492680 337232
rect 492732 337220 492738 337272
rect 326341 337195 326399 337201
rect 326341 337161 326353 337195
rect 326387 337192 326399 337195
rect 341334 337192 341340 337204
rect 326387 337164 341340 337192
rect 326387 337161 326399 337164
rect 326341 337155 326399 337161
rect 341334 337152 341340 337164
rect 341392 337152 341398 337204
rect 345658 337152 345664 337204
rect 345716 337192 345722 337204
rect 354766 337192 354772 337204
rect 345716 337164 354772 337192
rect 345716 337152 345722 337164
rect 354766 337152 354772 337164
rect 354824 337152 354830 337204
rect 362865 337195 362923 337201
rect 362865 337161 362877 337195
rect 362911 337192 362923 337195
rect 365530 337192 365536 337204
rect 362911 337164 365536 337192
rect 362911 337161 362923 337164
rect 362865 337155 362923 337161
rect 365530 337152 365536 337164
rect 365588 337152 365594 337204
rect 370498 337152 370504 337204
rect 370556 337192 370562 337204
rect 372706 337192 372712 337204
rect 370556 337164 372712 337192
rect 370556 337152 370562 337164
rect 372706 337152 372712 337164
rect 372764 337152 372770 337204
rect 383841 337195 383899 337201
rect 383841 337161 383853 337195
rect 383887 337192 383899 337195
rect 388533 337195 388591 337201
rect 388533 337192 388545 337195
rect 383887 337164 388545 337192
rect 383887 337161 383899 337164
rect 383841 337155 383899 337161
rect 388533 337161 388545 337164
rect 388579 337161 388591 337195
rect 388533 337155 388591 337161
rect 413094 337152 413100 337204
rect 413152 337192 413158 337204
rect 485774 337192 485780 337204
rect 413152 337164 485780 337192
rect 413152 337152 413158 337164
rect 485774 337152 485780 337164
rect 485832 337152 485838 337204
rect 343082 337124 343088 337136
rect 321520 337096 326292 337124
rect 326356 337096 343088 337124
rect 321520 337084 321526 337096
rect 107562 337016 107568 337068
rect 107620 337056 107626 337068
rect 270402 337056 270408 337068
rect 107620 337028 270408 337056
rect 107620 337016 107626 337028
rect 270402 337016 270408 337028
rect 270460 337016 270466 337068
rect 299385 337059 299443 337065
rect 299385 337025 299397 337059
rect 299431 337056 299443 337059
rect 299477 337059 299535 337065
rect 299477 337056 299489 337059
rect 299431 337028 299489 337056
rect 299431 337025 299443 337028
rect 299385 337019 299443 337025
rect 299477 337025 299489 337028
rect 299523 337025 299535 337059
rect 299477 337019 299535 337025
rect 105538 336948 105544 337000
rect 105596 336988 105602 337000
rect 262306 336988 262312 337000
rect 105596 336960 262312 336988
rect 105596 336948 105602 336960
rect 262306 336948 262312 336960
rect 262364 336948 262370 337000
rect 319530 336948 319536 337000
rect 319588 336988 319594 337000
rect 326356 336988 326384 337096
rect 343082 337084 343088 337096
rect 343140 337084 343146 337136
rect 346670 337124 346676 337136
rect 343192 337096 346676 337124
rect 326433 337059 326491 337065
rect 326433 337025 326445 337059
rect 326479 337056 326491 337059
rect 336553 337059 336611 337065
rect 336553 337056 336565 337059
rect 326479 337028 336565 337056
rect 326479 337025 326491 337028
rect 326433 337019 326491 337025
rect 336553 337025 336565 337028
rect 336599 337025 336611 337059
rect 336553 337019 336611 337025
rect 336645 337059 336703 337065
rect 336645 337025 336657 337059
rect 336691 337056 336703 337059
rect 339034 337056 339040 337068
rect 336691 337028 339040 337056
rect 336691 337025 336703 337028
rect 336645 337019 336703 337025
rect 339034 337016 339040 337028
rect 339092 337016 339098 337068
rect 343192 337056 343220 337096
rect 346670 337084 346676 337096
rect 346728 337084 346734 337136
rect 358722 337084 358728 337136
rect 358780 337124 358786 337136
rect 365070 337124 365076 337136
rect 358780 337096 365076 337124
rect 358780 337084 358786 337096
rect 365070 337084 365076 337096
rect 365128 337084 365134 337136
rect 393406 337084 393412 337136
rect 393464 337124 393470 337136
rect 394510 337124 394516 337136
rect 393464 337096 394516 337124
rect 393464 337084 393470 337096
rect 394510 337084 394516 337096
rect 394568 337084 394574 337136
rect 399662 337084 399668 337136
rect 399720 337124 399726 337136
rect 407761 337127 407819 337133
rect 407761 337124 407773 337127
rect 399720 337096 407773 337124
rect 399720 337084 399726 337096
rect 407761 337093 407773 337096
rect 407807 337093 407819 337127
rect 407761 337087 407819 337093
rect 410426 337084 410432 337136
rect 410484 337124 410490 337136
rect 477494 337124 477500 337136
rect 410484 337096 477500 337124
rect 410484 337084 410490 337096
rect 477494 337084 477500 337096
rect 477552 337084 477558 337136
rect 341904 337028 343220 337056
rect 345569 337059 345627 337065
rect 319588 336960 326384 336988
rect 319588 336948 319594 336960
rect 327718 336948 327724 337000
rect 327776 336988 327782 337000
rect 341705 336991 341763 336997
rect 341705 336988 341717 336991
rect 327776 336960 341717 336988
rect 327776 336948 327782 336960
rect 341705 336957 341717 336960
rect 341751 336957 341763 336991
rect 341705 336951 341763 336957
rect 99377 336923 99435 336929
rect 99377 336889 99389 336923
rect 99423 336920 99435 336923
rect 108945 336923 109003 336929
rect 108945 336920 108957 336923
rect 99423 336892 108957 336920
rect 99423 336889 99435 336892
rect 99377 336883 99435 336889
rect 108945 336889 108957 336892
rect 108991 336889 109003 336923
rect 108945 336883 109003 336889
rect 118602 336880 118608 336932
rect 118660 336920 118666 336932
rect 274450 336920 274456 336932
rect 118660 336892 274456 336920
rect 118660 336880 118666 336892
rect 274450 336880 274456 336892
rect 274508 336880 274514 336932
rect 316770 336880 316776 336932
rect 316828 336920 316834 336932
rect 336645 336923 336703 336929
rect 336645 336920 336657 336923
rect 316828 336892 336657 336920
rect 316828 336880 316834 336892
rect 336645 336889 336657 336892
rect 336691 336889 336703 336923
rect 341797 336923 341855 336929
rect 341797 336920 341809 336923
rect 336645 336883 336703 336889
rect 336752 336892 341809 336920
rect 102778 336812 102784 336864
rect 102836 336852 102842 336864
rect 255590 336852 255596 336864
rect 102836 336824 255596 336852
rect 102836 336812 102842 336824
rect 255590 336812 255596 336824
rect 255648 336812 255654 336864
rect 326338 336812 326344 336864
rect 326396 336852 326402 336864
rect 336752 336852 336780 336892
rect 341797 336889 341809 336892
rect 341843 336889 341855 336923
rect 341797 336883 341855 336889
rect 326396 336824 336780 336852
rect 326396 336812 326402 336824
rect 338758 336812 338764 336864
rect 338816 336852 338822 336864
rect 341904 336852 341932 337028
rect 345569 337025 345581 337059
rect 345615 337056 345627 337059
rect 353846 337056 353852 337068
rect 345615 337028 353852 337056
rect 345615 337025 345627 337028
rect 345569 337019 345627 337025
rect 353846 337016 353852 337028
rect 353904 337016 353910 337068
rect 359458 337016 359464 337068
rect 359516 337056 359522 337068
rect 364610 337056 364616 337068
rect 359516 337028 364616 337056
rect 359516 337016 359522 337028
rect 364610 337016 364616 337028
rect 364668 337016 364674 337068
rect 371786 337016 371792 337068
rect 371844 337056 371850 337068
rect 375650 337056 375656 337068
rect 371844 337028 375656 337056
rect 371844 337016 371850 337028
rect 375650 337016 375656 337028
rect 375708 337016 375714 337068
rect 389818 337016 389824 337068
rect 389876 337056 389882 337068
rect 390370 337056 390376 337068
rect 389876 337028 390376 337056
rect 389876 337016 389882 337028
rect 390370 337016 390376 337028
rect 390428 337016 390434 337068
rect 409966 337016 409972 337068
rect 410024 337056 410030 337068
rect 477586 337056 477592 337068
rect 410024 337028 477592 337056
rect 410024 337016 410030 337028
rect 477586 337016 477592 337028
rect 477644 337016 477650 337068
rect 341978 336948 341984 337000
rect 342036 336988 342042 337000
rect 348050 336988 348056 337000
rect 342036 336960 348056 336988
rect 342036 336948 342042 336960
rect 348050 336948 348056 336960
rect 348108 336948 348114 337000
rect 360102 336948 360108 337000
rect 360160 336988 360166 337000
rect 362865 336991 362923 336997
rect 362865 336988 362877 336991
rect 360160 336960 362877 336988
rect 360160 336948 360166 336960
rect 362865 336957 362877 336960
rect 362911 336957 362923 336991
rect 362865 336951 362923 336957
rect 364242 336948 364248 337000
rect 364300 336988 364306 337000
rect 366910 336988 366916 337000
rect 364300 336960 366916 336988
rect 364300 336948 364306 336960
rect 366910 336948 366916 336960
rect 366968 336948 366974 337000
rect 417421 336991 417479 336997
rect 417421 336957 417433 336991
rect 417467 336988 417479 336991
rect 470594 336988 470600 337000
rect 417467 336960 470600 336988
rect 417467 336957 417479 336960
rect 417421 336951 417479 336957
rect 470594 336948 470600 336960
rect 470652 336948 470658 337000
rect 344738 336880 344744 336932
rect 344796 336920 344802 336932
rect 350258 336920 350264 336932
rect 344796 336892 350264 336920
rect 344796 336880 344802 336892
rect 350258 336880 350264 336892
rect 350316 336880 350322 336932
rect 366358 336880 366364 336932
rect 366416 336920 366422 336932
rect 367370 336920 367376 336932
rect 366416 336892 367376 336920
rect 366416 336880 366422 336892
rect 367370 336880 367376 336892
rect 367428 336880 367434 336932
rect 373626 336880 373632 336932
rect 373684 336920 373690 336932
rect 374638 336920 374644 336932
rect 373684 336892 374644 336920
rect 373684 336880 373690 336892
rect 374638 336880 374644 336892
rect 374696 336880 374702 336932
rect 402330 336880 402336 336932
rect 402388 336920 402394 336932
rect 402388 336892 403204 336920
rect 402388 336880 402394 336892
rect 338816 336824 341932 336852
rect 338816 336812 338822 336824
rect 344646 336812 344652 336864
rect 344704 336852 344710 336864
rect 349338 336852 349344 336864
rect 344704 336824 349344 336852
rect 344704 336812 344710 336824
rect 349338 336812 349344 336824
rect 349396 336812 349402 336864
rect 362218 336812 362224 336864
rect 362276 336852 362282 336864
rect 365990 336852 365996 336864
rect 362276 336824 365996 336852
rect 362276 336812 362282 336824
rect 365990 336812 365996 336824
rect 366048 336812 366054 336864
rect 366910 336812 366916 336864
rect 366968 336852 366974 336864
rect 367830 336852 367836 336864
rect 366968 336824 367836 336852
rect 366968 336812 366974 336824
rect 367830 336812 367836 336824
rect 367888 336812 367894 336864
rect 403176 336852 403204 336892
rect 405366 336880 405372 336932
rect 405424 336920 405430 336932
rect 463694 336920 463700 336932
rect 405424 336892 463700 336920
rect 405424 336880 405430 336892
rect 463694 336880 463700 336892
rect 463752 336880 463758 336932
rect 456794 336852 456800 336864
rect 403176 336824 456800 336852
rect 456794 336812 456800 336824
rect 456852 336812 456858 336864
rect 118697 336787 118755 336793
rect 118697 336753 118709 336787
rect 118743 336784 118755 336787
rect 118743 336756 125456 336784
rect 118743 336753 118755 336756
rect 118697 336747 118755 336753
rect 125428 336716 125456 336756
rect 125502 336744 125508 336796
rect 125560 336784 125566 336796
rect 277118 336784 277124 336796
rect 125560 336756 277124 336784
rect 125560 336744 125566 336756
rect 277118 336744 277124 336756
rect 277176 336744 277182 336796
rect 322290 336744 322296 336796
rect 322348 336784 322354 336796
rect 326433 336787 326491 336793
rect 326433 336784 326445 336787
rect 322348 336756 326445 336784
rect 322348 336744 322354 336756
rect 326433 336753 326445 336756
rect 326479 336753 326491 336787
rect 326433 336747 326491 336753
rect 327810 336744 327816 336796
rect 327868 336784 327874 336796
rect 342622 336784 342628 336796
rect 327868 336756 342628 336784
rect 327868 336744 327874 336756
rect 342622 336744 342628 336756
rect 342680 336744 342686 336796
rect 345477 336787 345535 336793
rect 345477 336753 345489 336787
rect 345523 336784 345535 336787
rect 354306 336784 354312 336796
rect 345523 336756 354312 336784
rect 345523 336753 345535 336756
rect 345477 336747 345535 336753
rect 354306 336744 354312 336756
rect 354364 336744 354370 336796
rect 362862 336744 362868 336796
rect 362920 336784 362926 336796
rect 366450 336784 366456 336796
rect 362920 336756 366456 336784
rect 362920 336744 362926 336756
rect 366450 336744 366456 336756
rect 366508 336744 366514 336796
rect 367002 336744 367008 336796
rect 367060 336784 367066 336796
rect 368198 336784 368204 336796
rect 367060 336756 368204 336784
rect 367060 336744 367066 336756
rect 368198 336744 368204 336756
rect 368256 336744 368262 336796
rect 407761 336787 407819 336793
rect 407761 336753 407773 336787
rect 407807 336784 407819 336787
rect 437569 336787 437627 336793
rect 437569 336784 437581 336787
rect 407807 336756 437581 336784
rect 407807 336753 407819 336756
rect 407761 336747 407819 336753
rect 437569 336753 437581 336756
rect 437615 336753 437627 336787
rect 437569 336747 437627 336753
rect 437753 336787 437811 336793
rect 437753 336753 437765 336787
rect 437799 336784 437811 336787
rect 447045 336787 447103 336793
rect 437799 336756 446996 336784
rect 437799 336753 437811 336756
rect 437753 336747 437811 336753
rect 128265 336719 128323 336725
rect 128265 336716 128277 336719
rect 125428 336688 128277 336716
rect 128265 336685 128277 336688
rect 128311 336685 128323 336719
rect 239122 336716 239128 336728
rect 239083 336688 239128 336716
rect 128265 336679 128323 336685
rect 239122 336676 239128 336688
rect 239180 336676 239186 336728
rect 324682 336716 324688 336728
rect 324643 336688 324688 336716
rect 324682 336676 324688 336688
rect 324740 336676 324746 336728
rect 428093 336719 428151 336725
rect 428093 336685 428105 336719
rect 428139 336716 428151 336719
rect 435358 336716 435364 336728
rect 428139 336688 435364 336716
rect 428139 336685 428151 336688
rect 428093 336679 428151 336685
rect 435358 336676 435364 336688
rect 435416 336676 435422 336728
rect 446968 336716 446996 336756
rect 447045 336753 447057 336787
rect 447091 336784 447103 336787
rect 449989 336787 450047 336793
rect 449989 336784 450001 336787
rect 447091 336756 450001 336784
rect 447091 336753 447103 336756
rect 447045 336747 447103 336753
rect 449989 336753 450001 336756
rect 450035 336753 450047 336787
rect 449989 336747 450047 336753
rect 449894 336716 449900 336728
rect 446968 336688 449900 336716
rect 449894 336676 449900 336688
rect 449952 336676 449958 336728
rect 437293 336651 437351 336657
rect 437293 336617 437305 336651
rect 437339 336648 437351 336651
rect 438118 336648 438124 336660
rect 437339 336620 438124 336648
rect 437339 336617 437351 336620
rect 437293 336611 437351 336617
rect 438118 336608 438124 336620
rect 438176 336608 438182 336660
rect 435269 336515 435327 336521
rect 435269 336481 435281 336515
rect 435315 336512 435327 336515
rect 442258 336512 442264 336524
rect 435315 336484 442264 336512
rect 435315 336481 435327 336484
rect 435269 336475 435327 336481
rect 442258 336472 442264 336484
rect 442316 336472 442322 336524
rect 311894 335724 311900 335776
rect 311952 335764 311958 335776
rect 312262 335764 312268 335776
rect 311952 335736 312268 335764
rect 311952 335724 311958 335736
rect 312262 335724 312268 335736
rect 312320 335724 312326 335776
rect 232038 335656 232044 335708
rect 232096 335696 232102 335708
rect 232774 335696 232780 335708
rect 232096 335668 232780 335696
rect 232096 335656 232102 335668
rect 232774 335656 232780 335668
rect 232832 335656 232838 335708
rect 277394 335656 277400 335708
rect 277452 335696 277458 335708
rect 278130 335696 278136 335708
rect 277452 335668 278136 335696
rect 277452 335656 277458 335668
rect 278130 335656 278136 335668
rect 278188 335656 278194 335708
rect 285858 335656 285864 335708
rect 285916 335696 285922 335708
rect 286686 335696 286692 335708
rect 285916 335668 286692 335696
rect 285916 335656 285922 335668
rect 286686 335656 286692 335668
rect 286744 335656 286750 335708
rect 303706 335656 303712 335708
rect 303764 335696 303770 335708
rect 304626 335696 304632 335708
rect 303764 335668 304632 335696
rect 303764 335656 303770 335668
rect 304626 335656 304632 335668
rect 304684 335656 304690 335708
rect 306466 335656 306472 335708
rect 306524 335696 306530 335708
rect 307294 335696 307300 335708
rect 306524 335668 307300 335696
rect 306524 335656 306530 335668
rect 307294 335656 307300 335668
rect 307352 335656 307358 335708
rect 317414 335656 317420 335708
rect 317472 335696 317478 335708
rect 317598 335696 317604 335708
rect 317472 335668 317604 335696
rect 317472 335656 317478 335668
rect 317598 335656 317604 335668
rect 317656 335656 317662 335708
rect 323026 335656 323032 335708
rect 323084 335696 323090 335708
rect 323486 335696 323492 335708
rect 323084 335668 323492 335696
rect 323084 335656 323090 335668
rect 323486 335656 323492 335668
rect 323544 335656 323550 335708
rect 231946 335588 231952 335640
rect 232004 335628 232010 335640
rect 232406 335628 232412 335640
rect 232004 335600 232412 335628
rect 232004 335588 232010 335600
rect 232406 335588 232412 335600
rect 232464 335588 232470 335640
rect 234706 335588 234712 335640
rect 234764 335628 234770 335640
rect 234982 335628 234988 335640
rect 234764 335600 234988 335628
rect 234764 335588 234770 335600
rect 234982 335588 234988 335600
rect 235040 335588 235046 335640
rect 236086 335588 236092 335640
rect 236144 335628 236150 335640
rect 236454 335628 236460 335640
rect 236144 335600 236460 335628
rect 236144 335588 236150 335600
rect 236454 335588 236460 335600
rect 236512 335588 236518 335640
rect 237466 335588 237472 335640
rect 237524 335628 237530 335640
rect 238110 335628 238116 335640
rect 237524 335600 238116 335628
rect 237524 335588 237530 335600
rect 238110 335588 238116 335600
rect 238168 335588 238174 335640
rect 241514 335588 241520 335640
rect 241572 335628 241578 335640
rect 241790 335628 241796 335640
rect 241572 335600 241796 335628
rect 241572 335588 241578 335600
rect 241790 335588 241796 335600
rect 241848 335588 241854 335640
rect 247126 335588 247132 335640
rect 247184 335628 247190 335640
rect 247678 335628 247684 335640
rect 247184 335600 247684 335628
rect 247184 335588 247190 335600
rect 247678 335588 247684 335600
rect 247736 335588 247742 335640
rect 249886 335588 249892 335640
rect 249944 335628 249950 335640
rect 250806 335628 250812 335640
rect 249944 335600 250812 335628
rect 249944 335588 249950 335600
rect 250806 335588 250812 335600
rect 250864 335588 250870 335640
rect 251266 335588 251272 335640
rect 251324 335628 251330 335640
rect 252094 335628 252100 335640
rect 251324 335600 252100 335628
rect 251324 335588 251330 335600
rect 252094 335588 252100 335600
rect 252152 335588 252158 335640
rect 252646 335588 252652 335640
rect 252704 335628 252710 335640
rect 253382 335628 253388 335640
rect 252704 335600 253388 335628
rect 252704 335588 252710 335600
rect 253382 335588 253388 335600
rect 253440 335588 253446 335640
rect 255406 335588 255412 335640
rect 255464 335628 255470 335640
rect 256142 335628 256148 335640
rect 255464 335600 256148 335628
rect 255464 335588 255470 335600
rect 256142 335588 256148 335600
rect 256200 335588 256206 335640
rect 258166 335588 258172 335640
rect 258224 335628 258230 335640
rect 258902 335628 258908 335640
rect 258224 335600 258908 335628
rect 258224 335588 258230 335600
rect 258902 335588 258908 335600
rect 258960 335588 258966 335640
rect 259546 335588 259552 335640
rect 259604 335628 259610 335640
rect 260190 335628 260196 335640
rect 259604 335600 260196 335628
rect 259604 335588 259610 335600
rect 260190 335588 260196 335600
rect 260248 335588 260254 335640
rect 263686 335588 263692 335640
rect 263744 335628 263750 335640
rect 264238 335628 264244 335640
rect 263744 335600 264244 335628
rect 263744 335588 263750 335600
rect 264238 335588 264244 335600
rect 264296 335588 264302 335640
rect 266446 335588 266452 335640
rect 266504 335628 266510 335640
rect 266998 335628 267004 335640
rect 266504 335600 267004 335628
rect 266504 335588 266510 335600
rect 266998 335588 267004 335600
rect 267056 335588 267062 335640
rect 267826 335588 267832 335640
rect 267884 335628 267890 335640
rect 268286 335628 268292 335640
rect 267884 335600 268292 335628
rect 267884 335588 267890 335600
rect 268286 335588 268292 335600
rect 268344 335588 268350 335640
rect 269206 335588 269212 335640
rect 269264 335628 269270 335640
rect 269574 335628 269580 335640
rect 269264 335600 269580 335628
rect 269264 335588 269270 335600
rect 269574 335588 269580 335600
rect 269632 335588 269638 335640
rect 271966 335588 271972 335640
rect 272024 335628 272030 335640
rect 272334 335628 272340 335640
rect 272024 335600 272340 335628
rect 272024 335588 272030 335600
rect 272334 335588 272340 335600
rect 272392 335588 272398 335640
rect 274726 335588 274732 335640
rect 274784 335628 274790 335640
rect 274910 335628 274916 335640
rect 274784 335600 274916 335628
rect 274784 335588 274790 335600
rect 274910 335588 274916 335600
rect 274968 335588 274974 335640
rect 277486 335588 277492 335640
rect 277544 335628 277550 335640
rect 277670 335628 277676 335640
rect 277544 335600 277676 335628
rect 277544 335588 277550 335600
rect 277670 335588 277676 335600
rect 277728 335588 277734 335640
rect 278958 335588 278964 335640
rect 279016 335628 279022 335640
rect 279510 335628 279516 335640
rect 279016 335600 279516 335628
rect 279016 335588 279022 335600
rect 279510 335588 279516 335600
rect 279568 335588 279574 335640
rect 281718 335588 281724 335640
rect 281776 335628 281782 335640
rect 282178 335628 282184 335640
rect 281776 335600 282184 335628
rect 281776 335588 281782 335600
rect 282178 335588 282184 335600
rect 282236 335588 282242 335640
rect 283006 335588 283012 335640
rect 283064 335628 283070 335640
rect 283558 335628 283564 335640
rect 283064 335600 283564 335628
rect 283064 335588 283070 335600
rect 283558 335588 283564 335600
rect 283616 335588 283622 335640
rect 285766 335588 285772 335640
rect 285824 335628 285830 335640
rect 286134 335628 286140 335640
rect 285824 335600 286140 335628
rect 285824 335588 285830 335600
rect 286134 335588 286140 335600
rect 286192 335588 286198 335640
rect 294046 335588 294052 335640
rect 294104 335628 294110 335640
rect 294782 335628 294788 335640
rect 294104 335600 294788 335628
rect 294104 335588 294110 335600
rect 294782 335588 294788 335600
rect 294840 335588 294846 335640
rect 296806 335588 296812 335640
rect 296864 335628 296870 335640
rect 297358 335628 297364 335640
rect 296864 335600 297364 335628
rect 296864 335588 296870 335600
rect 297358 335588 297364 335600
rect 297416 335588 297422 335640
rect 302326 335588 302332 335640
rect 302384 335628 302390 335640
rect 302878 335628 302884 335640
rect 302384 335600 302884 335628
rect 302384 335588 302390 335600
rect 302878 335588 302884 335600
rect 302936 335588 302942 335640
rect 303798 335588 303804 335640
rect 303856 335628 303862 335640
rect 304166 335628 304172 335640
rect 303856 335600 304172 335628
rect 303856 335588 303862 335600
rect 304166 335588 304172 335600
rect 304224 335588 304230 335640
rect 306374 335588 306380 335640
rect 306432 335628 306438 335640
rect 306926 335628 306932 335640
rect 306432 335600 306932 335628
rect 306432 335588 306438 335600
rect 306926 335588 306932 335600
rect 306984 335588 306990 335640
rect 307754 335588 307760 335640
rect 307812 335628 307818 335640
rect 308214 335628 308220 335640
rect 307812 335600 308220 335628
rect 307812 335588 307818 335600
rect 308214 335588 308220 335600
rect 308272 335588 308278 335640
rect 309134 335588 309140 335640
rect 309192 335628 309198 335640
rect 309502 335628 309508 335640
rect 309192 335600 309508 335628
rect 309192 335588 309198 335600
rect 309502 335588 309508 335600
rect 309560 335588 309566 335640
rect 310514 335588 310520 335640
rect 310572 335628 310578 335640
rect 310974 335628 310980 335640
rect 310572 335600 310980 335628
rect 310572 335588 310578 335600
rect 310974 335588 310980 335600
rect 311032 335588 311038 335640
rect 313274 335588 313280 335640
rect 313332 335628 313338 335640
rect 313550 335628 313556 335640
rect 313332 335600 313556 335628
rect 313332 335588 313338 335600
rect 313550 335588 313556 335600
rect 313608 335588 313614 335640
rect 320266 335588 320272 335640
rect 320324 335628 320330 335640
rect 320726 335628 320732 335640
rect 320324 335600 320732 335628
rect 320324 335588 320330 335600
rect 320726 335588 320732 335600
rect 320784 335588 320790 335640
rect 321646 335588 321652 335640
rect 321704 335628 321710 335640
rect 322198 335628 322204 335640
rect 321704 335600 322204 335628
rect 321704 335588 321710 335600
rect 322198 335588 322204 335600
rect 322256 335588 322262 335640
rect 323210 335588 323216 335640
rect 323268 335628 323274 335640
rect 323854 335628 323860 335640
rect 323268 335600 323860 335628
rect 323268 335588 323274 335600
rect 323854 335588 323860 335600
rect 323912 335588 323918 335640
rect 325786 335588 325792 335640
rect 325844 335628 325850 335640
rect 326614 335628 326620 335640
rect 325844 335600 326620 335628
rect 325844 335588 325850 335600
rect 326614 335588 326620 335600
rect 326672 335588 326678 335640
rect 327166 335588 327172 335640
rect 327224 335628 327230 335640
rect 327902 335628 327908 335640
rect 327224 335600 327908 335628
rect 327224 335588 327230 335600
rect 327902 335588 327908 335600
rect 327960 335588 327966 335640
rect 329926 335588 329932 335640
rect 329984 335628 329990 335640
rect 330294 335628 330300 335640
rect 329984 335600 330300 335628
rect 329984 335588 329990 335600
rect 330294 335588 330300 335600
rect 330352 335588 330358 335640
rect 345106 335588 345112 335640
rect 345164 335628 345170 335640
rect 345934 335628 345940 335640
rect 345164 335600 345940 335628
rect 345164 335588 345170 335600
rect 345934 335588 345940 335600
rect 345992 335588 345998 335640
rect 435450 335588 435456 335640
rect 435508 335628 435514 335640
rect 436002 335628 436008 335640
rect 435508 335600 436008 335628
rect 435508 335588 435514 335600
rect 436002 335588 436008 335600
rect 436060 335588 436066 335640
rect 343821 335563 343879 335569
rect 343821 335529 343833 335563
rect 343867 335560 343879 335563
rect 344554 335560 344560 335572
rect 343867 335532 344560 335560
rect 343867 335529 343879 335532
rect 343821 335523 343879 335529
rect 344554 335520 344560 335532
rect 344612 335520 344618 335572
rect 273530 335424 273536 335436
rect 273456 335396 273536 335424
rect 273456 335232 273484 335396
rect 273530 335384 273536 335396
rect 273588 335384 273594 335436
rect 314654 335248 314660 335300
rect 314712 335288 314718 335300
rect 315022 335288 315028 335300
rect 314712 335260 315028 335288
rect 314712 335248 314718 335260
rect 315022 335248 315028 335260
rect 315080 335248 315086 335300
rect 273438 335180 273444 335232
rect 273496 335180 273502 335232
rect 324406 334976 324412 335028
rect 324464 335016 324470 335028
rect 325326 335016 325332 335028
rect 324464 334988 325332 335016
rect 324464 334976 324470 334988
rect 325326 334976 325332 334988
rect 325384 334976 325390 335028
rect 233513 334475 233571 334481
rect 233513 334441 233525 334475
rect 233559 334472 233571 334475
rect 234062 334472 234068 334484
rect 233559 334444 234068 334472
rect 233559 334441 233571 334444
rect 233513 334435 233571 334441
rect 234062 334432 234068 334444
rect 234120 334432 234126 334484
rect 265066 334296 265072 334348
rect 265124 334336 265130 334348
rect 265526 334336 265532 334348
rect 265124 334308 265532 334336
rect 265124 334296 265130 334308
rect 265526 334296 265532 334308
rect 265584 334296 265590 334348
rect 287425 334339 287483 334345
rect 287425 334305 287437 334339
rect 287471 334336 287483 334339
rect 287974 334336 287980 334348
rect 287471 334308 287980 334336
rect 287471 334305 287483 334308
rect 287425 334299 287483 334305
rect 287974 334296 287980 334308
rect 288032 334296 288038 334348
rect 312170 334296 312176 334348
rect 312228 334336 312234 334348
rect 312630 334336 312636 334348
rect 312228 334308 312636 334336
rect 312228 334296 312234 334308
rect 312630 334296 312636 334308
rect 312688 334296 312694 334348
rect 319165 334203 319223 334209
rect 319165 334169 319177 334203
rect 319211 334200 319223 334203
rect 319438 334200 319444 334212
rect 319211 334172 319444 334200
rect 319211 334169 319223 334172
rect 319165 334163 319223 334169
rect 319438 334160 319444 334172
rect 319496 334160 319502 334212
rect 256786 334024 256792 334076
rect 256844 334064 256850 334076
rect 257430 334064 257436 334076
rect 256844 334036 257436 334064
rect 256844 334024 256850 334036
rect 257430 334024 257436 334036
rect 257488 334024 257494 334076
rect 238662 333276 238668 333328
rect 238720 333316 238726 333328
rect 239030 333316 239036 333328
rect 238720 333288 239036 333316
rect 238720 333276 238726 333288
rect 239030 333276 239036 333288
rect 239088 333276 239094 333328
rect 273346 333276 273352 333328
rect 273404 333316 273410 333328
rect 273622 333316 273628 333328
rect 273404 333288 273628 333316
rect 273404 333276 273410 333288
rect 273622 333276 273628 333288
rect 273680 333276 273686 333328
rect 347866 333276 347872 333328
rect 347924 333316 347930 333328
rect 348694 333316 348700 333328
rect 347924 333288 348700 333316
rect 347924 333276 347930 333288
rect 348694 333276 348700 333288
rect 348752 333276 348758 333328
rect 284386 333140 284392 333192
rect 284444 333180 284450 333192
rect 284846 333180 284852 333192
rect 284444 333152 284852 333180
rect 284444 333140 284450 333152
rect 284846 333140 284852 333152
rect 284904 333140 284910 333192
rect 318794 333140 318800 333192
rect 318852 333180 318858 333192
rect 319070 333180 319076 333192
rect 318852 333152 319076 333180
rect 318852 333140 318858 333152
rect 319070 333140 319076 333152
rect 319128 333140 319134 333192
rect 300946 332800 300952 332852
rect 301004 332840 301010 332852
rect 301406 332840 301412 332852
rect 301004 332812 301412 332840
rect 301004 332800 301010 332812
rect 301406 332800 301412 332812
rect 301464 332800 301470 332852
rect 248598 332392 248604 332444
rect 248656 332432 248662 332444
rect 249334 332432 249340 332444
rect 248656 332404 249340 332432
rect 248656 332392 248662 332404
rect 249334 332392 249340 332404
rect 249392 332392 249398 332444
rect 235077 331959 235135 331965
rect 235077 331925 235089 331959
rect 235123 331956 235135 331959
rect 235442 331956 235448 331968
rect 235123 331928 235448 331956
rect 235123 331925 235135 331928
rect 235077 331919 235135 331925
rect 235442 331916 235448 331928
rect 235500 331916 235506 331968
rect 295426 331576 295432 331628
rect 295484 331616 295490 331628
rect 296070 331616 296076 331628
rect 295484 331588 296076 331616
rect 295484 331576 295490 331588
rect 296070 331576 296076 331588
rect 296128 331576 296134 331628
rect 298462 331440 298468 331492
rect 298520 331480 298526 331492
rect 298922 331480 298928 331492
rect 298520 331452 298928 331480
rect 298520 331440 298526 331452
rect 298922 331440 298928 331452
rect 298980 331440 298986 331492
rect 244458 331344 244464 331356
rect 244292 331316 244464 331344
rect 244292 331220 244320 331316
rect 244458 331304 244464 331316
rect 244516 331304 244522 331356
rect 244366 331236 244372 331288
rect 244424 331236 244430 331288
rect 244274 331168 244280 331220
rect 244332 331168 244338 331220
rect 244384 331152 244412 331236
rect 327442 331208 327448 331220
rect 327403 331180 327448 331208
rect 327442 331168 327448 331180
rect 327500 331168 327506 331220
rect 244366 331100 244372 331152
rect 244424 331100 244430 331152
rect 316034 330964 316040 331016
rect 316092 331004 316098 331016
rect 316310 331004 316316 331016
rect 316092 330976 316316 331004
rect 316092 330964 316098 330976
rect 316310 330964 316316 330976
rect 316368 330964 316374 331016
rect 314930 330216 314936 330268
rect 314988 330256 314994 330268
rect 315390 330256 315396 330268
rect 314988 330228 315396 330256
rect 314988 330216 314994 330228
rect 315390 330216 315396 330228
rect 315448 330216 315454 330268
rect 290458 329400 290464 329452
rect 290516 329440 290522 329452
rect 294049 329443 294107 329449
rect 294049 329440 294061 329443
rect 290516 329412 294061 329440
rect 290516 329400 290522 329412
rect 294049 329409 294061 329412
rect 294095 329409 294107 329443
rect 294049 329403 294107 329409
rect 233510 328488 233516 328500
rect 233471 328460 233516 328488
rect 233510 328448 233516 328460
rect 233568 328448 233574 328500
rect 262674 328448 262680 328500
rect 262732 328488 262738 328500
rect 263042 328488 263048 328500
rect 262732 328460 263048 328488
rect 262732 328448 262738 328460
rect 263042 328448 263048 328460
rect 263100 328448 263106 328500
rect 266998 328488 267004 328500
rect 266959 328460 267004 328488
rect 266998 328448 267004 328460
rect 267056 328448 267062 328500
rect 288802 328448 288808 328500
rect 288860 328488 288866 328500
rect 289538 328488 289544 328500
rect 288860 328460 289544 328488
rect 288860 328448 288866 328460
rect 289538 328448 289544 328460
rect 289596 328448 289602 328500
rect 289998 328448 290004 328500
rect 290056 328488 290062 328500
rect 290642 328488 290648 328500
rect 290056 328460 290648 328488
rect 290056 328448 290062 328460
rect 290642 328448 290648 328460
rect 290700 328448 290706 328500
rect 291562 328448 291568 328500
rect 291620 328488 291626 328500
rect 292114 328488 292120 328500
rect 291620 328460 292120 328488
rect 291620 328448 291626 328460
rect 292114 328448 292120 328460
rect 292172 328448 292178 328500
rect 292758 328448 292764 328500
rect 292816 328488 292822 328500
rect 293586 328488 293592 328500
rect 292816 328460 293592 328488
rect 292816 328448 292822 328460
rect 293586 328448 293592 328460
rect 293644 328448 293650 328500
rect 305362 328448 305368 328500
rect 305420 328488 305426 328500
rect 306098 328488 306104 328500
rect 305420 328460 306104 328488
rect 305420 328448 305426 328460
rect 306098 328448 306104 328460
rect 306156 328448 306162 328500
rect 308122 328448 308128 328500
rect 308180 328488 308186 328500
rect 308674 328488 308680 328500
rect 308180 328460 308680 328488
rect 308180 328448 308186 328460
rect 308674 328448 308680 328460
rect 308732 328448 308738 328500
rect 310882 328448 310888 328500
rect 310940 328488 310946 328500
rect 311434 328488 311440 328500
rect 310940 328460 311440 328488
rect 310940 328448 310946 328460
rect 311434 328448 311440 328460
rect 311492 328448 311498 328500
rect 316402 328448 316408 328500
rect 316460 328488 316466 328500
rect 316586 328488 316592 328500
rect 316460 328460 316592 328488
rect 316460 328448 316466 328460
rect 316586 328448 316592 328460
rect 316644 328448 316650 328500
rect 319162 328488 319168 328500
rect 319123 328460 319168 328488
rect 319162 328448 319168 328460
rect 319220 328448 319226 328500
rect 327442 328488 327448 328500
rect 327403 328460 327448 328488
rect 327442 328448 327448 328460
rect 327500 328448 327506 328500
rect 328546 328448 328552 328500
rect 328604 328488 328610 328500
rect 328822 328488 328828 328500
rect 328604 328460 328828 328488
rect 328604 328448 328610 328460
rect 328822 328448 328828 328460
rect 328880 328448 328886 328500
rect 343818 328488 343824 328500
rect 343779 328460 343824 328488
rect 343818 328448 343824 328460
rect 343876 328448 343882 328500
rect 346578 328448 346584 328500
rect 346636 328488 346642 328500
rect 347314 328488 347320 328500
rect 346636 328460 347320 328488
rect 346636 328448 346642 328460
rect 347314 328448 347320 328460
rect 347372 328448 347378 328500
rect 347958 328488 347964 328500
rect 347919 328460 347964 328488
rect 347958 328448 347964 328460
rect 348016 328448 348022 328500
rect 251450 328380 251456 328432
rect 251508 328420 251514 328432
rect 251634 328420 251640 328432
rect 251508 328392 251640 328420
rect 251508 328380 251514 328392
rect 251634 328380 251640 328392
rect 251692 328380 251698 328432
rect 254210 328380 254216 328432
rect 254268 328420 254274 328432
rect 254302 328420 254308 328432
rect 254268 328392 254308 328420
rect 254268 328380 254274 328392
rect 254302 328380 254308 328392
rect 254360 328380 254366 328432
rect 363230 328420 363236 328432
rect 363191 328392 363236 328420
rect 363230 328380 363236 328392
rect 363288 328380 363294 328432
rect 324685 328355 324743 328361
rect 324685 328321 324697 328355
rect 324731 328352 324743 328355
rect 324774 328352 324780 328364
rect 324731 328324 324780 328352
rect 324731 328321 324743 328324
rect 324685 328315 324743 328321
rect 324774 328312 324780 328324
rect 324832 328312 324838 328364
rect 347958 328352 347964 328364
rect 347919 328324 347964 328352
rect 347958 328312 347964 328324
rect 348016 328312 348022 328364
rect 235074 327128 235080 327140
rect 235035 327100 235080 327128
rect 235074 327088 235080 327100
rect 235132 327088 235138 327140
rect 240410 327088 240416 327140
rect 240468 327128 240474 327140
rect 240870 327128 240876 327140
rect 240468 327100 240876 327128
rect 240468 327088 240474 327100
rect 240870 327088 240876 327100
rect 240928 327088 240934 327140
rect 241882 327088 241888 327140
rect 241940 327128 241946 327140
rect 242158 327128 242164 327140
rect 241940 327100 242164 327128
rect 241940 327088 241946 327100
rect 242158 327088 242164 327100
rect 242216 327088 242222 327140
rect 245930 327088 245936 327140
rect 245988 327128 245994 327140
rect 246206 327128 246212 327140
rect 245988 327100 246212 327128
rect 245988 327088 245994 327100
rect 246206 327088 246212 327100
rect 246264 327088 246270 327140
rect 287422 327128 287428 327140
rect 287383 327100 287428 327128
rect 287422 327088 287428 327100
rect 287480 327088 287486 327140
rect 234798 327060 234804 327072
rect 234759 327032 234804 327060
rect 234798 327020 234804 327032
rect 234856 327020 234862 327072
rect 248874 325660 248880 325712
rect 248932 325700 248938 325712
rect 249242 325700 249248 325712
rect 248932 325672 249248 325700
rect 248932 325660 248938 325672
rect 249242 325660 249248 325672
rect 249300 325660 249306 325712
rect 577590 322872 577596 322924
rect 577648 322912 577654 322924
rect 579890 322912 579896 322924
rect 577648 322884 579896 322912
rect 577648 322872 577654 322884
rect 579890 322872 579896 322884
rect 579948 322872 579954 322924
rect 248782 322192 248788 322244
rect 248840 322232 248846 322244
rect 249242 322232 249248 322244
rect 248840 322204 249248 322232
rect 248840 322192 248846 322204
rect 249242 322192 249248 322204
rect 249300 322192 249306 322244
rect 255682 321580 255688 321632
rect 255740 321580 255746 321632
rect 261202 321580 261208 321632
rect 261260 321580 261266 321632
rect 267090 321620 267096 321632
rect 267016 321592 267096 321620
rect 229278 321512 229284 321564
rect 229336 321552 229342 321564
rect 229462 321552 229468 321564
rect 229336 321524 229468 321552
rect 229336 321512 229342 321524
rect 229462 321512 229468 321524
rect 229520 321512 229526 321564
rect 238754 321512 238760 321564
rect 238812 321552 238818 321564
rect 238938 321552 238944 321564
rect 238812 321524 238944 321552
rect 238812 321512 238818 321524
rect 238938 321512 238944 321524
rect 238996 321512 239002 321564
rect 255700 321428 255728 321580
rect 255682 321376 255688 321428
rect 255740 321376 255746 321428
rect 261220 321416 261248 321580
rect 267016 321428 267044 321592
rect 267090 321580 267096 321592
rect 267148 321580 267154 321632
rect 289998 321580 290004 321632
rect 290056 321580 290062 321632
rect 292758 321580 292764 321632
rect 292816 321580 292822 321632
rect 325970 321580 325976 321632
rect 326028 321580 326034 321632
rect 290016 321484 290044 321580
rect 290090 321484 290096 321496
rect 290016 321456 290096 321484
rect 290090 321444 290096 321456
rect 290148 321444 290154 321496
rect 292776 321484 292804 321580
rect 292850 321484 292856 321496
rect 292776 321456 292856 321484
rect 292850 321444 292856 321456
rect 292908 321444 292914 321496
rect 261294 321416 261300 321428
rect 261220 321388 261300 321416
rect 261294 321376 261300 321388
rect 261352 321376 261358 321428
rect 266998 321376 267004 321428
rect 267056 321376 267062 321428
rect 325988 321416 326016 321580
rect 326062 321416 326068 321428
rect 325988 321388 326068 321416
rect 326062 321376 326068 321388
rect 326120 321376 326126 321428
rect 251634 318900 251640 318912
rect 251468 318872 251640 318900
rect 239122 318832 239128 318844
rect 239083 318804 239128 318832
rect 239122 318792 239128 318804
rect 239180 318792 239186 318844
rect 251468 318776 251496 318872
rect 251634 318860 251640 318872
rect 251692 318860 251698 318912
rect 316402 318900 316408 318912
rect 316328 318872 316408 318900
rect 280522 318792 280528 318844
rect 280580 318832 280586 318844
rect 280614 318832 280620 318844
rect 280580 318804 280620 318832
rect 280580 318792 280586 318804
rect 280614 318792 280620 318804
rect 280672 318792 280678 318844
rect 316328 318776 316356 318872
rect 316402 318860 316408 318872
rect 316460 318860 316466 318912
rect 317874 318900 317880 318912
rect 317800 318872 317880 318900
rect 317800 318844 317828 318872
rect 317874 318860 317880 318872
rect 317932 318860 317938 318912
rect 317782 318792 317788 318844
rect 317840 318792 317846 318844
rect 347958 318832 347964 318844
rect 347919 318804 347964 318832
rect 347958 318792 347964 318804
rect 348016 318792 348022 318844
rect 363233 318835 363291 318841
rect 363233 318801 363245 318835
rect 363279 318832 363291 318835
rect 363322 318832 363328 318844
rect 363279 318804 363328 318832
rect 363279 318801 363291 318804
rect 363233 318795 363291 318801
rect 363322 318792 363328 318804
rect 363380 318792 363386 318844
rect 434346 318792 434352 318844
rect 434404 318832 434410 318844
rect 434438 318832 434444 318844
rect 434404 318804 434444 318832
rect 434404 318792 434410 318804
rect 434438 318792 434444 318804
rect 434496 318792 434502 318844
rect 444098 318792 444104 318844
rect 444156 318832 444162 318844
rect 444190 318832 444196 318844
rect 444156 318804 444196 318832
rect 444156 318792 444162 318804
rect 444190 318792 444196 318804
rect 444248 318792 444254 318844
rect 251450 318724 251456 318776
rect 251508 318724 251514 318776
rect 262674 318764 262680 318776
rect 262635 318736 262680 318764
rect 262674 318724 262680 318736
rect 262732 318724 262738 318776
rect 292850 318764 292856 318776
rect 292811 318736 292856 318764
rect 292850 318724 292856 318736
rect 292908 318724 292914 318776
rect 298462 318724 298468 318776
rect 298520 318764 298526 318776
rect 298554 318764 298560 318776
rect 298520 318736 298560 318764
rect 298520 318724 298526 318736
rect 298554 318724 298560 318736
rect 298612 318724 298618 318776
rect 316310 318724 316316 318776
rect 316368 318724 316374 318776
rect 327442 318764 327448 318776
rect 327403 318736 327448 318764
rect 327442 318724 327448 318736
rect 327500 318724 327506 318776
rect 328546 318724 328552 318776
rect 328604 318764 328610 318776
rect 328730 318764 328736 318776
rect 328604 318736 328736 318764
rect 328604 318724 328610 318736
rect 328730 318724 328736 318736
rect 328788 318724 328794 318776
rect 342530 318764 342536 318776
rect 342491 318736 342536 318764
rect 342530 318724 342536 318736
rect 342588 318724 342594 318776
rect 345198 318764 345204 318776
rect 345159 318736 345204 318764
rect 345198 318724 345204 318736
rect 345256 318724 345262 318776
rect 324590 318656 324596 318708
rect 324648 318696 324654 318708
rect 324774 318696 324780 318708
rect 324648 318668 324780 318696
rect 324648 318656 324654 318668
rect 324774 318656 324780 318668
rect 324832 318656 324838 318708
rect 234801 317475 234859 317481
rect 234801 317441 234813 317475
rect 234847 317472 234859 317475
rect 234890 317472 234896 317484
rect 234847 317444 234896 317472
rect 234847 317441 234859 317444
rect 234801 317435 234859 317441
rect 234890 317432 234896 317444
rect 234948 317432 234954 317484
rect 287330 317404 287336 317416
rect 287291 317376 287336 317404
rect 287330 317364 287336 317376
rect 287388 317364 287394 317416
rect 298462 317404 298468 317416
rect 298423 317376 298468 317404
rect 298462 317364 298468 317376
rect 298520 317364 298526 317416
rect 435358 316684 435364 316736
rect 435416 316724 435422 316736
rect 435542 316724 435548 316736
rect 435416 316696 435548 316724
rect 435416 316684 435422 316696
rect 435542 316684 435548 316696
rect 435600 316684 435606 316736
rect 249978 316072 249984 316124
rect 250036 316112 250042 316124
rect 250162 316112 250168 316124
rect 250036 316084 250168 316112
rect 250036 316072 250042 316084
rect 250162 316072 250168 316084
rect 250220 316072 250226 316124
rect 250073 315979 250131 315985
rect 250073 315945 250085 315979
rect 250119 315976 250131 315979
rect 250162 315976 250168 315988
rect 250119 315948 250168 315976
rect 250119 315945 250131 315948
rect 250073 315939 250131 315945
rect 250162 315936 250168 315948
rect 250220 315936 250226 315988
rect 290090 315908 290096 315920
rect 290051 315880 290096 315908
rect 290090 315868 290096 315880
rect 290148 315868 290154 315920
rect 229462 313896 229468 313948
rect 229520 313936 229526 313948
rect 229646 313936 229652 313948
rect 229520 313908 229652 313936
rect 229520 313896 229526 313908
rect 229646 313896 229652 313908
rect 229704 313896 229710 313948
rect 305362 312740 305368 312792
rect 305420 312780 305426 312792
rect 305638 312780 305644 312792
rect 305420 312752 305644 312780
rect 305420 312740 305426 312752
rect 305638 312740 305644 312752
rect 305696 312740 305702 312792
rect 262674 312168 262680 312180
rect 262635 312140 262680 312168
rect 262674 312128 262680 312140
rect 262732 312128 262738 312180
rect 248785 311967 248843 311973
rect 248785 311933 248797 311967
rect 248831 311964 248843 311967
rect 248874 311964 248880 311976
rect 248831 311936 248880 311964
rect 248831 311933 248843 311936
rect 248785 311927 248843 311933
rect 248874 311924 248880 311936
rect 248932 311924 248938 311976
rect 444098 311924 444104 311976
rect 444156 311964 444162 311976
rect 444190 311964 444196 311976
rect 444156 311936 444196 311964
rect 444156 311924 444162 311936
rect 444190 311924 444196 311936
rect 444248 311924 444254 311976
rect 328638 311856 328644 311908
rect 328696 311856 328702 311908
rect 287330 311828 287336 311840
rect 287291 311800 287336 311828
rect 287330 311788 287336 311800
rect 287388 311788 287394 311840
rect 328656 311704 328684 311856
rect 328638 311652 328644 311704
rect 328696 311652 328702 311704
rect 238846 309748 238852 309800
rect 238904 309748 238910 309800
rect 238864 309664 238892 309748
rect 238846 309612 238852 309664
rect 238904 309612 238910 309664
rect 347958 309272 347964 309324
rect 348016 309272 348022 309324
rect 347976 309188 348004 309272
rect 266906 309136 266912 309188
rect 266964 309176 266970 309188
rect 266998 309176 267004 309188
rect 266964 309148 267004 309176
rect 266964 309136 266970 309148
rect 266998 309136 267004 309148
rect 267056 309136 267062 309188
rect 291470 309136 291476 309188
rect 291528 309176 291534 309188
rect 291562 309176 291568 309188
rect 291528 309148 291568 309176
rect 291528 309136 291534 309148
rect 291562 309136 291568 309148
rect 291620 309136 291626 309188
rect 292850 309176 292856 309188
rect 292811 309148 292856 309176
rect 292850 309136 292856 309148
rect 292908 309136 292914 309188
rect 327442 309176 327448 309188
rect 327403 309148 327448 309176
rect 327442 309136 327448 309148
rect 327500 309136 327506 309188
rect 342530 309176 342536 309188
rect 342491 309148 342536 309176
rect 342530 309136 342536 309148
rect 342588 309136 342594 309188
rect 345201 309179 345259 309185
rect 345201 309145 345213 309179
rect 345247 309176 345259 309179
rect 345290 309176 345296 309188
rect 345247 309148 345296 309176
rect 345247 309145 345259 309148
rect 345201 309139 345259 309145
rect 345290 309136 345296 309148
rect 345348 309136 345354 309188
rect 347958 309136 347964 309188
rect 348016 309136 348022 309188
rect 362954 309136 362960 309188
rect 363012 309176 363018 309188
rect 363322 309176 363328 309188
rect 363012 309148 363328 309176
rect 363012 309136 363018 309148
rect 363322 309136 363328 309148
rect 363380 309136 363386 309188
rect 229462 309068 229468 309120
rect 229520 309108 229526 309120
rect 229646 309108 229652 309120
rect 229520 309080 229652 309108
rect 229520 309068 229526 309080
rect 229646 309068 229652 309080
rect 229704 309068 229710 309120
rect 235074 309108 235080 309120
rect 235035 309080 235080 309108
rect 235074 309068 235080 309080
rect 235132 309068 235138 309120
rect 308030 309068 308036 309120
rect 308088 309108 308094 309120
rect 308214 309108 308220 309120
rect 308088 309080 308220 309108
rect 308088 309068 308094 309080
rect 308214 309068 308220 309080
rect 308272 309068 308278 309120
rect 434257 309111 434315 309117
rect 434257 309077 434269 309111
rect 434303 309108 434315 309111
rect 434530 309108 434536 309120
rect 434303 309080 434536 309108
rect 434303 309077 434315 309080
rect 434257 309071 434315 309077
rect 434530 309068 434536 309080
rect 434588 309068 434594 309120
rect 266998 309040 267004 309052
rect 266959 309012 267004 309040
rect 266998 309000 267004 309012
rect 267056 309000 267062 309052
rect 347958 309040 347964 309052
rect 347919 309012 347964 309040
rect 347958 309000 347964 309012
rect 348016 309000 348022 309052
rect 290093 307819 290151 307825
rect 290093 307785 290105 307819
rect 290139 307816 290151 307819
rect 290274 307816 290280 307828
rect 290139 307788 290280 307816
rect 290139 307785 290151 307788
rect 290093 307779 290151 307785
rect 290274 307776 290280 307788
rect 290332 307776 290338 307828
rect 298462 307816 298468 307828
rect 298423 307788 298468 307816
rect 298462 307776 298468 307788
rect 298520 307776 298526 307828
rect 234890 307748 234896 307760
rect 234851 307720 234896 307748
rect 234890 307708 234896 307720
rect 234948 307708 234954 307760
rect 305457 307751 305515 307757
rect 305457 307717 305469 307751
rect 305503 307748 305515 307751
rect 305546 307748 305552 307760
rect 305503 307720 305552 307748
rect 305503 307717 305515 307720
rect 305457 307711 305515 307717
rect 305546 307708 305552 307720
rect 305604 307708 305610 307760
rect 316310 307748 316316 307760
rect 316271 307720 316316 307748
rect 316310 307708 316316 307720
rect 316368 307708 316374 307760
rect 342438 307748 342444 307760
rect 342399 307720 342444 307748
rect 342438 307708 342444 307720
rect 342496 307708 342502 307760
rect 254118 306416 254124 306468
rect 254176 306456 254182 306468
rect 254302 306456 254308 306468
rect 254176 306428 254308 306456
rect 254176 306416 254182 306428
rect 254302 306416 254308 306428
rect 254360 306416 254366 306468
rect 313458 306348 313464 306400
rect 313516 306388 313522 306400
rect 313550 306388 313556 306400
rect 313516 306360 313556 306388
rect 313516 306348 313522 306360
rect 313550 306348 313556 306360
rect 313608 306348 313614 306400
rect 288710 302268 288716 302320
rect 288768 302268 288774 302320
rect 233326 302200 233332 302252
rect 233384 302240 233390 302252
rect 233510 302240 233516 302252
rect 233384 302212 233516 302240
rect 233384 302200 233390 302212
rect 233510 302200 233516 302212
rect 233568 302200 233574 302252
rect 280430 302200 280436 302252
rect 280488 302240 280494 302252
rect 280614 302240 280620 302252
rect 280488 302212 280620 302240
rect 280488 302200 280494 302212
rect 280614 302200 280620 302212
rect 280672 302200 280678 302252
rect 288728 302184 288756 302268
rect 435358 302200 435364 302252
rect 435416 302240 435422 302252
rect 435542 302240 435548 302252
rect 435416 302212 435548 302240
rect 435416 302200 435422 302212
rect 435542 302200 435548 302212
rect 435600 302200 435606 302252
rect 444006 302200 444012 302252
rect 444064 302240 444070 302252
rect 444190 302240 444196 302252
rect 444064 302212 444196 302240
rect 444064 302200 444070 302212
rect 444190 302200 444196 302212
rect 444248 302200 444254 302252
rect 288710 302132 288716 302184
rect 288768 302132 288774 302184
rect 362954 302064 362960 302116
rect 363012 302104 363018 302116
rect 363230 302104 363236 302116
rect 363012 302076 363236 302104
rect 363012 302064 363018 302076
rect 363230 302064 363236 302076
rect 363288 302064 363294 302116
rect 229281 299591 229339 299597
rect 229281 299557 229293 299591
rect 229327 299588 229339 299591
rect 229462 299588 229468 299600
rect 229327 299560 229468 299588
rect 229327 299557 229339 299560
rect 229281 299551 229339 299557
rect 229462 299548 229468 299560
rect 229520 299548 229526 299600
rect 244182 299548 244188 299600
rect 244240 299588 244246 299600
rect 347958 299588 347964 299600
rect 244240 299560 244320 299588
rect 347919 299560 347964 299588
rect 244240 299548 244246 299560
rect 244292 299532 244320 299560
rect 347958 299548 347964 299560
rect 348016 299548 348022 299600
rect 235074 299520 235080 299532
rect 235035 299492 235080 299520
rect 235074 299480 235080 299492
rect 235132 299480 235138 299532
rect 244274 299480 244280 299532
rect 244332 299480 244338 299532
rect 248782 299520 248788 299532
rect 248743 299492 248788 299520
rect 248782 299480 248788 299492
rect 248840 299480 248846 299532
rect 250070 299520 250076 299532
rect 250031 299492 250076 299520
rect 250070 299480 250076 299492
rect 250128 299480 250134 299532
rect 267001 299523 267059 299529
rect 267001 299489 267013 299523
rect 267047 299520 267059 299523
rect 267274 299520 267280 299532
rect 267047 299492 267280 299520
rect 267047 299489 267059 299492
rect 267001 299483 267059 299489
rect 267274 299480 267280 299492
rect 267332 299480 267338 299532
rect 290090 299480 290096 299532
rect 290148 299520 290154 299532
rect 290274 299520 290280 299532
rect 290148 299492 290280 299520
rect 290148 299480 290154 299492
rect 290274 299480 290280 299492
rect 290332 299480 290338 299532
rect 434254 299520 434260 299532
rect 434215 299492 434260 299520
rect 434254 299480 434260 299492
rect 434312 299480 434318 299532
rect 262585 299455 262643 299461
rect 262585 299421 262597 299455
rect 262631 299452 262643 299455
rect 262674 299452 262680 299464
rect 262631 299424 262680 299452
rect 262631 299421 262643 299424
rect 262585 299415 262643 299421
rect 262674 299412 262680 299424
rect 262732 299412 262738 299464
rect 287330 299452 287336 299464
rect 287291 299424 287336 299452
rect 287330 299412 287336 299424
rect 287388 299412 287394 299464
rect 291470 299412 291476 299464
rect 291528 299452 291534 299464
rect 291562 299452 291568 299464
rect 291528 299424 291568 299452
rect 291528 299412 291534 299424
rect 291562 299412 291568 299424
rect 291620 299412 291626 299464
rect 298465 299455 298523 299461
rect 298465 299421 298477 299455
rect 298511 299452 298523 299455
rect 298554 299452 298560 299464
rect 298511 299424 298560 299452
rect 298511 299421 298523 299424
rect 298465 299415 298523 299421
rect 298554 299412 298560 299424
rect 298612 299412 298618 299464
rect 324593 299455 324651 299461
rect 324593 299421 324605 299455
rect 324639 299452 324651 299455
rect 324682 299452 324688 299464
rect 324639 299424 324688 299452
rect 324639 299421 324651 299424
rect 324593 299415 324651 299421
rect 324682 299412 324688 299424
rect 324740 299412 324746 299464
rect 327258 299412 327264 299464
rect 327316 299452 327322 299464
rect 327442 299452 327448 299464
rect 327316 299424 327448 299452
rect 327316 299412 327322 299424
rect 327442 299412 327448 299424
rect 327500 299412 327506 299464
rect 347958 299412 347964 299464
rect 348016 299452 348022 299464
rect 348050 299452 348056 299464
rect 348016 299424 348056 299452
rect 348016 299412 348022 299424
rect 348050 299412 348056 299424
rect 348108 299412 348114 299464
rect 577498 299412 577504 299464
rect 577556 299452 577562 299464
rect 579890 299452 579896 299464
rect 577556 299424 579896 299452
rect 577556 299412 577562 299424
rect 579890 299412 579896 299424
rect 579948 299412 579954 299464
rect 229278 298160 229284 298172
rect 229239 298132 229284 298160
rect 229278 298120 229284 298132
rect 229336 298120 229342 298172
rect 234890 298160 234896 298172
rect 234851 298132 234896 298160
rect 234890 298120 234896 298132
rect 234948 298120 234954 298172
rect 305454 298160 305460 298172
rect 305415 298132 305460 298160
rect 305454 298120 305460 298132
rect 305512 298120 305518 298172
rect 310793 298163 310851 298169
rect 310793 298129 310805 298163
rect 310839 298160 310851 298163
rect 310882 298160 310888 298172
rect 310839 298132 310888 298160
rect 310839 298129 310851 298132
rect 310793 298123 310851 298129
rect 310882 298120 310888 298132
rect 310940 298120 310946 298172
rect 316310 298160 316316 298172
rect 316271 298132 316316 298160
rect 316310 298120 316316 298132
rect 316368 298120 316374 298172
rect 342441 298163 342499 298169
rect 342441 298129 342453 298163
rect 342487 298160 342499 298163
rect 342530 298160 342536 298172
rect 342487 298132 342536 298160
rect 342487 298129 342499 298132
rect 342441 298123 342499 298129
rect 342530 298120 342536 298132
rect 342588 298120 342594 298172
rect 235074 298092 235080 298104
rect 235035 298064 235080 298092
rect 235074 298052 235080 298064
rect 235132 298052 235138 298104
rect 239030 298052 239036 298104
rect 239088 298092 239094 298104
rect 239122 298092 239128 298104
rect 239088 298064 239128 298092
rect 239088 298052 239094 298064
rect 239122 298052 239128 298064
rect 239180 298052 239186 298104
rect 240410 298092 240416 298104
rect 240371 298064 240416 298092
rect 240410 298052 240416 298064
rect 240468 298052 240474 298104
rect 241882 298092 241888 298104
rect 241843 298064 241888 298092
rect 241882 298052 241888 298064
rect 241940 298052 241946 298104
rect 291470 298092 291476 298104
rect 291431 298064 291476 298092
rect 291470 298052 291476 298064
rect 291528 298052 291534 298104
rect 308122 298052 308128 298104
rect 308180 298092 308186 298104
rect 308214 298092 308220 298104
rect 308180 298064 308220 298092
rect 308180 298052 308186 298064
rect 308214 298052 308220 298064
rect 308272 298052 308278 298104
rect 327258 298092 327264 298104
rect 327219 298064 327264 298092
rect 327258 298052 327264 298064
rect 327316 298052 327322 298104
rect 435358 297372 435364 297424
rect 435416 297412 435422 297424
rect 435542 297412 435548 297424
rect 435416 297384 435548 297412
rect 435416 297372 435422 297384
rect 435542 297372 435548 297384
rect 435600 297372 435606 297424
rect 253934 296692 253940 296744
rect 253992 296732 253998 296744
rect 254210 296732 254216 296744
rect 253992 296704 254216 296732
rect 253992 296692 253998 296704
rect 254210 296692 254216 296704
rect 254268 296692 254274 296744
rect 310790 296732 310796 296744
rect 310751 296704 310796 296732
rect 310790 296692 310796 296704
rect 310848 296692 310854 296744
rect 310790 295740 310796 295792
rect 310848 295780 310854 295792
rect 310974 295780 310980 295792
rect 310848 295752 310980 295780
rect 310848 295740 310854 295752
rect 310974 295740 310980 295752
rect 311032 295740 311038 295792
rect 2774 295196 2780 295248
rect 2832 295236 2838 295248
rect 5258 295236 5264 295248
rect 2832 295208 5264 295236
rect 2832 295196 2838 295208
rect 5258 295196 5264 295208
rect 5316 295196 5322 295248
rect 325973 294695 326031 294701
rect 325973 294661 325985 294695
rect 326019 294692 326031 294695
rect 326062 294692 326068 294704
rect 326019 294664 326068 294692
rect 326019 294661 326031 294664
rect 325973 294655 326031 294661
rect 326062 294652 326068 294664
rect 326120 294652 326126 294704
rect 254210 292612 254216 292664
rect 254268 292612 254274 292664
rect 342530 292612 342536 292664
rect 342588 292612 342594 292664
rect 254228 292528 254256 292612
rect 266998 292544 267004 292596
rect 267056 292584 267062 292596
rect 267274 292584 267280 292596
rect 267056 292556 267280 292584
rect 267056 292544 267062 292556
rect 267274 292544 267280 292556
rect 267332 292544 267338 292596
rect 328546 292544 328552 292596
rect 328604 292584 328610 292596
rect 328730 292584 328736 292596
rect 328604 292556 328736 292584
rect 328604 292544 328610 292556
rect 328730 292544 328736 292556
rect 328788 292544 328794 292596
rect 342548 292528 342576 292612
rect 254210 292476 254216 292528
rect 254268 292476 254274 292528
rect 342530 292476 342536 292528
rect 342588 292476 342594 292528
rect 229370 292408 229376 292460
rect 229428 292448 229434 292460
rect 229554 292448 229560 292460
rect 229428 292420 229560 292448
rect 229428 292408 229434 292420
rect 229554 292408 229560 292420
rect 229612 292408 229618 292460
rect 262582 289932 262588 289944
rect 262543 289904 262588 289932
rect 262582 289892 262588 289904
rect 262640 289892 262646 289944
rect 324590 289932 324596 289944
rect 324551 289904 324596 289932
rect 324590 289892 324596 289904
rect 324648 289892 324654 289944
rect 261202 289824 261208 289876
rect 261260 289864 261266 289876
rect 261294 289864 261300 289876
rect 261260 289836 261300 289864
rect 261260 289824 261266 289836
rect 261294 289824 261300 289836
rect 261352 289824 261358 289876
rect 287330 289864 287336 289876
rect 287291 289836 287336 289864
rect 287330 289824 287336 289836
rect 287388 289824 287394 289876
rect 288710 289824 288716 289876
rect 288768 289864 288774 289876
rect 288986 289864 288992 289876
rect 288768 289836 288992 289864
rect 288768 289824 288774 289836
rect 288986 289824 288992 289836
rect 289044 289824 289050 289876
rect 298462 289864 298468 289876
rect 298423 289836 298468 289864
rect 298462 289824 298468 289836
rect 298520 289824 298526 289876
rect 305454 289824 305460 289876
rect 305512 289824 305518 289876
rect 325970 289864 325976 289876
rect 325931 289836 325976 289864
rect 325970 289824 325976 289836
rect 326028 289824 326034 289876
rect 266998 289756 267004 289808
rect 267056 289796 267062 289808
rect 267274 289796 267280 289808
rect 267056 289768 267280 289796
rect 267056 289756 267062 289768
rect 267274 289756 267280 289768
rect 267332 289756 267338 289808
rect 305472 289740 305500 289824
rect 324590 289756 324596 289808
rect 324648 289756 324654 289808
rect 345198 289796 345204 289808
rect 345159 289768 345204 289796
rect 345198 289756 345204 289768
rect 345256 289756 345262 289808
rect 347774 289756 347780 289808
rect 347832 289796 347838 289808
rect 347958 289796 347964 289808
rect 347832 289768 347964 289796
rect 347832 289756 347838 289768
rect 347958 289756 347964 289768
rect 348016 289756 348022 289808
rect 434257 289799 434315 289805
rect 434257 289765 434269 289799
rect 434303 289796 434315 289799
rect 434346 289796 434352 289808
rect 434303 289768 434352 289796
rect 434303 289765 434315 289768
rect 434257 289759 434315 289765
rect 434346 289756 434352 289768
rect 434404 289756 434410 289808
rect 288710 289728 288716 289740
rect 288671 289700 288716 289728
rect 288710 289688 288716 289700
rect 288768 289688 288774 289740
rect 305454 289688 305460 289740
rect 305512 289688 305518 289740
rect 324608 289728 324636 289756
rect 324774 289728 324780 289740
rect 324608 289700 324780 289728
rect 324774 289688 324780 289700
rect 324832 289688 324838 289740
rect 316221 288507 316279 288513
rect 316221 288473 316233 288507
rect 316267 288504 316279 288507
rect 316310 288504 316316 288516
rect 316267 288476 316316 288504
rect 316267 288473 316279 288476
rect 316221 288467 316279 288473
rect 316310 288464 316316 288476
rect 316368 288464 316374 288516
rect 240410 288436 240416 288448
rect 240371 288408 240416 288436
rect 240410 288396 240416 288408
rect 240468 288396 240474 288448
rect 241882 288436 241888 288448
rect 241843 288408 241888 288436
rect 241882 288396 241888 288408
rect 241940 288396 241946 288448
rect 291470 288436 291476 288448
rect 291431 288408 291476 288436
rect 291470 288396 291476 288408
rect 291528 288396 291534 288448
rect 327261 288439 327319 288445
rect 327261 288405 327273 288439
rect 327307 288436 327319 288439
rect 327534 288436 327540 288448
rect 327307 288408 327540 288436
rect 327307 288405 327319 288408
rect 327261 288399 327319 288405
rect 327534 288396 327540 288408
rect 327592 288396 327598 288448
rect 262493 288371 262551 288377
rect 262493 288337 262505 288371
rect 262539 288368 262551 288371
rect 262582 288368 262588 288380
rect 262539 288340 262588 288368
rect 262539 288337 262551 288340
rect 262493 288331 262551 288337
rect 262582 288328 262588 288340
rect 262640 288328 262646 288380
rect 316218 287076 316224 287088
rect 316179 287048 316224 287076
rect 316218 287036 316224 287048
rect 316276 287036 316282 287088
rect 229370 282956 229376 283008
rect 229428 282956 229434 283008
rect 229388 282804 229416 282956
rect 233326 282888 233332 282940
rect 233384 282928 233390 282940
rect 233510 282928 233516 282940
rect 233384 282900 233516 282928
rect 233384 282888 233390 282900
rect 233510 282888 233516 282900
rect 233568 282888 233574 282940
rect 280430 282888 280436 282940
rect 280488 282928 280494 282940
rect 280614 282928 280620 282940
rect 280488 282900 280620 282928
rect 280488 282888 280494 282900
rect 280614 282888 280620 282900
rect 280672 282888 280678 282940
rect 298462 282888 298468 282940
rect 298520 282888 298526 282940
rect 435358 282888 435364 282940
rect 435416 282928 435422 282940
rect 435542 282928 435548 282940
rect 435416 282900 435548 282928
rect 435416 282888 435422 282900
rect 435542 282888 435548 282900
rect 435600 282888 435606 282940
rect 444006 282888 444012 282940
rect 444064 282928 444070 282940
rect 444190 282928 444196 282940
rect 444064 282900 444196 282928
rect 444064 282888 444070 282900
rect 444190 282888 444196 282900
rect 444248 282888 444254 282940
rect 288710 282860 288716 282872
rect 288671 282832 288716 282860
rect 288710 282820 288716 282832
rect 288768 282820 288774 282872
rect 229370 282752 229376 282804
rect 229428 282752 229434 282804
rect 298480 282792 298508 282888
rect 298554 282792 298560 282804
rect 298480 282764 298560 282792
rect 298554 282752 298560 282764
rect 298612 282752 298618 282804
rect 345198 280276 345204 280288
rect 345159 280248 345204 280276
rect 345198 280236 345204 280248
rect 345256 280236 345262 280288
rect 235074 280208 235080 280220
rect 235035 280180 235080 280208
rect 235074 280168 235080 280180
rect 235132 280168 235138 280220
rect 434254 280208 434260 280220
rect 434215 280180 434260 280208
rect 434254 280168 434260 280180
rect 434312 280168 434318 280220
rect 3142 280100 3148 280152
rect 3200 280140 3206 280152
rect 6270 280140 6276 280152
rect 3200 280112 6276 280140
rect 3200 280100 3206 280112
rect 6270 280100 6276 280112
rect 6328 280100 6334 280152
rect 229370 280140 229376 280152
rect 229331 280112 229376 280140
rect 229370 280100 229376 280112
rect 229428 280100 229434 280152
rect 254210 280140 254216 280152
rect 254171 280112 254216 280140
rect 254210 280100 254216 280112
rect 254268 280100 254274 280152
rect 287330 280140 287336 280152
rect 287291 280112 287336 280140
rect 287330 280100 287336 280112
rect 287388 280100 287394 280152
rect 290090 280140 290096 280152
rect 290051 280112 290096 280140
rect 290090 280100 290096 280112
rect 290148 280100 290154 280152
rect 291470 280100 291476 280152
rect 291528 280140 291534 280152
rect 291562 280140 291568 280152
rect 291528 280112 291568 280140
rect 291528 280100 291534 280112
rect 291562 280100 291568 280112
rect 291620 280100 291626 280152
rect 298465 280143 298523 280149
rect 298465 280109 298477 280143
rect 298511 280140 298523 280143
rect 298554 280140 298560 280152
rect 298511 280112 298560 280140
rect 298511 280109 298523 280112
rect 298465 280103 298523 280109
rect 298554 280100 298560 280112
rect 298612 280100 298618 280152
rect 305454 280140 305460 280152
rect 305288 280112 305460 280140
rect 305288 280084 305316 280112
rect 305454 280100 305460 280112
rect 305512 280100 305518 280152
rect 324498 280100 324504 280152
rect 324556 280140 324562 280152
rect 324774 280140 324780 280152
rect 324556 280112 324780 280140
rect 324556 280100 324562 280112
rect 324774 280100 324780 280112
rect 324832 280100 324838 280152
rect 327534 280140 327540 280152
rect 327368 280112 327540 280140
rect 327368 280084 327396 280112
rect 327534 280100 327540 280112
rect 327592 280100 327598 280152
rect 342530 280140 342536 280152
rect 342491 280112 342536 280140
rect 342530 280100 342536 280112
rect 342588 280100 342594 280152
rect 347958 280100 347964 280152
rect 348016 280140 348022 280152
rect 348050 280140 348056 280152
rect 348016 280112 348056 280140
rect 348016 280100 348022 280112
rect 348050 280100 348056 280112
rect 348108 280100 348114 280152
rect 363138 280140 363144 280152
rect 363099 280112 363144 280140
rect 363138 280100 363144 280112
rect 363196 280100 363202 280152
rect 305270 280032 305276 280084
rect 305328 280032 305334 280084
rect 327350 280032 327356 280084
rect 327408 280032 327414 280084
rect 262398 278916 262404 278928
rect 262324 278888 262404 278916
rect 239122 278740 239128 278792
rect 239180 278780 239186 278792
rect 239306 278780 239312 278792
rect 239180 278752 239312 278780
rect 239180 278740 239186 278752
rect 239306 278740 239312 278752
rect 239364 278740 239370 278792
rect 251174 278740 251180 278792
rect 251232 278780 251238 278792
rect 251450 278780 251456 278792
rect 251232 278752 251456 278780
rect 251232 278740 251238 278752
rect 251450 278740 251456 278752
rect 251508 278740 251514 278792
rect 255498 278740 255504 278792
rect 255556 278780 255562 278792
rect 255866 278780 255872 278792
rect 255556 278752 255872 278780
rect 255556 278740 255562 278752
rect 255866 278740 255872 278752
rect 255924 278740 255930 278792
rect 262324 278780 262352 278888
rect 262398 278876 262404 278888
rect 262456 278876 262462 278928
rect 262490 278848 262496 278860
rect 262451 278820 262496 278848
rect 262490 278808 262496 278820
rect 262548 278808 262554 278860
rect 262398 278780 262404 278792
rect 262324 278752 262404 278780
rect 262398 278740 262404 278752
rect 262456 278740 262462 278792
rect 307938 278740 307944 278792
rect 307996 278780 308002 278792
rect 308214 278780 308220 278792
rect 307996 278752 308220 278780
rect 307996 278740 308002 278752
rect 308214 278740 308220 278752
rect 308272 278740 308278 278792
rect 316218 278740 316224 278792
rect 316276 278780 316282 278792
rect 316310 278780 316316 278792
rect 316276 278752 316316 278780
rect 316276 278740 316282 278752
rect 316310 278740 316316 278752
rect 316368 278740 316374 278792
rect 235074 278712 235080 278724
rect 235035 278684 235080 278712
rect 235074 278672 235080 278684
rect 235132 278672 235138 278724
rect 262490 278712 262496 278724
rect 262451 278684 262496 278712
rect 262490 278672 262496 278684
rect 262548 278672 262554 278724
rect 324498 278712 324504 278724
rect 324459 278684 324504 278712
rect 324498 278672 324504 278684
rect 324556 278672 324562 278724
rect 435358 278060 435364 278112
rect 435416 278100 435422 278112
rect 435542 278100 435548 278112
rect 435416 278072 435548 278100
rect 435416 278060 435422 278072
rect 435542 278060 435548 278072
rect 435600 278060 435606 278112
rect 310698 277380 310704 277432
rect 310756 277420 310762 277432
rect 310790 277420 310796 277432
rect 310756 277392 310796 277420
rect 310756 277380 310762 277392
rect 310790 277380 310796 277392
rect 310848 277380 310854 277432
rect 239122 274048 239128 274100
rect 239180 274088 239186 274100
rect 239309 274091 239367 274097
rect 239309 274088 239321 274091
rect 239180 274060 239321 274088
rect 239180 274048 239186 274060
rect 239309 274057 239321 274060
rect 239355 274057 239367 274091
rect 239309 274051 239367 274057
rect 251450 273884 251456 273896
rect 251411 273856 251456 273884
rect 251450 273844 251456 273856
rect 251508 273844 251514 273896
rect 310698 273408 310704 273420
rect 310659 273380 310704 273408
rect 310698 273368 310704 273380
rect 310756 273368 310762 273420
rect 261202 273164 261208 273216
rect 261260 273164 261266 273216
rect 299842 273164 299848 273216
rect 299900 273164 299906 273216
rect 309410 273204 309416 273216
rect 309371 273176 309416 273204
rect 309410 273164 309416 273176
rect 309468 273164 309474 273216
rect 325970 273164 325976 273216
rect 326028 273164 326034 273216
rect 229370 273136 229376 273148
rect 229331 273108 229376 273136
rect 229370 273096 229376 273108
rect 229428 273096 229434 273148
rect 261220 273080 261248 273164
rect 299860 273080 299888 273164
rect 325988 273080 326016 273164
rect 261202 273028 261208 273080
rect 261260 273028 261266 273080
rect 299842 273028 299848 273080
rect 299900 273028 299906 273080
rect 325970 273028 325976 273080
rect 326028 273028 326034 273080
rect 290090 273000 290096 273012
rect 290051 272972 290096 273000
rect 290090 272960 290096 272972
rect 290148 272960 290154 273012
rect 298462 270620 298468 270632
rect 298423 270592 298468 270620
rect 298462 270580 298468 270592
rect 298520 270580 298526 270632
rect 254210 270552 254216 270564
rect 254171 270524 254216 270552
rect 254210 270512 254216 270524
rect 254268 270512 254274 270564
rect 255590 270512 255596 270564
rect 255648 270552 255654 270564
rect 255866 270552 255872 270564
rect 255648 270524 255872 270552
rect 255648 270512 255654 270524
rect 255866 270512 255872 270524
rect 255924 270512 255930 270564
rect 287330 270552 287336 270564
rect 287291 270524 287336 270552
rect 287330 270512 287336 270524
rect 287388 270512 287394 270564
rect 288618 270512 288624 270564
rect 288676 270552 288682 270564
rect 288710 270552 288716 270564
rect 288676 270524 288716 270552
rect 288676 270512 288682 270524
rect 288710 270512 288716 270524
rect 288768 270512 288774 270564
rect 342530 270552 342536 270564
rect 342491 270524 342536 270552
rect 342530 270512 342536 270524
rect 342588 270512 342594 270564
rect 363141 270555 363199 270561
rect 363141 270521 363153 270555
rect 363187 270552 363199 270555
rect 363230 270552 363236 270564
rect 363187 270524 363236 270552
rect 363187 270521 363199 270524
rect 363141 270515 363199 270521
rect 363230 270512 363236 270524
rect 363288 270512 363294 270564
rect 229370 270484 229376 270496
rect 229331 270456 229376 270484
rect 229370 270444 229376 270456
rect 229428 270444 229434 270496
rect 244274 270484 244280 270496
rect 244235 270456 244280 270484
rect 244274 270444 244280 270456
rect 244332 270444 244338 270496
rect 245930 270484 245936 270496
rect 245891 270456 245936 270484
rect 245930 270444 245936 270456
rect 245988 270444 245994 270496
rect 307938 270484 307944 270496
rect 307899 270456 307944 270484
rect 307938 270444 307944 270456
rect 307996 270444 308002 270496
rect 345198 270484 345204 270496
rect 345159 270456 345204 270484
rect 345198 270444 345204 270456
rect 345256 270444 345262 270496
rect 347958 270484 347964 270496
rect 347919 270456 347964 270484
rect 347958 270444 347964 270456
rect 348016 270444 348022 270496
rect 434257 270487 434315 270493
rect 434257 270453 434269 270487
rect 434303 270484 434315 270487
rect 434346 270484 434352 270496
rect 434303 270456 434352 270484
rect 434303 270453 434315 270456
rect 434257 270447 434315 270453
rect 434346 270444 434352 270456
rect 434404 270444 434410 270496
rect 255590 270416 255596 270428
rect 255551 270388 255596 270416
rect 255590 270376 255596 270388
rect 255648 270376 255654 270428
rect 288710 270416 288716 270428
rect 288671 270388 288716 270416
rect 288710 270376 288716 270388
rect 288768 270376 288774 270428
rect 240226 269084 240232 269136
rect 240284 269124 240290 269136
rect 240410 269124 240416 269136
rect 240284 269096 240416 269124
rect 240284 269084 240290 269096
rect 240410 269084 240416 269096
rect 240468 269084 240474 269136
rect 241882 269084 241888 269136
rect 241940 269124 241946 269136
rect 242066 269124 242072 269136
rect 241940 269096 242072 269124
rect 241940 269084 241946 269096
rect 242066 269084 242072 269096
rect 242124 269084 242130 269136
rect 291470 269084 291476 269136
rect 291528 269124 291534 269136
rect 291654 269124 291660 269136
rect 291528 269096 291660 269124
rect 291528 269084 291534 269096
rect 291654 269084 291660 269096
rect 291712 269084 291718 269136
rect 310701 267835 310759 267841
rect 310701 267801 310713 267835
rect 310747 267832 310759 267835
rect 310790 267832 310796 267844
rect 310747 267804 310796 267832
rect 310747 267801 310759 267804
rect 310701 267795 310759 267801
rect 310790 267792 310796 267804
rect 310848 267792 310854 267844
rect 239306 267724 239312 267776
rect 239364 267764 239370 267776
rect 309410 267764 309416 267776
rect 239364 267736 239409 267764
rect 309371 267736 309416 267764
rect 239364 267724 239370 267736
rect 309410 267724 309416 267736
rect 309468 267724 309474 267776
rect 310790 263644 310796 263696
rect 310848 263644 310854 263696
rect 233326 263576 233332 263628
rect 233384 263616 233390 263628
rect 233510 263616 233516 263628
rect 233384 263588 233516 263616
rect 233384 263576 233390 263588
rect 233510 263576 233516 263588
rect 233568 263576 233574 263628
rect 280430 263576 280436 263628
rect 280488 263616 280494 263628
rect 280614 263616 280620 263628
rect 280488 263588 280620 263616
rect 280488 263576 280494 263588
rect 280614 263576 280620 263588
rect 280672 263576 280678 263628
rect 291470 263576 291476 263628
rect 291528 263576 291534 263628
rect 298462 263576 298468 263628
rect 298520 263576 298526 263628
rect 288710 263548 288716 263560
rect 288671 263520 288716 263548
rect 288710 263508 288716 263520
rect 288768 263508 288774 263560
rect 229370 263480 229376 263492
rect 229331 263452 229376 263480
rect 229370 263440 229376 263452
rect 229428 263440 229434 263492
rect 262493 263483 262551 263489
rect 262493 263449 262505 263483
rect 262539 263480 262551 263483
rect 262674 263480 262680 263492
rect 262539 263452 262680 263480
rect 262539 263449 262551 263452
rect 262493 263443 262551 263449
rect 262674 263440 262680 263452
rect 262732 263440 262738 263492
rect 291488 263480 291516 263576
rect 291562 263480 291568 263492
rect 291488 263452 291568 263480
rect 291562 263440 291568 263452
rect 291620 263440 291626 263492
rect 298480 263480 298508 263576
rect 310808 263560 310836 263644
rect 435358 263576 435364 263628
rect 435416 263616 435422 263628
rect 435542 263616 435548 263628
rect 435416 263588 435548 263616
rect 435416 263576 435422 263588
rect 435542 263576 435548 263588
rect 435600 263576 435606 263628
rect 444006 263576 444012 263628
rect 444064 263616 444070 263628
rect 444190 263616 444196 263628
rect 444064 263588 444196 263616
rect 444064 263576 444070 263588
rect 444190 263576 444196 263588
rect 444248 263576 444254 263628
rect 310790 263508 310796 263560
rect 310848 263508 310854 263560
rect 298554 263480 298560 263492
rect 298480 263452 298560 263480
rect 298554 263440 298560 263452
rect 298612 263440 298618 263492
rect 324501 263483 324559 263489
rect 324501 263449 324513 263483
rect 324547 263480 324559 263483
rect 324682 263480 324688 263492
rect 324547 263452 324688 263480
rect 324547 263449 324559 263452
rect 324501 263443 324559 263449
rect 324682 263440 324688 263452
rect 324740 263440 324746 263492
rect 345198 260964 345204 260976
rect 345159 260936 345204 260964
rect 345198 260924 345204 260936
rect 345256 260924 345262 260976
rect 347958 260964 347964 260976
rect 347919 260936 347964 260964
rect 347958 260924 347964 260936
rect 348016 260924 348022 260976
rect 235074 260896 235080 260908
rect 235035 260868 235080 260896
rect 235074 260856 235080 260868
rect 235132 260856 235138 260908
rect 244274 260896 244280 260908
rect 244235 260868 244280 260896
rect 244274 260856 244280 260868
rect 244332 260856 244338 260908
rect 245930 260896 245936 260908
rect 245891 260868 245936 260896
rect 245930 260856 245936 260868
rect 245988 260856 245994 260908
rect 251450 260896 251456 260908
rect 251411 260868 251456 260896
rect 251450 260856 251456 260868
rect 251508 260856 251514 260908
rect 255593 260899 255651 260905
rect 255593 260865 255605 260899
rect 255639 260896 255651 260899
rect 255682 260896 255688 260908
rect 255639 260868 255688 260896
rect 255639 260865 255651 260868
rect 255593 260859 255651 260865
rect 255682 260856 255688 260868
rect 255740 260856 255746 260908
rect 434254 260896 434260 260908
rect 434215 260868 434260 260896
rect 434254 260856 434260 260868
rect 434312 260856 434318 260908
rect 229370 260828 229376 260840
rect 229331 260800 229376 260828
rect 229370 260788 229376 260800
rect 229428 260788 229434 260840
rect 254210 260828 254216 260840
rect 254171 260800 254216 260828
rect 254210 260788 254216 260800
rect 254268 260788 254274 260840
rect 262585 260831 262643 260837
rect 262585 260797 262597 260831
rect 262631 260828 262643 260831
rect 262674 260828 262680 260840
rect 262631 260800 262680 260828
rect 262631 260797 262643 260800
rect 262585 260791 262643 260797
rect 262674 260788 262680 260800
rect 262732 260788 262738 260840
rect 287330 260828 287336 260840
rect 287291 260800 287336 260828
rect 287330 260788 287336 260800
rect 287388 260788 287394 260840
rect 290090 260828 290096 260840
rect 290051 260800 290096 260828
rect 290090 260788 290096 260800
rect 290148 260788 290154 260840
rect 291473 260831 291531 260837
rect 291473 260797 291485 260831
rect 291519 260828 291531 260831
rect 291562 260828 291568 260840
rect 291519 260800 291568 260828
rect 291519 260797 291531 260800
rect 291473 260791 291531 260797
rect 291562 260788 291568 260800
rect 291620 260788 291626 260840
rect 298465 260831 298523 260837
rect 298465 260797 298477 260831
rect 298511 260828 298523 260831
rect 298554 260828 298560 260840
rect 298511 260800 298560 260828
rect 298511 260797 298523 260800
rect 298465 260791 298523 260797
rect 298554 260788 298560 260800
rect 298612 260788 298618 260840
rect 324593 260831 324651 260837
rect 324593 260797 324605 260831
rect 324639 260828 324651 260831
rect 324682 260828 324688 260840
rect 324639 260800 324688 260828
rect 324639 260797 324651 260800
rect 324593 260791 324651 260797
rect 324682 260788 324688 260800
rect 324740 260788 324746 260840
rect 342530 260828 342536 260840
rect 342491 260800 342536 260828
rect 342530 260788 342536 260800
rect 342588 260788 342594 260840
rect 347958 260788 347964 260840
rect 348016 260828 348022 260840
rect 363138 260828 363144 260840
rect 348016 260800 348096 260828
rect 363099 260800 363144 260828
rect 348016 260788 348022 260800
rect 348068 260772 348096 260800
rect 363138 260788 363144 260800
rect 363196 260788 363202 260840
rect 435266 260828 435272 260840
rect 435227 260800 435272 260828
rect 435266 260788 435272 260800
rect 435324 260788 435330 260840
rect 255593 260763 255651 260769
rect 255593 260729 255605 260763
rect 255639 260760 255651 260763
rect 255682 260760 255688 260772
rect 255639 260732 255688 260760
rect 255639 260729 255651 260732
rect 255593 260723 255651 260729
rect 255682 260720 255688 260732
rect 255740 260720 255746 260772
rect 348050 260720 348056 260772
rect 348108 260720 348114 260772
rect 234614 259428 234620 259480
rect 234672 259468 234678 259480
rect 234890 259468 234896 259480
rect 234672 259440 234896 259468
rect 234672 259428 234678 259440
rect 234890 259428 234896 259440
rect 234948 259428 234954 259480
rect 239122 259428 239128 259480
rect 239180 259468 239186 259480
rect 239306 259468 239312 259480
rect 239180 259440 239312 259468
rect 239180 259428 239186 259440
rect 239306 259428 239312 259440
rect 239364 259428 239370 259480
rect 267182 259428 267188 259480
rect 267240 259468 267246 259480
rect 267274 259468 267280 259480
rect 267240 259440 267280 259468
rect 267240 259428 267246 259440
rect 267274 259428 267280 259440
rect 267332 259428 267338 259480
rect 235074 259400 235080 259412
rect 235035 259372 235080 259400
rect 235074 259360 235080 259372
rect 235132 259360 235138 259412
rect 251450 259400 251456 259412
rect 251411 259372 251456 259400
rect 251450 259360 251456 259372
rect 251508 259360 251514 259412
rect 307938 258108 307944 258120
rect 307899 258080 307944 258108
rect 307938 258068 307944 258080
rect 307996 258068 308002 258120
rect 310793 256683 310851 256689
rect 310793 256649 310805 256683
rect 310839 256680 310851 256683
rect 310882 256680 310888 256692
rect 310839 256652 310888 256680
rect 310839 256649 310851 256652
rect 310793 256643 310851 256649
rect 310882 256640 310888 256652
rect 310940 256640 310946 256692
rect 261202 253852 261208 253904
rect 261260 253852 261266 253904
rect 299842 253852 299848 253904
rect 299900 253852 299906 253904
rect 325970 253852 325976 253904
rect 326028 253852 326034 253904
rect 229370 253824 229376 253836
rect 229331 253796 229376 253824
rect 229370 253784 229376 253796
rect 229428 253784 229434 253836
rect 261220 253768 261248 253852
rect 299860 253768 299888 253852
rect 325988 253768 326016 253852
rect 261202 253716 261208 253768
rect 261260 253716 261266 253768
rect 299842 253716 299848 253768
rect 299900 253716 299906 253768
rect 325970 253716 325976 253768
rect 326028 253716 326034 253768
rect 290090 252872 290096 252884
rect 290051 252844 290096 252872
rect 290090 252832 290096 252844
rect 290148 252832 290154 252884
rect 291470 251308 291476 251320
rect 291431 251280 291476 251308
rect 291470 251268 291476 251280
rect 291528 251268 291534 251320
rect 298462 251308 298468 251320
rect 298423 251280 298468 251308
rect 298462 251268 298468 251280
rect 298520 251268 298526 251320
rect 435266 251308 435272 251320
rect 435227 251280 435272 251308
rect 435266 251268 435272 251280
rect 435324 251268 435330 251320
rect 234890 251200 234896 251252
rect 234948 251200 234954 251252
rect 254210 251240 254216 251252
rect 254171 251212 254216 251240
rect 254210 251200 254216 251212
rect 254268 251200 254274 251252
rect 255590 251240 255596 251252
rect 255551 251212 255596 251240
rect 255590 251200 255596 251212
rect 255648 251200 255654 251252
rect 262582 251240 262588 251252
rect 262543 251212 262588 251240
rect 262582 251200 262588 251212
rect 262640 251200 262646 251252
rect 287330 251240 287336 251252
rect 287291 251212 287336 251240
rect 287330 251200 287336 251212
rect 287388 251200 287394 251252
rect 288618 251200 288624 251252
rect 288676 251240 288682 251252
rect 288710 251240 288716 251252
rect 288676 251212 288716 251240
rect 288676 251200 288682 251212
rect 288710 251200 288716 251212
rect 288768 251200 288774 251252
rect 324590 251240 324596 251252
rect 324551 251212 324596 251240
rect 324590 251200 324596 251212
rect 324648 251200 324654 251252
rect 342530 251240 342536 251252
rect 342491 251212 342536 251240
rect 342530 251200 342536 251212
rect 342588 251200 342594 251252
rect 363141 251243 363199 251249
rect 363141 251209 363153 251243
rect 363187 251240 363199 251243
rect 363230 251240 363236 251252
rect 363187 251212 363236 251240
rect 363187 251209 363199 251212
rect 363141 251203 363199 251209
rect 363230 251200 363236 251212
rect 363288 251200 363294 251252
rect 234908 251104 234936 251200
rect 244274 251172 244280 251184
rect 244235 251144 244280 251172
rect 244274 251132 244280 251144
rect 244332 251132 244338 251184
rect 245930 251172 245936 251184
rect 245891 251144 245936 251172
rect 245930 251132 245936 251144
rect 245988 251132 245994 251184
rect 291470 251172 291476 251184
rect 291431 251144 291476 251172
rect 291470 251132 291476 251144
rect 291528 251132 291534 251184
rect 298462 251172 298468 251184
rect 298423 251144 298468 251172
rect 298462 251132 298468 251144
rect 298520 251132 298526 251184
rect 305181 251175 305239 251181
rect 305181 251141 305193 251175
rect 305227 251172 305239 251175
rect 305270 251172 305276 251184
rect 305227 251144 305276 251172
rect 305227 251141 305239 251144
rect 305181 251135 305239 251141
rect 305270 251132 305276 251144
rect 305328 251132 305334 251184
rect 307938 251172 307944 251184
rect 307899 251144 307944 251172
rect 307938 251132 307944 251144
rect 307996 251132 308002 251184
rect 327261 251175 327319 251181
rect 327261 251141 327273 251175
rect 327307 251172 327319 251175
rect 327350 251172 327356 251184
rect 327307 251144 327356 251172
rect 327307 251141 327319 251144
rect 327261 251135 327319 251141
rect 327350 251132 327356 251144
rect 327408 251132 327414 251184
rect 345198 251172 345204 251184
rect 345159 251144 345204 251172
rect 345198 251132 345204 251144
rect 345256 251132 345262 251184
rect 347958 251172 347964 251184
rect 347919 251144 347964 251172
rect 347958 251132 347964 251144
rect 348016 251132 348022 251184
rect 434257 251175 434315 251181
rect 434257 251141 434269 251175
rect 434303 251172 434315 251175
rect 434346 251172 434352 251184
rect 434303 251144 434352 251172
rect 434303 251141 434315 251144
rect 434257 251135 434315 251141
rect 434346 251132 434352 251144
rect 434404 251132 434410 251184
rect 435085 251175 435143 251181
rect 435085 251141 435097 251175
rect 435131 251172 435143 251175
rect 435174 251172 435180 251184
rect 435131 251144 435180 251172
rect 435131 251141 435143 251144
rect 435085 251135 435143 251141
rect 435174 251132 435180 251144
rect 435232 251132 435238 251184
rect 234982 251104 234988 251116
rect 234908 251076 234988 251104
rect 234982 251064 234988 251076
rect 235040 251064 235046 251116
rect 251453 251107 251511 251113
rect 251453 251073 251465 251107
rect 251499 251104 251511 251107
rect 251542 251104 251548 251116
rect 251499 251076 251548 251104
rect 251499 251073 251511 251076
rect 251453 251067 251511 251073
rect 251542 251064 251548 251076
rect 251600 251064 251606 251116
rect 239125 249883 239183 249889
rect 239125 249849 239137 249883
rect 239171 249880 239183 249883
rect 239214 249880 239220 249892
rect 239171 249852 239220 249880
rect 239171 249849 239183 249852
rect 239125 249843 239183 249849
rect 239214 249840 239220 249852
rect 239272 249840 239278 249892
rect 240226 249772 240232 249824
rect 240284 249812 240290 249824
rect 240410 249812 240416 249824
rect 240284 249784 240416 249812
rect 240284 249772 240290 249784
rect 240410 249772 240416 249784
rect 240468 249772 240474 249824
rect 241882 249772 241888 249824
rect 241940 249812 241946 249824
rect 242066 249812 242072 249824
rect 241940 249784 242072 249812
rect 241940 249772 241946 249784
rect 242066 249772 242072 249784
rect 242124 249772 242130 249824
rect 266998 249772 267004 249824
rect 267056 249812 267062 249824
rect 267274 249812 267280 249824
rect 267056 249784 267280 249812
rect 267056 249772 267062 249784
rect 267274 249772 267280 249784
rect 267332 249772 267338 249824
rect 229370 244372 229376 244384
rect 229296 244344 229376 244372
rect 229296 244248 229324 244344
rect 229370 244332 229376 244344
rect 229428 244332 229434 244384
rect 233326 244264 233332 244316
rect 233384 244304 233390 244316
rect 233510 244304 233516 244316
rect 233384 244276 233516 244304
rect 233384 244264 233390 244276
rect 233510 244264 233516 244276
rect 233568 244264 233574 244316
rect 288710 244264 288716 244316
rect 288768 244264 288774 244316
rect 444006 244264 444012 244316
rect 444064 244304 444070 244316
rect 444190 244304 444196 244316
rect 444064 244276 444196 244304
rect 444064 244264 444070 244276
rect 444190 244264 444196 244276
rect 444248 244264 444254 244316
rect 229278 244196 229284 244248
rect 229336 244196 229342 244248
rect 288728 244168 288756 244264
rect 307941 244239 307999 244245
rect 307941 244205 307953 244239
rect 307987 244236 307999 244239
rect 308030 244236 308036 244248
rect 307987 244208 308036 244236
rect 307987 244205 307999 244208
rect 307941 244199 307999 244205
rect 308030 244196 308036 244208
rect 308088 244196 308094 244248
rect 288802 244168 288808 244180
rect 288728 244140 288808 244168
rect 288802 244128 288808 244140
rect 288860 244128 288866 244180
rect 327258 242672 327264 242684
rect 327219 242644 327264 242672
rect 327258 242632 327264 242644
rect 327316 242632 327322 242684
rect 234890 241476 234896 241528
rect 234948 241516 234954 241528
rect 234982 241516 234988 241528
rect 234948 241488 234988 241516
rect 234948 241476 234954 241488
rect 234982 241476 234988 241488
rect 235040 241476 235046 241528
rect 235074 241476 235080 241528
rect 235132 241516 235138 241528
rect 244274 241516 244280 241528
rect 235132 241488 235177 241516
rect 244235 241488 244280 241516
rect 235132 241476 235138 241488
rect 244274 241476 244280 241488
rect 244332 241476 244338 241528
rect 245930 241516 245936 241528
rect 245891 241488 245936 241516
rect 245930 241476 245936 241488
rect 245988 241476 245994 241528
rect 251450 241516 251456 241528
rect 251411 241488 251456 241516
rect 251450 241476 251456 241488
rect 251508 241476 251514 241528
rect 255774 241476 255780 241528
rect 255832 241516 255838 241528
rect 255866 241516 255872 241528
rect 255832 241488 255872 241516
rect 255832 241476 255838 241488
rect 255866 241476 255872 241488
rect 255924 241476 255930 241528
rect 262766 241476 262772 241528
rect 262824 241516 262830 241528
rect 262858 241516 262864 241528
rect 262824 241488 262864 241516
rect 262824 241476 262830 241488
rect 262858 241476 262864 241488
rect 262916 241476 262922 241528
rect 266998 241476 267004 241528
rect 267056 241476 267062 241528
rect 291473 241519 291531 241525
rect 291473 241485 291485 241519
rect 291519 241516 291531 241519
rect 291562 241516 291568 241528
rect 291519 241488 291568 241516
rect 291519 241485 291531 241488
rect 291473 241479 291531 241485
rect 291562 241476 291568 241488
rect 291620 241476 291626 241528
rect 298465 241519 298523 241525
rect 298465 241485 298477 241519
rect 298511 241516 298523 241519
rect 298554 241516 298560 241528
rect 298511 241488 298560 241516
rect 298511 241485 298523 241488
rect 298465 241479 298523 241485
rect 298554 241476 298560 241488
rect 298612 241476 298618 241528
rect 305178 241516 305184 241528
rect 305139 241488 305184 241516
rect 305178 241476 305184 241488
rect 305236 241476 305242 241528
rect 324774 241476 324780 241528
rect 324832 241516 324838 241528
rect 324866 241516 324872 241528
rect 324832 241488 324872 241516
rect 324832 241476 324838 241488
rect 324866 241476 324872 241488
rect 324924 241476 324930 241528
rect 345198 241516 345204 241528
rect 345159 241488 345204 241516
rect 345198 241476 345204 241488
rect 345256 241476 345262 241528
rect 347958 241516 347964 241528
rect 347919 241488 347964 241516
rect 347958 241476 347964 241488
rect 348016 241476 348022 241528
rect 434254 241516 434260 241528
rect 434215 241488 434260 241516
rect 434254 241476 434260 241488
rect 434312 241476 434318 241528
rect 435082 241516 435088 241528
rect 435043 241488 435088 241516
rect 435082 241476 435088 241488
rect 435140 241476 435146 241528
rect 267016 241392 267044 241476
rect 266998 241340 267004 241392
rect 267056 241340 267062 241392
rect 239122 240156 239128 240168
rect 239083 240128 239128 240156
rect 239122 240116 239128 240128
rect 239180 240116 239186 240168
rect 251450 240156 251456 240168
rect 251411 240128 251456 240156
rect 251450 240116 251456 240128
rect 251508 240116 251514 240168
rect 234890 240088 234896 240100
rect 234851 240060 234896 240088
rect 234890 240048 234896 240060
rect 234948 240048 234954 240100
rect 288710 240088 288716 240100
rect 288671 240060 288716 240088
rect 288710 240048 288716 240060
rect 288768 240048 288774 240100
rect 327258 240048 327264 240100
rect 327316 240088 327322 240100
rect 327350 240088 327356 240100
rect 327316 240060 327356 240088
rect 327316 240048 327322 240060
rect 327350 240048 327356 240060
rect 327408 240048 327414 240100
rect 251450 240020 251456 240032
rect 251411 239992 251456 240020
rect 251450 239980 251456 239992
rect 251508 239980 251514 240032
rect 310790 240020 310796 240032
rect 310751 239992 310796 240020
rect 310790 239980 310796 239992
rect 310848 239980 310854 240032
rect 310698 238688 310704 238740
rect 310756 238728 310762 238740
rect 310790 238728 310796 238740
rect 310756 238700 310796 238728
rect 310756 238688 310762 238700
rect 310790 238688 310796 238700
rect 310848 238688 310854 238740
rect 280614 234716 280620 234728
rect 280540 234688 280620 234716
rect 280540 234592 280568 234688
rect 280614 234676 280620 234688
rect 280672 234676 280678 234728
rect 434254 234608 434260 234660
rect 434312 234608 434318 234660
rect 435082 234608 435088 234660
rect 435140 234608 435146 234660
rect 261202 234540 261208 234592
rect 261260 234540 261266 234592
rect 280522 234540 280528 234592
rect 280580 234540 280586 234592
rect 287330 234540 287336 234592
rect 287388 234540 287394 234592
rect 299842 234540 299848 234592
rect 299900 234540 299906 234592
rect 325970 234540 325976 234592
rect 326028 234540 326034 234592
rect 261220 234456 261248 234540
rect 287348 234456 287376 234540
rect 299860 234456 299888 234540
rect 325988 234456 326016 234540
rect 434272 234512 434300 234608
rect 434346 234512 434352 234524
rect 434272 234484 434352 234512
rect 434346 234472 434352 234484
rect 434404 234472 434410 234524
rect 435100 234512 435128 234608
rect 435174 234512 435180 234524
rect 435100 234484 435180 234512
rect 435174 234472 435180 234484
rect 435232 234472 435238 234524
rect 261202 234404 261208 234456
rect 261260 234404 261266 234456
rect 287330 234404 287336 234456
rect 287388 234404 287394 234456
rect 299842 234404 299848 234456
rect 299900 234404 299906 234456
rect 325970 234404 325976 234456
rect 326028 234404 326034 234456
rect 308030 231956 308036 232008
rect 308088 231956 308094 232008
rect 308048 231872 308076 231956
rect 345382 231888 345388 231940
rect 345440 231888 345446 231940
rect 254210 231820 254216 231872
rect 254268 231860 254274 231872
rect 254394 231860 254400 231872
rect 254268 231832 254400 231860
rect 254268 231820 254274 231832
rect 254394 231820 254400 231832
rect 254452 231820 254458 231872
rect 262582 231820 262588 231872
rect 262640 231860 262646 231872
rect 262858 231860 262864 231872
rect 262640 231832 262864 231860
rect 262640 231820 262646 231832
rect 262858 231820 262864 231832
rect 262916 231820 262922 231872
rect 288713 231863 288771 231869
rect 288713 231829 288725 231863
rect 288759 231860 288771 231863
rect 288802 231860 288808 231872
rect 288759 231832 288808 231860
rect 288759 231829 288771 231832
rect 288713 231823 288771 231829
rect 288802 231820 288808 231832
rect 288860 231820 288866 231872
rect 298554 231820 298560 231872
rect 298612 231820 298618 231872
rect 305178 231820 305184 231872
rect 305236 231860 305242 231872
rect 305270 231860 305276 231872
rect 305236 231832 305276 231860
rect 305236 231820 305242 231832
rect 305270 231820 305276 231832
rect 305328 231820 305334 231872
rect 308030 231820 308036 231872
rect 308088 231820 308094 231872
rect 324590 231820 324596 231872
rect 324648 231860 324654 231872
rect 324866 231860 324872 231872
rect 324648 231832 324872 231860
rect 324648 231820 324654 231832
rect 324866 231820 324872 231832
rect 324924 231820 324930 231872
rect 342346 231820 342352 231872
rect 342404 231860 342410 231872
rect 342530 231860 342536 231872
rect 342404 231832 342536 231860
rect 342404 231820 342410 231832
rect 342530 231820 342536 231832
rect 342588 231820 342594 231872
rect 345290 231820 345296 231872
rect 345348 231860 345354 231872
rect 345400 231860 345428 231888
rect 345348 231832 345428 231860
rect 345348 231820 345354 231832
rect 362954 231820 362960 231872
rect 363012 231860 363018 231872
rect 363230 231860 363236 231872
rect 363012 231832 363236 231860
rect 363012 231820 363018 231832
rect 363230 231820 363236 231832
rect 363288 231820 363294 231872
rect 244458 231752 244464 231804
rect 244516 231792 244522 231804
rect 244550 231792 244556 231804
rect 244516 231764 244556 231792
rect 244516 231752 244522 231764
rect 244550 231752 244556 231764
rect 244608 231752 244614 231804
rect 298572 231736 298600 231820
rect 298554 231684 298560 231736
rect 298612 231684 298618 231736
rect 229370 230460 229376 230512
rect 229428 230500 229434 230512
rect 229554 230500 229560 230512
rect 229428 230472 229560 230500
rect 229428 230460 229434 230472
rect 229554 230460 229560 230472
rect 229612 230460 229618 230512
rect 234890 230500 234896 230512
rect 234851 230472 234896 230500
rect 234890 230460 234896 230472
rect 234948 230460 234954 230512
rect 235074 230460 235080 230512
rect 235132 230500 235138 230512
rect 235258 230500 235264 230512
rect 235132 230472 235264 230500
rect 235132 230460 235138 230472
rect 235258 230460 235264 230472
rect 235316 230460 235322 230512
rect 240226 230460 240232 230512
rect 240284 230500 240290 230512
rect 240410 230500 240416 230512
rect 240284 230472 240416 230500
rect 240284 230460 240290 230472
rect 240410 230460 240416 230472
rect 240468 230460 240474 230512
rect 241882 230460 241888 230512
rect 241940 230500 241946 230512
rect 242066 230500 242072 230512
rect 241940 230472 242072 230500
rect 241940 230460 241946 230472
rect 242066 230460 242072 230472
rect 242124 230460 242130 230512
rect 251450 230500 251456 230512
rect 251411 230472 251456 230500
rect 251450 230460 251456 230472
rect 251508 230460 251514 230512
rect 255774 230460 255780 230512
rect 255832 230500 255838 230512
rect 255866 230500 255872 230512
rect 255832 230472 255872 230500
rect 255832 230460 255838 230472
rect 255866 230460 255872 230472
rect 255924 230460 255930 230512
rect 266814 230460 266820 230512
rect 266872 230500 266878 230512
rect 266998 230500 267004 230512
rect 266872 230472 267004 230500
rect 266872 230460 266878 230472
rect 266998 230460 267004 230472
rect 267056 230460 267062 230512
rect 291562 230460 291568 230512
rect 291620 230500 291626 230512
rect 291654 230500 291660 230512
rect 291620 230472 291660 230500
rect 291620 230460 291626 230472
rect 291654 230460 291660 230472
rect 291712 230460 291718 230512
rect 298554 229032 298560 229084
rect 298612 229072 298618 229084
rect 298646 229072 298652 229084
rect 298612 229044 298652 229072
rect 298612 229032 298618 229044
rect 298646 229032 298652 229044
rect 298704 229032 298710 229084
rect 229370 225060 229376 225072
rect 229296 225032 229376 225060
rect 229296 224936 229324 225032
rect 229370 225020 229376 225032
rect 229428 225020 229434 225072
rect 434346 225060 434352 225072
rect 434272 225032 434352 225060
rect 233326 224952 233332 225004
rect 233384 224992 233390 225004
rect 233510 224992 233516 225004
rect 233384 224964 233516 224992
rect 233384 224952 233390 224964
rect 233510 224952 233516 224964
rect 233568 224952 233574 225004
rect 288802 224952 288808 225004
rect 288860 224952 288866 225004
rect 229278 224884 229284 224936
rect 229336 224884 229342 224936
rect 288820 224868 288848 224952
rect 434272 224936 434300 225032
rect 434346 225020 434352 225032
rect 434404 225020 434410 225072
rect 435082 224992 435088 225004
rect 435043 224964 435088 224992
rect 435082 224952 435088 224964
rect 435140 224952 435146 225004
rect 444006 224952 444012 225004
rect 444064 224992 444070 225004
rect 444190 224992 444196 225004
rect 444064 224964 444196 224992
rect 444064 224952 444070 224964
rect 444190 224952 444196 224964
rect 444248 224952 444254 225004
rect 434254 224884 434260 224936
rect 434312 224884 434318 224936
rect 288802 224816 288808 224868
rect 288860 224816 288866 224868
rect 251174 224204 251180 224256
rect 251232 224244 251238 224256
rect 251450 224244 251456 224256
rect 251232 224216 251456 224244
rect 251232 224204 251238 224216
rect 251450 224204 251456 224216
rect 251508 224204 251514 224256
rect 235074 222300 235080 222352
rect 235132 222300 235138 222352
rect 235092 222216 235120 222300
rect 235074 222164 235080 222216
rect 235132 222164 235138 222216
rect 244182 222164 244188 222216
rect 244240 222204 244246 222216
rect 244274 222204 244280 222216
rect 244240 222176 244280 222204
rect 244240 222164 244246 222176
rect 244274 222164 244280 222176
rect 244332 222164 244338 222216
rect 245746 222164 245752 222216
rect 245804 222204 245810 222216
rect 245930 222204 245936 222216
rect 245804 222176 245936 222204
rect 245804 222164 245810 222176
rect 245930 222164 245936 222176
rect 245988 222164 245994 222216
rect 262490 222164 262496 222216
rect 262548 222204 262554 222216
rect 262858 222204 262864 222216
rect 262548 222176 262864 222204
rect 262548 222164 262554 222176
rect 262858 222164 262864 222176
rect 262916 222164 262922 222216
rect 345198 222164 345204 222216
rect 345256 222204 345262 222216
rect 345290 222204 345296 222216
rect 345256 222176 345296 222204
rect 345256 222164 345262 222176
rect 345290 222164 345296 222176
rect 345348 222164 345354 222216
rect 347958 222164 347964 222216
rect 348016 222204 348022 222216
rect 348142 222204 348148 222216
rect 348016 222176 348148 222204
rect 348016 222164 348022 222176
rect 348142 222164 348148 222176
rect 348200 222164 348206 222216
rect 435082 222204 435088 222216
rect 435043 222176 435088 222204
rect 435082 222164 435088 222176
rect 435140 222164 435146 222216
rect 291378 220872 291384 220924
rect 291436 220912 291442 220924
rect 291746 220912 291752 220924
rect 291436 220884 291752 220912
rect 291436 220872 291442 220884
rect 291746 220872 291752 220884
rect 291804 220872 291810 220924
rect 239122 220804 239128 220856
rect 239180 220844 239186 220856
rect 239214 220844 239220 220856
rect 239180 220816 239220 220844
rect 239180 220804 239186 220816
rect 239214 220804 239220 220816
rect 239272 220804 239278 220856
rect 266906 220804 266912 220856
rect 266964 220844 266970 220856
rect 266998 220844 267004 220856
rect 266964 220816 267004 220844
rect 266964 220804 266970 220816
rect 266998 220804 267004 220816
rect 267056 220804 267062 220856
rect 316218 220804 316224 220856
rect 316276 220844 316282 220856
rect 316310 220844 316316 220856
rect 316276 220816 316316 220844
rect 316276 220804 316282 220816
rect 316310 220804 316316 220816
rect 316368 220804 316374 220856
rect 327350 220804 327356 220856
rect 327408 220844 327414 220856
rect 327534 220844 327540 220856
rect 327408 220816 327540 220844
rect 327408 220804 327414 220816
rect 327534 220804 327540 220816
rect 327592 220804 327598 220856
rect 229278 220776 229284 220788
rect 229239 220748 229284 220776
rect 229278 220736 229284 220748
rect 229336 220736 229342 220788
rect 235074 220776 235080 220788
rect 235035 220748 235080 220776
rect 235074 220736 235080 220748
rect 235132 220736 235138 220788
rect 291378 220776 291384 220788
rect 291339 220748 291384 220776
rect 291378 220736 291384 220748
rect 291436 220736 291442 220788
rect 434254 220776 434260 220788
rect 434215 220748 434260 220776
rect 434254 220736 434260 220748
rect 434312 220736 434318 220788
rect 310882 219416 310888 219428
rect 310843 219388 310888 219416
rect 310882 219376 310888 219388
rect 310940 219376 310946 219428
rect 308030 217444 308036 217456
rect 307991 217416 308036 217444
rect 308030 217404 308036 217416
rect 308088 217404 308094 217456
rect 261202 215976 261208 216028
rect 261260 216016 261266 216028
rect 261386 216016 261392 216028
rect 261260 215988 261392 216016
rect 261260 215976 261266 215988
rect 261386 215976 261392 215988
rect 261444 215976 261450 216028
rect 327350 215364 327356 215416
rect 327408 215364 327414 215416
rect 266998 215336 267004 215348
rect 266959 215308 267004 215336
rect 266998 215296 267004 215308
rect 267056 215296 267062 215348
rect 288710 215336 288716 215348
rect 288671 215308 288716 215336
rect 288710 215296 288716 215308
rect 288768 215296 288774 215348
rect 305362 215336 305368 215348
rect 305288 215308 305368 215336
rect 305288 215280 305316 215308
rect 305362 215296 305368 215308
rect 305420 215296 305426 215348
rect 327368 215280 327396 215364
rect 435082 215296 435088 215348
rect 435140 215296 435146 215348
rect 229278 215268 229284 215280
rect 229239 215240 229284 215268
rect 229278 215228 229284 215240
rect 229336 215228 229342 215280
rect 273346 215228 273352 215280
rect 273404 215268 273410 215280
rect 273530 215268 273536 215280
rect 273404 215240 273536 215268
rect 273404 215228 273410 215240
rect 273530 215228 273536 215240
rect 273588 215228 273594 215280
rect 299842 215228 299848 215280
rect 299900 215228 299906 215280
rect 305270 215228 305276 215280
rect 305328 215228 305334 215280
rect 325970 215228 325976 215280
rect 326028 215228 326034 215280
rect 327350 215228 327356 215280
rect 327408 215228 327414 215280
rect 434254 215268 434260 215280
rect 434215 215240 434260 215268
rect 434254 215228 434260 215240
rect 434312 215228 434318 215280
rect 299860 215144 299888 215228
rect 325988 215144 326016 215228
rect 435100 215200 435128 215296
rect 435174 215200 435180 215212
rect 435100 215172 435180 215200
rect 435174 215160 435180 215172
rect 435232 215160 435238 215212
rect 299842 215092 299848 215144
rect 299900 215092 299906 215144
rect 325970 215092 325976 215144
rect 326028 215092 326034 215144
rect 310882 214588 310888 214600
rect 310843 214560 310888 214588
rect 310882 214548 310888 214560
rect 310940 214548 310946 214600
rect 345382 212576 345388 212628
rect 345440 212576 345446 212628
rect 254210 212508 254216 212560
rect 254268 212548 254274 212560
rect 254394 212548 254400 212560
rect 254268 212520 254400 212548
rect 254268 212508 254274 212520
rect 254394 212508 254400 212520
rect 254452 212508 254458 212560
rect 262582 212508 262588 212560
rect 262640 212548 262646 212560
rect 262858 212548 262864 212560
rect 262640 212520 262864 212548
rect 262640 212508 262646 212520
rect 262858 212508 262864 212520
rect 262916 212508 262922 212560
rect 266998 212548 267004 212560
rect 266959 212520 267004 212548
rect 266998 212508 267004 212520
rect 267056 212508 267062 212560
rect 287330 212508 287336 212560
rect 287388 212548 287394 212560
rect 287514 212548 287520 212560
rect 287388 212520 287520 212548
rect 287388 212508 287394 212520
rect 287514 212508 287520 212520
rect 287572 212508 287578 212560
rect 288713 212551 288771 212557
rect 288713 212517 288725 212551
rect 288759 212548 288771 212551
rect 288802 212548 288808 212560
rect 288759 212520 288808 212548
rect 288759 212517 288771 212520
rect 288713 212511 288771 212517
rect 288802 212508 288808 212520
rect 288860 212508 288866 212560
rect 308030 212548 308036 212560
rect 307991 212520 308036 212548
rect 308030 212508 308036 212520
rect 308088 212508 308094 212560
rect 324590 212508 324596 212560
rect 324648 212548 324654 212560
rect 324866 212548 324872 212560
rect 324648 212520 324872 212548
rect 324648 212508 324654 212520
rect 324866 212508 324872 212520
rect 324924 212508 324930 212560
rect 342346 212508 342352 212560
rect 342404 212548 342410 212560
rect 342530 212548 342536 212560
rect 342404 212520 342536 212548
rect 342404 212508 342410 212520
rect 342530 212508 342536 212520
rect 342588 212508 342594 212560
rect 343818 212548 343824 212560
rect 343744 212520 343824 212548
rect 343744 212492 343772 212520
rect 343818 212508 343824 212520
rect 343876 212508 343882 212560
rect 345290 212508 345296 212560
rect 345348 212548 345354 212560
rect 345400 212548 345428 212576
rect 345348 212520 345428 212548
rect 345348 212508 345354 212520
rect 362954 212508 362960 212560
rect 363012 212548 363018 212560
rect 363230 212548 363236 212560
rect 363012 212520 363236 212548
rect 363012 212508 363018 212520
rect 363230 212508 363236 212520
rect 363288 212508 363294 212560
rect 343726 212440 343732 212492
rect 343784 212440 343790 212492
rect 239030 211216 239036 211268
rect 239088 211256 239094 211268
rect 239122 211256 239128 211268
rect 239088 211228 239128 211256
rect 239088 211216 239094 211228
rect 239122 211216 239128 211228
rect 239180 211216 239186 211268
rect 235074 211188 235080 211200
rect 235035 211160 235080 211188
rect 235074 211148 235080 211160
rect 235132 211148 235138 211200
rect 239122 211120 239128 211132
rect 239083 211092 239128 211120
rect 239122 211080 239128 211092
rect 239180 211080 239186 211132
rect 266998 211120 267004 211132
rect 266959 211092 267004 211120
rect 266998 211080 267004 211092
rect 267056 211080 267062 211132
rect 316310 211080 316316 211132
rect 316368 211120 316374 211132
rect 316494 211120 316500 211132
rect 316368 211092 316500 211120
rect 316368 211080 316374 211092
rect 316494 211080 316500 211092
rect 316552 211080 316558 211132
rect 327350 211080 327356 211132
rect 327408 211120 327414 211132
rect 327534 211120 327540 211132
rect 327408 211092 327540 211120
rect 327408 211080 327414 211092
rect 327534 211080 327540 211092
rect 327592 211080 327598 211132
rect 343726 211120 343732 211132
rect 343687 211092 343732 211120
rect 343726 211080 343732 211092
rect 343784 211080 343790 211132
rect 251358 209720 251364 209772
rect 251416 209760 251422 209772
rect 251726 209760 251732 209772
rect 251416 209732 251732 209760
rect 251416 209720 251422 209732
rect 251726 209720 251732 209732
rect 251784 209720 251790 209772
rect 2774 208156 2780 208208
rect 2832 208196 2838 208208
rect 5166 208196 5172 208208
rect 2832 208168 5172 208196
rect 2832 208156 2838 208168
rect 5166 208156 5172 208168
rect 5224 208156 5230 208208
rect 233326 205640 233332 205692
rect 233384 205680 233390 205692
rect 233510 205680 233516 205692
rect 233384 205652 233516 205680
rect 233384 205640 233390 205652
rect 233510 205640 233516 205652
rect 233568 205640 233574 205692
rect 288802 205680 288808 205692
rect 288763 205652 288808 205680
rect 288802 205640 288808 205652
rect 288860 205640 288866 205692
rect 305270 205680 305276 205692
rect 305231 205652 305276 205680
rect 305270 205640 305276 205652
rect 305328 205640 305334 205692
rect 444006 205640 444012 205692
rect 444064 205680 444070 205692
rect 444190 205680 444196 205692
rect 444064 205652 444196 205680
rect 444064 205640 444070 205652
rect 444190 205640 444196 205652
rect 444248 205640 444254 205692
rect 308030 205504 308036 205556
rect 308088 205544 308094 205556
rect 308214 205544 308220 205556
rect 308088 205516 308220 205544
rect 308088 205504 308094 205516
rect 308214 205504 308220 205516
rect 308272 205504 308278 205556
rect 238754 204552 238760 204604
rect 238812 204592 238818 204604
rect 238938 204592 238944 204604
rect 238812 204564 238944 204592
rect 238812 204552 238818 204564
rect 238938 204552 238944 204564
rect 238996 204552 239002 204604
rect 255590 202920 255596 202972
rect 255648 202960 255654 202972
rect 255682 202960 255688 202972
rect 255648 202932 255688 202960
rect 255648 202920 255654 202932
rect 255682 202920 255688 202932
rect 255740 202920 255746 202972
rect 291378 202960 291384 202972
rect 291339 202932 291384 202960
rect 291378 202920 291384 202932
rect 291436 202920 291442 202972
rect 229278 202852 229284 202904
rect 229336 202892 229342 202904
rect 229370 202892 229376 202904
rect 229336 202864 229376 202892
rect 229336 202852 229342 202864
rect 229370 202852 229376 202864
rect 229428 202852 229434 202904
rect 234798 202852 234804 202904
rect 234856 202892 234862 202904
rect 234890 202892 234896 202904
rect 234856 202864 234896 202892
rect 234856 202852 234862 202864
rect 234890 202852 234896 202864
rect 234948 202852 234954 202904
rect 288802 202892 288808 202904
rect 288763 202864 288808 202892
rect 288802 202852 288808 202864
rect 288860 202852 288866 202904
rect 305270 202892 305276 202904
rect 305231 202864 305276 202892
rect 305270 202852 305276 202864
rect 305328 202852 305334 202904
rect 347958 202852 347964 202904
rect 348016 202892 348022 202904
rect 348142 202892 348148 202904
rect 348016 202864 348148 202892
rect 348016 202852 348022 202864
rect 348142 202852 348148 202864
rect 348200 202852 348206 202904
rect 434346 202852 434352 202904
rect 434404 202892 434410 202904
rect 434530 202892 434536 202904
rect 434404 202864 434536 202892
rect 434404 202852 434410 202864
rect 434530 202852 434536 202864
rect 434588 202852 434594 202904
rect 239122 202824 239128 202836
rect 239083 202796 239128 202824
rect 239122 202784 239128 202796
rect 239180 202784 239186 202836
rect 267001 202827 267059 202833
rect 267001 202793 267013 202827
rect 267047 202824 267059 202827
rect 267090 202824 267096 202836
rect 267047 202796 267096 202824
rect 267047 202793 267059 202796
rect 267001 202787 267059 202793
rect 267090 202784 267096 202796
rect 267148 202784 267154 202836
rect 343726 202824 343732 202836
rect 343687 202796 343732 202824
rect 343726 202784 343732 202796
rect 343784 202784 343790 202836
rect 298554 201492 298560 201544
rect 298612 201532 298618 201544
rect 298646 201532 298652 201544
rect 298612 201504 298652 201532
rect 298612 201492 298618 201504
rect 298646 201492 298652 201504
rect 298704 201492 298710 201544
rect 234798 201464 234804 201476
rect 234759 201436 234804 201464
rect 234798 201424 234804 201436
rect 234856 201424 234862 201476
rect 240410 201464 240416 201476
rect 240371 201436 240416 201464
rect 240410 201424 240416 201436
rect 240468 201424 240474 201476
rect 291378 201424 291384 201476
rect 291436 201464 291442 201476
rect 291654 201464 291660 201476
rect 291436 201436 291660 201464
rect 291436 201424 291442 201436
rect 291654 201424 291660 201436
rect 291712 201424 291718 201476
rect 305270 201464 305276 201476
rect 305231 201436 305276 201464
rect 305270 201424 305276 201436
rect 305328 201424 305334 201476
rect 309318 201424 309324 201476
rect 309376 201424 309382 201476
rect 310790 201424 310796 201476
rect 310848 201464 310854 201476
rect 310882 201464 310888 201476
rect 310848 201436 310888 201464
rect 310848 201424 310854 201436
rect 310882 201424 310888 201436
rect 310940 201424 310946 201476
rect 313550 201424 313556 201476
rect 313608 201464 313614 201476
rect 313642 201464 313648 201476
rect 313608 201436 313648 201464
rect 313608 201424 313614 201436
rect 313642 201424 313648 201436
rect 313700 201424 313706 201476
rect 345017 201467 345075 201473
rect 345017 201433 345029 201467
rect 345063 201464 345075 201467
rect 345198 201464 345204 201476
rect 345063 201436 345204 201464
rect 345063 201433 345075 201436
rect 345017 201427 345075 201433
rect 345198 201424 345204 201436
rect 345256 201424 345262 201476
rect 309336 201396 309364 201424
rect 309410 201396 309416 201408
rect 309336 201368 309416 201396
rect 309410 201356 309416 201368
rect 309468 201356 309474 201408
rect 267001 200107 267059 200113
rect 267001 200073 267013 200107
rect 267047 200104 267059 200107
rect 267090 200104 267096 200116
rect 267047 200076 267096 200104
rect 267047 200073 267059 200076
rect 267001 200067 267059 200073
rect 267090 200064 267096 200076
rect 267148 200064 267154 200116
rect 310790 200104 310796 200116
rect 310751 200076 310796 200104
rect 310790 200064 310796 200076
rect 310848 200064 310854 200116
rect 238846 198472 238852 198484
rect 238807 198444 238852 198472
rect 238846 198432 238852 198444
rect 238904 198432 238910 198484
rect 238846 198064 238852 198076
rect 238807 198036 238852 198064
rect 238846 198024 238852 198036
rect 238904 198024 238910 198076
rect 254210 196596 254216 196648
rect 254268 196636 254274 196648
rect 254394 196636 254400 196648
rect 254268 196608 254400 196636
rect 254268 196596 254274 196608
rect 254394 196596 254400 196608
rect 254452 196596 254458 196648
rect 298465 196095 298523 196101
rect 298465 196061 298477 196095
rect 298511 196092 298523 196095
rect 298554 196092 298560 196104
rect 298511 196064 298560 196092
rect 298511 196061 298523 196064
rect 298465 196055 298523 196061
rect 298554 196052 298560 196064
rect 298612 196052 298618 196104
rect 327350 196052 327356 196104
rect 327408 196052 327414 196104
rect 273346 195984 273352 196036
rect 273404 196024 273410 196036
rect 273530 196024 273536 196036
rect 273404 195996 273536 196024
rect 273404 195984 273410 195996
rect 273530 195984 273536 195996
rect 273588 195984 273594 196036
rect 288710 196024 288716 196036
rect 288671 195996 288716 196024
rect 288710 195984 288716 195996
rect 288768 195984 288774 196036
rect 308030 196024 308036 196036
rect 307991 195996 308036 196024
rect 308030 195984 308036 195996
rect 308088 195984 308094 196036
rect 327368 195968 327396 196052
rect 434438 196024 434444 196036
rect 434399 195996 434444 196024
rect 434438 195984 434444 195996
rect 434496 195984 434502 196036
rect 299842 195916 299848 195968
rect 299900 195916 299906 195968
rect 305270 195956 305276 195968
rect 305231 195928 305276 195956
rect 305270 195916 305276 195928
rect 305328 195916 305334 195968
rect 325970 195916 325976 195968
rect 326028 195916 326034 195968
rect 327350 195916 327356 195968
rect 327408 195916 327414 195968
rect 299860 195832 299888 195916
rect 325988 195832 326016 195916
rect 435174 195848 435180 195900
rect 435232 195888 435238 195900
rect 435358 195888 435364 195900
rect 435232 195860 435364 195888
rect 435232 195848 435238 195860
rect 435358 195848 435364 195860
rect 435416 195848 435422 195900
rect 299842 195780 299848 195832
rect 299900 195780 299906 195832
rect 325970 195780 325976 195832
rect 326028 195780 326034 195832
rect 262582 193332 262588 193384
rect 262640 193332 262646 193384
rect 262600 193248 262628 193332
rect 345106 193264 345112 193316
rect 345164 193264 345170 193316
rect 229370 193196 229376 193248
rect 229428 193236 229434 193248
rect 229554 193236 229560 193248
rect 229428 193208 229560 193236
rect 229428 193196 229434 193208
rect 229554 193196 229560 193208
rect 229612 193196 229618 193248
rect 235074 193196 235080 193248
rect 235132 193196 235138 193248
rect 239122 193196 239128 193248
rect 239180 193196 239186 193248
rect 244090 193196 244096 193248
rect 244148 193236 244154 193248
rect 244274 193236 244280 193248
rect 244148 193208 244280 193236
rect 244148 193196 244154 193208
rect 244274 193196 244280 193208
rect 244332 193196 244338 193248
rect 262582 193196 262588 193248
rect 262640 193196 262646 193248
rect 287330 193196 287336 193248
rect 287388 193236 287394 193248
rect 287514 193236 287520 193248
rect 287388 193208 287520 193236
rect 287388 193196 287394 193208
rect 287514 193196 287520 193208
rect 287572 193196 287578 193248
rect 288713 193239 288771 193245
rect 288713 193205 288725 193239
rect 288759 193236 288771 193239
rect 288802 193236 288808 193248
rect 288759 193208 288808 193236
rect 288759 193205 288771 193208
rect 288713 193199 288771 193205
rect 288802 193196 288808 193208
rect 288860 193196 288866 193248
rect 298462 193236 298468 193248
rect 298423 193208 298468 193236
rect 298462 193196 298468 193208
rect 298520 193196 298526 193248
rect 308030 193236 308036 193248
rect 307991 193208 308036 193236
rect 308030 193196 308036 193208
rect 308088 193196 308094 193248
rect 324590 193196 324596 193248
rect 324648 193236 324654 193248
rect 324682 193236 324688 193248
rect 324648 193208 324688 193236
rect 324648 193196 324654 193208
rect 324682 193196 324688 193208
rect 324740 193196 324746 193248
rect 235092 193168 235120 193196
rect 235258 193168 235264 193180
rect 235092 193140 235264 193168
rect 235258 193128 235264 193140
rect 235316 193128 235322 193180
rect 239140 193168 239168 193196
rect 345124 193180 345152 193264
rect 362954 193196 362960 193248
rect 363012 193236 363018 193248
rect 363230 193236 363236 193248
rect 363012 193208 363236 193236
rect 363012 193196 363018 193208
rect 363230 193196 363236 193208
rect 363288 193196 363294 193248
rect 434438 193236 434444 193248
rect 434399 193208 434444 193236
rect 434438 193196 434444 193208
rect 434496 193196 434502 193248
rect 239214 193168 239220 193180
rect 239140 193140 239220 193168
rect 239214 193128 239220 193140
rect 239272 193128 239278 193180
rect 240413 193171 240471 193177
rect 240413 193137 240425 193171
rect 240459 193168 240471 193171
rect 240502 193168 240508 193180
rect 240459 193140 240508 193168
rect 240459 193137 240471 193140
rect 240413 193131 240471 193137
rect 240502 193128 240508 193140
rect 240560 193128 240566 193180
rect 345106 193128 345112 193180
rect 345164 193128 345170 193180
rect 345014 192760 345020 192772
rect 344975 192732 345020 192760
rect 345014 192720 345020 192732
rect 345072 192720 345078 192772
rect 234798 192284 234804 192296
rect 234759 192256 234804 192284
rect 234798 192244 234804 192256
rect 234856 192244 234862 192296
rect 251450 191836 251456 191888
rect 251508 191876 251514 191888
rect 251542 191876 251548 191888
rect 251508 191848 251548 191876
rect 251508 191836 251514 191848
rect 251542 191836 251548 191848
rect 251600 191836 251606 191888
rect 316221 191879 316279 191885
rect 316221 191845 316233 191879
rect 316267 191876 316279 191879
rect 316310 191876 316316 191888
rect 316267 191848 316316 191876
rect 316267 191845 316279 191848
rect 316221 191839 316279 191845
rect 316310 191836 316316 191848
rect 316368 191836 316374 191888
rect 255590 191808 255596 191820
rect 255551 191780 255596 191808
rect 255590 191768 255596 191780
rect 255648 191768 255654 191820
rect 262582 191808 262588 191820
rect 262543 191780 262588 191808
rect 262582 191768 262588 191780
rect 262640 191768 262646 191820
rect 345014 190612 345020 190664
rect 345072 190652 345078 190664
rect 345290 190652 345296 190664
rect 345072 190624 345296 190652
rect 345072 190612 345078 190624
rect 345290 190612 345296 190624
rect 345348 190612 345354 190664
rect 266998 190516 267004 190528
rect 266959 190488 267004 190516
rect 266998 190476 267004 190488
rect 267056 190476 267062 190528
rect 316218 190516 316224 190528
rect 316179 190488 316224 190516
rect 316218 190476 316224 190488
rect 316276 190476 316282 190528
rect 244274 189388 244280 189440
rect 244332 189428 244338 189440
rect 244458 189428 244464 189440
rect 244332 189400 244464 189428
rect 244332 189388 244338 189400
rect 244458 189388 244464 189400
rect 244516 189388 244522 189440
rect 261202 186396 261208 186448
rect 261260 186396 261266 186448
rect 276290 186436 276296 186448
rect 276124 186408 276296 186436
rect 233326 186328 233332 186380
rect 233384 186368 233390 186380
rect 233510 186368 233516 186380
rect 233384 186340 233516 186368
rect 233384 186328 233390 186340
rect 233510 186328 233516 186340
rect 233568 186328 233574 186380
rect 238754 186328 238760 186380
rect 238812 186368 238818 186380
rect 238938 186368 238944 186380
rect 238812 186340 238944 186368
rect 238812 186328 238818 186340
rect 238938 186328 238944 186340
rect 238996 186328 239002 186380
rect 261220 186312 261248 186396
rect 276124 186380 276152 186408
rect 276290 186396 276296 186408
rect 276348 186396 276354 186448
rect 276106 186328 276112 186380
rect 276164 186328 276170 186380
rect 288802 186368 288808 186380
rect 288763 186340 288808 186368
rect 288802 186328 288808 186340
rect 288860 186328 288866 186380
rect 327350 186328 327356 186380
rect 327408 186328 327414 186380
rect 346578 186328 346584 186380
rect 346636 186328 346642 186380
rect 444006 186328 444012 186380
rect 444064 186368 444070 186380
rect 444190 186368 444196 186380
rect 444064 186340 444196 186368
rect 444064 186328 444070 186340
rect 444190 186328 444196 186340
rect 444248 186328 444254 186380
rect 255590 186300 255596 186312
rect 255551 186272 255596 186300
rect 255590 186260 255596 186272
rect 255648 186260 255654 186312
rect 261202 186260 261208 186312
rect 261260 186260 261266 186312
rect 280430 186260 280436 186312
rect 280488 186300 280494 186312
rect 280614 186300 280620 186312
rect 280488 186272 280620 186300
rect 280488 186260 280494 186272
rect 280614 186260 280620 186272
rect 280672 186260 280678 186312
rect 327368 186232 327396 186328
rect 327442 186232 327448 186244
rect 327368 186204 327448 186232
rect 327442 186192 327448 186204
rect 327500 186192 327506 186244
rect 346596 186232 346624 186328
rect 346670 186232 346676 186244
rect 346596 186204 346676 186232
rect 346670 186192 346676 186204
rect 346728 186192 346734 186244
rect 310422 185580 310428 185632
rect 310480 185620 310486 185632
rect 310793 185623 310851 185629
rect 310793 185620 310805 185623
rect 310480 185592 310805 185620
rect 310480 185580 310486 185592
rect 310793 185589 310805 185592
rect 310839 185589 310851 185623
rect 310793 185583 310851 185589
rect 241882 183648 241888 183660
rect 241808 183620 241888 183648
rect 241808 183592 241836 183620
rect 241882 183608 241888 183620
rect 241940 183608 241946 183660
rect 434438 183648 434444 183660
rect 434272 183620 434444 183648
rect 434272 183592 434300 183620
rect 434438 183608 434444 183620
rect 434496 183608 434502 183660
rect 234982 183540 234988 183592
rect 235040 183580 235046 183592
rect 235258 183580 235264 183592
rect 235040 183552 235264 183580
rect 235040 183540 235046 183552
rect 235258 183540 235264 183552
rect 235316 183540 235322 183592
rect 239122 183540 239128 183592
rect 239180 183580 239186 183592
rect 239214 183580 239220 183592
rect 239180 183552 239220 183580
rect 239180 183540 239186 183552
rect 239214 183540 239220 183552
rect 239272 183540 239278 183592
rect 241790 183540 241796 183592
rect 241848 183540 241854 183592
rect 288802 183580 288808 183592
rect 288763 183552 288808 183580
rect 288802 183540 288808 183552
rect 288860 183540 288866 183592
rect 305178 183540 305184 183592
rect 305236 183580 305242 183592
rect 305454 183580 305460 183592
rect 305236 183552 305460 183580
rect 305236 183540 305242 183552
rect 305454 183540 305460 183552
rect 305512 183540 305518 183592
rect 308122 183540 308128 183592
rect 308180 183580 308186 183592
rect 308306 183580 308312 183592
rect 308180 183552 308312 183580
rect 308180 183540 308186 183552
rect 308306 183540 308312 183552
rect 308364 183540 308370 183592
rect 342346 183540 342352 183592
rect 342404 183580 342410 183592
rect 342530 183580 342536 183592
rect 342404 183552 342536 183580
rect 342404 183540 342410 183552
rect 342530 183540 342536 183552
rect 342588 183540 342594 183592
rect 347958 183540 347964 183592
rect 348016 183580 348022 183592
rect 348142 183580 348148 183592
rect 348016 183552 348148 183580
rect 348016 183540 348022 183552
rect 348142 183540 348148 183552
rect 348200 183540 348206 183592
rect 434254 183540 434260 183592
rect 434312 183540 434318 183592
rect 262582 183512 262588 183524
rect 262543 183484 262588 183512
rect 262582 183472 262588 183484
rect 262640 183472 262646 183524
rect 343818 183472 343824 183524
rect 343876 183512 343882 183524
rect 343910 183512 343916 183524
rect 343876 183484 343916 183512
rect 343876 183472 343882 183484
rect 343910 183472 343916 183484
rect 343968 183472 343974 183524
rect 316218 182180 316224 182232
rect 316276 182220 316282 182232
rect 316310 182220 316316 182232
rect 316276 182192 316316 182220
rect 316276 182180 316282 182192
rect 316310 182180 316316 182192
rect 316368 182180 316374 182232
rect 239122 182152 239128 182164
rect 239083 182124 239128 182152
rect 239122 182112 239128 182124
rect 239180 182112 239186 182164
rect 255593 182155 255651 182161
rect 255593 182121 255605 182155
rect 255639 182152 255651 182155
rect 255682 182152 255688 182164
rect 255639 182124 255688 182152
rect 255639 182121 255651 182124
rect 255593 182115 255651 182121
rect 255682 182112 255688 182124
rect 255740 182112 255746 182164
rect 324498 182112 324504 182164
rect 324556 182152 324562 182164
rect 324682 182152 324688 182164
rect 324556 182124 324688 182152
rect 324556 182112 324562 182124
rect 324682 182112 324688 182124
rect 324740 182112 324746 182164
rect 343910 182112 343916 182164
rect 343968 182152 343974 182164
rect 344094 182152 344100 182164
rect 343968 182124 344100 182152
rect 343968 182112 343974 182124
rect 344094 182112 344100 182124
rect 344152 182112 344158 182164
rect 309042 181024 309048 181076
rect 309100 181064 309106 181076
rect 312078 181064 312084 181076
rect 309100 181036 312084 181064
rect 309100 181024 309106 181036
rect 312078 181024 312084 181036
rect 312136 181024 312142 181076
rect 398466 180956 398472 181008
rect 398524 180996 398530 181008
rect 399018 180996 399024 181008
rect 398524 180968 399024 180996
rect 398524 180956 398530 180968
rect 399018 180956 399024 180968
rect 399076 180956 399082 181008
rect 417878 180956 417884 181008
rect 417936 180996 417942 181008
rect 418338 180996 418344 181008
rect 417936 180968 418344 180996
rect 417936 180956 417942 180968
rect 418338 180956 418344 180968
rect 418396 180956 418402 181008
rect 338022 180888 338028 180940
rect 338080 180888 338086 180940
rect 454402 180888 454408 180940
rect 454460 180928 454466 180940
rect 458358 180928 458364 180940
rect 454460 180900 458364 180928
rect 454460 180888 454466 180900
rect 458358 180888 458364 180900
rect 458416 180888 458422 180940
rect 270494 180820 270500 180872
rect 270552 180860 270558 180872
rect 275370 180860 275376 180872
rect 270552 180832 275376 180860
rect 270552 180820 270558 180832
rect 275370 180820 275376 180832
rect 275428 180820 275434 180872
rect 338040 180804 338068 180888
rect 313642 180752 313648 180804
rect 313700 180792 313706 180804
rect 313734 180792 313740 180804
rect 313700 180764 313740 180792
rect 313700 180752 313706 180764
rect 313734 180752 313740 180764
rect 313792 180752 313798 180804
rect 327353 180795 327411 180801
rect 327353 180761 327365 180795
rect 327399 180792 327411 180795
rect 327442 180792 327448 180804
rect 327399 180764 327448 180792
rect 327399 180761 327411 180764
rect 327353 180755 327411 180761
rect 327442 180752 327448 180764
rect 327500 180752 327506 180804
rect 338022 180752 338028 180804
rect 338080 180752 338086 180804
rect 2774 179800 2780 179852
rect 2832 179840 2838 179852
rect 5074 179840 5080 179852
rect 2832 179812 5080 179840
rect 2832 179800 2838 179812
rect 5074 179800 5080 179812
rect 5132 179800 5138 179852
rect 234982 179324 234988 179376
rect 235040 179364 235046 179376
rect 235166 179364 235172 179376
rect 235040 179336 235172 179364
rect 235040 179324 235046 179336
rect 235166 179324 235172 179336
rect 235224 179324 235230 179376
rect 310790 179364 310796 179376
rect 310751 179336 310796 179364
rect 310790 179324 310796 179336
rect 310848 179324 310854 179376
rect 241790 178820 241796 178832
rect 241751 178792 241796 178820
rect 241790 178780 241796 178792
rect 241848 178780 241854 178832
rect 248782 176780 248788 176792
rect 248708 176752 248788 176780
rect 248708 176656 248736 176752
rect 248782 176740 248788 176752
rect 248840 176740 248846 176792
rect 288802 176740 288808 176792
rect 288860 176740 288866 176792
rect 287238 176672 287244 176724
rect 287296 176712 287302 176724
rect 287296 176684 287376 176712
rect 287296 176672 287302 176684
rect 287348 176656 287376 176684
rect 288820 176656 288848 176740
rect 238754 176604 238760 176656
rect 238812 176644 238818 176656
rect 238938 176644 238944 176656
rect 238812 176616 238944 176644
rect 238812 176604 238818 176616
rect 238938 176604 238944 176616
rect 238996 176604 239002 176656
rect 248690 176604 248696 176656
rect 248748 176604 248754 176656
rect 276106 176604 276112 176656
rect 276164 176604 276170 176656
rect 287330 176604 287336 176656
rect 287388 176604 287394 176656
rect 288802 176604 288808 176656
rect 288860 176604 288866 176656
rect 276124 176576 276152 176604
rect 276290 176576 276296 176588
rect 276124 176548 276296 176576
rect 276290 176536 276296 176548
rect 276348 176536 276354 176588
rect 267090 173992 267096 174004
rect 267016 173964 267096 173992
rect 267016 173936 267044 173964
rect 267090 173952 267096 173964
rect 267148 173952 267154 174004
rect 299842 173992 299848 174004
rect 299768 173964 299848 173992
rect 299768 173936 299796 173964
rect 299842 173952 299848 173964
rect 299900 173952 299906 174004
rect 229370 173884 229376 173936
rect 229428 173924 229434 173936
rect 229554 173924 229560 173936
rect 229428 173896 229560 173924
rect 229428 173884 229434 173896
rect 229554 173884 229560 173896
rect 229612 173884 229618 173936
rect 234798 173884 234804 173936
rect 234856 173924 234862 173936
rect 234890 173924 234896 173936
rect 234856 173896 234896 173924
rect 234856 173884 234862 173896
rect 234890 173884 234896 173896
rect 234948 173884 234954 173936
rect 240410 173884 240416 173936
rect 240468 173924 240474 173936
rect 240502 173924 240508 173936
rect 240468 173896 240508 173924
rect 240468 173884 240474 173896
rect 240502 173884 240508 173896
rect 240560 173884 240566 173936
rect 241790 173924 241796 173936
rect 241751 173896 241796 173924
rect 241790 173884 241796 173896
rect 241848 173884 241854 173936
rect 244274 173884 244280 173936
rect 244332 173924 244338 173936
rect 244458 173924 244464 173936
rect 244332 173896 244464 173924
rect 244332 173884 244338 173896
rect 244458 173884 244464 173896
rect 244516 173884 244522 173936
rect 261202 173884 261208 173936
rect 261260 173924 261266 173936
rect 261294 173924 261300 173936
rect 261260 173896 261300 173924
rect 261260 173884 261266 173896
rect 261294 173884 261300 173896
rect 261352 173884 261358 173936
rect 262674 173884 262680 173936
rect 262732 173884 262738 173936
rect 266998 173884 267004 173936
rect 267056 173884 267062 173936
rect 291378 173884 291384 173936
rect 291436 173924 291442 173936
rect 291470 173924 291476 173936
rect 291436 173896 291476 173924
rect 291436 173884 291442 173896
rect 291470 173884 291476 173896
rect 291528 173884 291534 173936
rect 299750 173884 299756 173936
rect 299808 173884 299814 173936
rect 305362 173884 305368 173936
rect 305420 173924 305426 173936
rect 305454 173924 305460 173936
rect 305420 173896 305460 173924
rect 305420 173884 305426 173896
rect 305454 173884 305460 173896
rect 305512 173884 305518 173936
rect 308030 173884 308036 173936
rect 308088 173924 308094 173936
rect 308214 173924 308220 173936
rect 308088 173896 308220 173924
rect 308088 173884 308094 173896
rect 308214 173884 308220 173896
rect 308272 173884 308278 173936
rect 362954 173884 362960 173936
rect 363012 173924 363018 173936
rect 363230 173924 363236 173936
rect 363012 173896 363236 173924
rect 363012 173884 363018 173896
rect 363230 173884 363236 173896
rect 363288 173884 363294 173936
rect 443914 173884 443920 173936
rect 443972 173924 443978 173936
rect 444098 173924 444104 173936
rect 443972 173896 444104 173924
rect 443972 173884 443978 173896
rect 444098 173884 444104 173896
rect 444156 173884 444162 173936
rect 239122 173856 239128 173868
rect 239083 173828 239128 173856
rect 239122 173816 239128 173828
rect 239180 173816 239186 173868
rect 262692 173788 262720 173884
rect 262766 173788 262772 173800
rect 262692 173760 262772 173788
rect 262766 173748 262772 173760
rect 262824 173748 262830 173800
rect 255590 172564 255596 172576
rect 255551 172536 255596 172564
rect 255590 172524 255596 172536
rect 255648 172524 255654 172576
rect 251358 172456 251364 172508
rect 251416 172496 251422 172508
rect 251450 172496 251456 172508
rect 251416 172468 251456 172496
rect 251416 172456 251422 172468
rect 251450 172456 251456 172468
rect 251508 172456 251514 172508
rect 299750 172456 299756 172508
rect 299808 172496 299814 172508
rect 300026 172496 300032 172508
rect 299808 172468 300032 172496
rect 299808 172456 299814 172468
rect 300026 172456 300032 172468
rect 300084 172456 300090 172508
rect 327350 171136 327356 171148
rect 327311 171108 327356 171136
rect 327350 171096 327356 171108
rect 327408 171096 327414 171148
rect 251358 171068 251364 171080
rect 251319 171040 251364 171068
rect 251358 171028 251364 171040
rect 251416 171028 251422 171080
rect 313550 171068 313556 171080
rect 313511 171040 313556 171068
rect 313550 171028 313556 171040
rect 313608 171028 313614 171080
rect 345014 171028 345020 171080
rect 345072 171068 345078 171080
rect 345198 171068 345204 171080
rect 345072 171040 345204 171068
rect 345072 171028 345078 171040
rect 345198 171028 345204 171040
rect 345256 171028 345262 171080
rect 310793 169779 310851 169785
rect 310793 169745 310805 169779
rect 310839 169776 310851 169779
rect 310882 169776 310888 169788
rect 310839 169748 310888 169776
rect 310839 169745 310851 169748
rect 310793 169739 310851 169745
rect 310882 169736 310888 169748
rect 310940 169736 310946 169788
rect 239122 169056 239128 169108
rect 239180 169096 239186 169108
rect 239306 169096 239312 169108
rect 239180 169068 239312 169096
rect 239180 169056 239186 169068
rect 239306 169056 239312 169068
rect 239364 169056 239370 169108
rect 233326 167016 233332 167068
rect 233384 167056 233390 167068
rect 233510 167056 233516 167068
rect 233384 167028 233516 167056
rect 233384 167016 233390 167028
rect 233510 167016 233516 167028
rect 233568 167016 233574 167068
rect 238754 167016 238760 167068
rect 238812 167056 238818 167068
rect 238938 167056 238944 167068
rect 238812 167028 238944 167056
rect 238812 167016 238818 167028
rect 238938 167016 238944 167028
rect 238996 167016 239002 167068
rect 346486 167016 346492 167068
rect 346544 167056 346550 167068
rect 346670 167056 346676 167068
rect 346544 167028 346676 167056
rect 346544 167016 346550 167028
rect 346670 167016 346676 167028
rect 346728 167016 346734 167068
rect 435174 167016 435180 167068
rect 435232 167056 435238 167068
rect 435358 167056 435364 167068
rect 435232 167028 435364 167056
rect 435232 167016 435238 167028
rect 435358 167016 435364 167028
rect 435416 167016 435422 167068
rect 2774 165452 2780 165504
rect 2832 165492 2838 165504
rect 4982 165492 4988 165504
rect 2832 165464 4988 165492
rect 2832 165452 2838 165464
rect 4982 165452 4988 165464
rect 5040 165452 5046 165504
rect 435174 165044 435180 165096
rect 435232 165084 435238 165096
rect 435542 165084 435548 165096
rect 435232 165056 435548 165084
rect 435232 165044 435238 165056
rect 435542 165044 435548 165056
rect 435600 165044 435606 165096
rect 255590 164228 255596 164280
rect 255648 164228 255654 164280
rect 262674 164228 262680 164280
rect 262732 164268 262738 164280
rect 262766 164268 262772 164280
rect 262732 164240 262772 164268
rect 262732 164228 262738 164240
rect 262766 164228 262772 164240
rect 262824 164228 262830 164280
rect 254210 164160 254216 164212
rect 254268 164200 254274 164212
rect 254394 164200 254400 164212
rect 254268 164172 254400 164200
rect 254268 164160 254274 164172
rect 254394 164160 254400 164172
rect 254452 164160 254458 164212
rect 255608 164132 255636 164228
rect 287330 164200 287336 164212
rect 287291 164172 287336 164200
rect 287330 164160 287336 164172
rect 287388 164160 287394 164212
rect 324593 164203 324651 164209
rect 324593 164169 324605 164203
rect 324639 164200 324651 164203
rect 324682 164200 324688 164212
rect 324639 164172 324688 164200
rect 324639 164169 324651 164172
rect 324593 164163 324651 164169
rect 324682 164160 324688 164172
rect 324740 164160 324746 164212
rect 362954 164160 362960 164212
rect 363012 164200 363018 164212
rect 363138 164200 363144 164212
rect 363012 164172 363144 164200
rect 363012 164160 363018 164172
rect 363138 164160 363144 164172
rect 363196 164160 363202 164212
rect 444098 164200 444104 164212
rect 444059 164172 444104 164200
rect 444098 164160 444104 164172
rect 444156 164160 444162 164212
rect 255682 164132 255688 164144
rect 255608 164104 255688 164132
rect 255682 164092 255688 164104
rect 255740 164092 255746 164144
rect 234982 162936 234988 162988
rect 235040 162976 235046 162988
rect 235166 162976 235172 162988
rect 235040 162948 235172 162976
rect 235040 162936 235046 162948
rect 235166 162936 235172 162948
rect 235224 162936 235230 162988
rect 241882 162840 241888 162852
rect 241843 162812 241888 162840
rect 241882 162800 241888 162812
rect 241940 162800 241946 162852
rect 261297 162843 261355 162849
rect 261297 162809 261309 162843
rect 261343 162840 261355 162843
rect 261386 162840 261392 162852
rect 261343 162812 261392 162840
rect 261343 162809 261355 162812
rect 261297 162803 261355 162809
rect 261386 162800 261392 162812
rect 261444 162800 261450 162852
rect 262493 162843 262551 162849
rect 262493 162809 262505 162843
rect 262539 162840 262551 162843
rect 262674 162840 262680 162852
rect 262539 162812 262680 162840
rect 262539 162809 262551 162812
rect 262493 162803 262551 162809
rect 262674 162800 262680 162812
rect 262732 162800 262738 162852
rect 288710 162800 288716 162852
rect 288768 162840 288774 162852
rect 288802 162840 288808 162852
rect 288768 162812 288808 162840
rect 288768 162800 288774 162812
rect 288802 162800 288808 162812
rect 288860 162800 288866 162852
rect 305273 162843 305331 162849
rect 305273 162809 305285 162843
rect 305319 162840 305331 162843
rect 305362 162840 305368 162852
rect 305319 162812 305368 162840
rect 305319 162809 305331 162812
rect 305273 162803 305331 162809
rect 305362 162800 305368 162812
rect 305420 162800 305426 162852
rect 342530 162800 342536 162852
rect 342588 162840 342594 162852
rect 342622 162840 342628 162852
rect 342588 162812 342628 162840
rect 342588 162800 342594 162812
rect 342622 162800 342628 162812
rect 342680 162800 342686 162852
rect 343910 162840 343916 162852
rect 343871 162812 343916 162840
rect 343910 162800 343916 162812
rect 343968 162800 343974 162852
rect 345198 162840 345204 162852
rect 345159 162812 345204 162840
rect 345198 162800 345204 162812
rect 345256 162800 345262 162852
rect 251361 161483 251419 161489
rect 251361 161449 251373 161483
rect 251407 161480 251419 161483
rect 251450 161480 251456 161492
rect 251407 161452 251456 161480
rect 251407 161449 251419 161452
rect 251361 161443 251419 161449
rect 251450 161440 251456 161452
rect 251508 161440 251514 161492
rect 313553 161483 313611 161489
rect 313553 161449 313565 161483
rect 313599 161480 313611 161483
rect 313826 161480 313832 161492
rect 313599 161452 313832 161480
rect 313599 161449 313611 161452
rect 313553 161443 313611 161449
rect 313826 161440 313832 161452
rect 313884 161440 313890 161492
rect 234982 161412 234988 161424
rect 234943 161384 234988 161412
rect 234982 161372 234988 161384
rect 235040 161372 235046 161424
rect 288710 161412 288716 161424
rect 288671 161384 288716 161412
rect 288710 161372 288716 161384
rect 288768 161372 288774 161424
rect 308033 161415 308091 161421
rect 308033 161381 308045 161415
rect 308079 161412 308091 161415
rect 308122 161412 308128 161424
rect 308079 161384 308128 161412
rect 308079 161381 308091 161384
rect 308033 161375 308091 161381
rect 308122 161372 308128 161384
rect 308180 161372 308186 161424
rect 310882 161372 310888 161424
rect 310940 161412 310946 161424
rect 310974 161412 310980 161424
rect 310940 161384 310980 161412
rect 310940 161372 310946 161384
rect 310974 161372 310980 161384
rect 311032 161372 311038 161424
rect 234890 161344 234896 161356
rect 234851 161316 234896 161344
rect 234890 161304 234896 161316
rect 234948 161304 234954 161356
rect 238846 159712 238852 159724
rect 238807 159684 238852 159712
rect 238846 159672 238852 159684
rect 238904 159672 238910 159724
rect 238846 159372 238852 159384
rect 238807 159344 238852 159372
rect 238846 159332 238852 159344
rect 238904 159332 238910 159384
rect 434438 159168 434444 159180
rect 434399 159140 434444 159168
rect 434438 159128 434444 159140
rect 434496 159128 434502 159180
rect 229278 157360 229284 157412
rect 229336 157360 229342 157412
rect 280522 157360 280528 157412
rect 280580 157360 280586 157412
rect 229296 157332 229324 157360
rect 229370 157332 229376 157344
rect 229296 157304 229376 157332
rect 229370 157292 229376 157304
rect 229428 157292 229434 157344
rect 280540 157264 280568 157360
rect 325970 157292 325976 157344
rect 326028 157292 326034 157344
rect 444098 157332 444104 157344
rect 444059 157304 444104 157332
rect 444098 157292 444104 157304
rect 444156 157292 444162 157344
rect 280614 157264 280620 157276
rect 280540 157236 280620 157264
rect 280614 157224 280620 157236
rect 280672 157224 280678 157276
rect 325988 157208 326016 157292
rect 325970 157156 325976 157208
rect 326028 157156 326034 157208
rect 239033 154683 239091 154689
rect 239033 154649 239045 154683
rect 239079 154680 239091 154683
rect 239122 154680 239128 154692
rect 239079 154652 239128 154680
rect 239079 154649 239091 154652
rect 239033 154643 239091 154649
rect 239122 154640 239128 154652
rect 239180 154640 239186 154692
rect 255590 154640 255596 154692
rect 255648 154680 255654 154692
rect 255682 154680 255688 154692
rect 255648 154652 255688 154680
rect 255648 154640 255654 154652
rect 255682 154640 255688 154652
rect 255740 154640 255746 154692
rect 240413 154615 240471 154621
rect 240413 154581 240425 154615
rect 240459 154612 240471 154615
rect 240502 154612 240508 154624
rect 240459 154584 240508 154612
rect 240459 154581 240471 154584
rect 240413 154575 240471 154581
rect 240502 154572 240508 154584
rect 240560 154572 240566 154624
rect 287330 154612 287336 154624
rect 287291 154584 287336 154612
rect 287330 154572 287336 154584
rect 287388 154572 287394 154624
rect 324590 154612 324596 154624
rect 324551 154584 324596 154612
rect 324590 154572 324596 154584
rect 324648 154572 324654 154624
rect 434438 154612 434444 154624
rect 434399 154584 434444 154612
rect 434438 154572 434444 154584
rect 434496 154572 434502 154624
rect 229370 154504 229376 154556
rect 229428 154544 229434 154556
rect 229554 154544 229560 154556
rect 229428 154516 229560 154544
rect 229428 154504 229434 154516
rect 229554 154504 229560 154516
rect 229612 154504 229618 154556
rect 245746 154504 245752 154556
rect 245804 154544 245810 154556
rect 245930 154544 245936 154556
rect 245804 154516 245936 154544
rect 245804 154504 245810 154516
rect 245930 154504 245936 154516
rect 245988 154504 245994 154556
rect 290090 154504 290096 154556
rect 290148 154544 290154 154556
rect 290182 154544 290188 154556
rect 290148 154516 290188 154544
rect 290148 154504 290154 154516
rect 290182 154504 290188 154516
rect 290240 154504 290246 154556
rect 316310 154504 316316 154556
rect 316368 154544 316374 154556
rect 316402 154544 316408 154556
rect 316368 154516 316408 154544
rect 316368 154504 316374 154516
rect 316402 154504 316408 154516
rect 316460 154504 316466 154556
rect 347958 154504 347964 154556
rect 348016 154544 348022 154556
rect 348142 154544 348148 154556
rect 348016 154516 348148 154544
rect 348016 154504 348022 154516
rect 348142 154504 348148 154516
rect 348200 154504 348206 154556
rect 444101 154547 444159 154553
rect 444101 154513 444113 154547
rect 444147 154544 444159 154547
rect 444190 154544 444196 154556
rect 444147 154516 444196 154544
rect 444147 154513 444159 154516
rect 444101 154507 444159 154513
rect 444190 154504 444196 154516
rect 444248 154504 444254 154556
rect 288713 153867 288771 153873
rect 288713 153833 288725 153867
rect 288759 153864 288771 153867
rect 288802 153864 288808 153876
rect 288759 153836 288808 153864
rect 288759 153833 288771 153836
rect 288713 153827 288771 153833
rect 288802 153824 288808 153836
rect 288860 153824 288866 153876
rect 327350 153524 327356 153536
rect 327311 153496 327356 153524
rect 327350 153484 327356 153496
rect 327408 153484 327414 153536
rect 240410 153320 240416 153332
rect 240371 153292 240416 153320
rect 240410 153280 240416 153292
rect 240468 153280 240474 153332
rect 241882 153252 241888 153264
rect 241843 153224 241888 153252
rect 241882 153212 241888 153224
rect 241940 153212 241946 153264
rect 261294 153252 261300 153264
rect 261255 153224 261300 153252
rect 261294 153212 261300 153224
rect 261352 153212 261358 153264
rect 262490 153252 262496 153264
rect 262451 153224 262496 153252
rect 262490 153212 262496 153224
rect 262548 153212 262554 153264
rect 305270 153252 305276 153264
rect 305231 153224 305276 153252
rect 305270 153212 305276 153224
rect 305328 153212 305334 153264
rect 343910 153252 343916 153264
rect 343871 153224 343916 153252
rect 343910 153212 343916 153224
rect 343968 153212 343974 153264
rect 240321 153187 240379 153193
rect 240321 153153 240333 153187
rect 240367 153184 240379 153187
rect 240410 153184 240416 153196
rect 240367 153156 240416 153184
rect 240367 153153 240379 153156
rect 240321 153147 240379 153153
rect 240410 153144 240416 153156
rect 240468 153144 240474 153196
rect 255314 153144 255320 153196
rect 255372 153184 255378 153196
rect 255590 153184 255596 153196
rect 255372 153156 255596 153184
rect 255372 153144 255378 153156
rect 255590 153144 255596 153156
rect 255648 153144 255654 153196
rect 305270 153116 305276 153128
rect 305231 153088 305276 153116
rect 305270 153076 305276 153088
rect 305328 153076 305334 153128
rect 234985 151827 235043 151833
rect 234985 151793 234997 151827
rect 235031 151824 235043 151827
rect 235074 151824 235080 151836
rect 235031 151796 235080 151824
rect 235031 151793 235043 151796
rect 234985 151787 235043 151793
rect 235074 151784 235080 151796
rect 235132 151784 235138 151836
rect 239030 151824 239036 151836
rect 238991 151796 239036 151824
rect 239030 151784 239036 151796
rect 239088 151784 239094 151836
rect 251174 151784 251180 151836
rect 251232 151824 251238 151836
rect 251358 151824 251364 151836
rect 251232 151796 251364 151824
rect 251232 151784 251238 151796
rect 251358 151784 251364 151796
rect 251416 151784 251422 151836
rect 308030 151824 308036 151836
rect 307991 151796 308036 151824
rect 308030 151784 308036 151796
rect 308088 151784 308094 151836
rect 313645 150603 313703 150609
rect 313645 150569 313657 150603
rect 313691 150600 313703 150603
rect 313826 150600 313832 150612
rect 313691 150572 313832 150600
rect 313691 150569 313703 150572
rect 313645 150563 313703 150569
rect 313826 150560 313832 150572
rect 313884 150560 313890 150612
rect 313642 150464 313648 150476
rect 313603 150436 313648 150464
rect 313642 150424 313648 150436
rect 313700 150424 313706 150476
rect 288802 149036 288808 149048
rect 288763 149008 288808 149036
rect 288802 148996 288808 149008
rect 288860 148996 288866 149048
rect 309502 149036 309508 149048
rect 309463 149008 309508 149036
rect 309502 148996 309508 149008
rect 309560 148996 309566 149048
rect 343821 148359 343879 148365
rect 343821 148325 343833 148359
rect 343867 148356 343879 148359
rect 343910 148356 343916 148368
rect 343867 148328 343916 148356
rect 343867 148325 343879 148328
rect 343821 148319 343879 148325
rect 343910 148316 343916 148328
rect 343968 148316 343974 148368
rect 238938 147772 238944 147824
rect 238996 147772 239002 147824
rect 435542 147772 435548 147824
rect 435600 147772 435606 147824
rect 238846 147704 238852 147756
rect 238904 147704 238910 147756
rect 233326 147636 233332 147688
rect 233384 147676 233390 147688
rect 233510 147676 233516 147688
rect 233384 147648 233516 147676
rect 233384 147636 233390 147648
rect 233510 147636 233516 147648
rect 233568 147636 233574 147688
rect 238864 147620 238892 147704
rect 238956 147620 238984 147772
rect 324590 147704 324596 147756
rect 324648 147704 324654 147756
rect 435450 147704 435456 147756
rect 435508 147704 435514 147756
rect 280430 147636 280436 147688
rect 280488 147676 280494 147688
rect 280614 147676 280620 147688
rect 280488 147648 280620 147676
rect 280488 147636 280494 147648
rect 280614 147636 280620 147648
rect 280672 147636 280678 147688
rect 324608 147620 324636 147704
rect 435468 147620 435496 147704
rect 435560 147620 435588 147772
rect 238846 147568 238852 147620
rect 238904 147568 238910 147620
rect 238938 147568 238944 147620
rect 238996 147568 239002 147620
rect 324590 147568 324596 147620
rect 324648 147568 324654 147620
rect 327350 147608 327356 147620
rect 327311 147580 327356 147608
rect 327350 147568 327356 147580
rect 327408 147568 327414 147620
rect 434438 147568 434444 147620
rect 434496 147608 434502 147620
rect 434714 147608 434720 147620
rect 434496 147580 434720 147608
rect 434496 147568 434502 147580
rect 434714 147568 434720 147580
rect 434772 147568 434778 147620
rect 435450 147568 435456 147620
rect 435508 147568 435514 147620
rect 435542 147568 435548 147620
rect 435600 147568 435606 147620
rect 287238 144984 287244 145036
rect 287296 145024 287302 145036
rect 287330 145024 287336 145036
rect 287296 144996 287336 145024
rect 287296 144984 287302 144996
rect 287330 144984 287336 144996
rect 287388 144984 287394 145036
rect 444098 145024 444104 145036
rect 444059 144996 444104 145024
rect 444098 144984 444104 144996
rect 444156 144984 444162 145036
rect 345201 144959 345259 144965
rect 345201 144925 345213 144959
rect 345247 144956 345259 144959
rect 345290 144956 345296 144968
rect 345247 144928 345296 144956
rect 345247 144925 345259 144928
rect 345201 144919 345259 144925
rect 345290 144916 345296 144928
rect 345348 144916 345354 144968
rect 241790 144848 241796 144900
rect 241848 144888 241854 144900
rect 241974 144888 241980 144900
rect 241848 144860 241980 144888
rect 241848 144848 241854 144860
rect 241974 144848 241980 144860
rect 242032 144848 242038 144900
rect 244090 144848 244096 144900
rect 244148 144888 244154 144900
rect 244274 144888 244280 144900
rect 244148 144860 244280 144888
rect 244148 144848 244154 144860
rect 244274 144848 244280 144860
rect 244332 144848 244338 144900
rect 254210 144848 254216 144900
rect 254268 144888 254274 144900
rect 254394 144888 254400 144900
rect 254268 144860 254400 144888
rect 254268 144848 254274 144860
rect 254394 144848 254400 144860
rect 254452 144848 254458 144900
rect 240318 143596 240324 143608
rect 240279 143568 240324 143596
rect 240318 143556 240324 143568
rect 240376 143556 240382 143608
rect 238754 143488 238760 143540
rect 238812 143528 238818 143540
rect 238938 143528 238944 143540
rect 238812 143500 238944 143528
rect 238812 143488 238818 143500
rect 238938 143488 238944 143500
rect 238996 143488 239002 143540
rect 239030 143488 239036 143540
rect 239088 143528 239094 143540
rect 239122 143528 239128 143540
rect 239088 143500 239128 143528
rect 239088 143488 239094 143500
rect 239122 143488 239128 143500
rect 239180 143488 239186 143540
rect 251358 143488 251364 143540
rect 251416 143528 251422 143540
rect 251545 143531 251603 143537
rect 251545 143528 251557 143531
rect 251416 143500 251557 143528
rect 251416 143488 251422 143500
rect 251545 143497 251557 143500
rect 251591 143497 251603 143531
rect 287238 143528 287244 143540
rect 287199 143500 287244 143528
rect 251545 143491 251603 143497
rect 287238 143488 287244 143500
rect 287296 143488 287302 143540
rect 345198 143488 345204 143540
rect 345256 143528 345262 143540
rect 345382 143528 345388 143540
rect 345256 143500 345388 143528
rect 345256 143488 345262 143500
rect 345382 143488 345388 143500
rect 345440 143488 345446 143540
rect 434438 143528 434444 143540
rect 434399 143500 434444 143528
rect 434438 143488 434444 143500
rect 434496 143488 434502 143540
rect 444098 143528 444104 143540
rect 444059 143500 444104 143528
rect 444098 143488 444104 143500
rect 444156 143488 444162 143540
rect 305273 142171 305331 142177
rect 305273 142137 305285 142171
rect 305319 142168 305331 142171
rect 305362 142168 305368 142180
rect 305319 142140 305368 142168
rect 305319 142137 305331 142140
rect 305273 142131 305331 142137
rect 305362 142128 305368 142140
rect 305420 142128 305426 142180
rect 239122 142100 239128 142112
rect 239083 142072 239128 142100
rect 239122 142060 239128 142072
rect 239180 142060 239186 142112
rect 240318 142100 240324 142112
rect 240279 142072 240324 142100
rect 240318 142060 240324 142072
rect 240376 142060 240382 142112
rect 316310 142100 316316 142112
rect 316271 142072 316316 142100
rect 316310 142060 316316 142072
rect 316368 142060 316374 142112
rect 234798 140836 234804 140888
rect 234856 140876 234862 140888
rect 234893 140879 234951 140885
rect 234893 140876 234905 140879
rect 234856 140848 234905 140876
rect 234856 140836 234862 140848
rect 234893 140845 234905 140848
rect 234939 140845 234951 140879
rect 234893 140839 234951 140845
rect 234798 140740 234804 140752
rect 234759 140712 234804 140740
rect 234798 140700 234804 140712
rect 234856 140700 234862 140752
rect 288802 139516 288808 139528
rect 288763 139488 288808 139516
rect 288802 139476 288808 139488
rect 288860 139476 288866 139528
rect 309502 139448 309508 139460
rect 309463 139420 309508 139448
rect 309502 139408 309508 139420
rect 309560 139408 309566 139460
rect 262674 139380 262680 139392
rect 262635 139352 262680 139380
rect 262674 139340 262680 139352
rect 262732 139340 262738 139392
rect 288802 139340 288808 139392
rect 288860 139380 288866 139392
rect 288894 139380 288900 139392
rect 288860 139352 288900 139380
rect 288860 139340 288866 139352
rect 288894 139340 288900 139352
rect 288952 139340 288958 139392
rect 267182 138088 267188 138100
rect 267108 138060 267188 138088
rect 229278 137980 229284 138032
rect 229336 137980 229342 138032
rect 229296 137952 229324 137980
rect 267108 137964 267136 138060
rect 267182 138048 267188 138060
rect 267240 138048 267246 138100
rect 435358 137980 435364 138032
rect 435416 138020 435422 138032
rect 435542 138020 435548 138032
rect 435416 137992 435548 138020
rect 435416 137980 435422 137992
rect 435542 137980 435548 137992
rect 435600 137980 435606 138032
rect 229370 137952 229376 137964
rect 229296 137924 229376 137952
rect 229370 137912 229376 137924
rect 229428 137912 229434 137964
rect 267090 137912 267096 137964
rect 267148 137912 267154 137964
rect 434441 137955 434499 137961
rect 434441 137921 434453 137955
rect 434487 137952 434499 137955
rect 434530 137952 434536 137964
rect 434487 137924 434536 137952
rect 434487 137921 434499 137924
rect 434441 137915 434499 137921
rect 434530 137912 434536 137924
rect 434588 137912 434594 137964
rect 287241 137819 287299 137825
rect 287241 137785 287253 137819
rect 287287 137816 287299 137819
rect 287422 137816 287428 137828
rect 287287 137788 287428 137816
rect 287287 137785 287299 137788
rect 287241 137779 287299 137785
rect 287422 137776 287428 137788
rect 287480 137776 287486 137828
rect 2774 136348 2780 136400
rect 2832 136388 2838 136400
rect 4890 136388 4896 136400
rect 2832 136360 4896 136388
rect 2832 136348 2838 136360
rect 4890 136348 4896 136360
rect 4948 136348 4954 136400
rect 343818 135300 343824 135312
rect 343779 135272 343824 135300
rect 343818 135260 343824 135272
rect 343876 135260 343882 135312
rect 346578 135260 346584 135312
rect 346636 135300 346642 135312
rect 346670 135300 346676 135312
rect 346636 135272 346676 135300
rect 346636 135260 346642 135272
rect 346670 135260 346676 135272
rect 346728 135260 346734 135312
rect 229370 135192 229376 135244
rect 229428 135232 229434 135244
rect 229554 135232 229560 135244
rect 229428 135204 229560 135232
rect 229428 135192 229434 135204
rect 229554 135192 229560 135204
rect 229612 135192 229618 135244
rect 241882 135232 241888 135244
rect 241843 135204 241888 135232
rect 241882 135192 241888 135204
rect 241940 135192 241946 135244
rect 245746 135192 245752 135244
rect 245804 135232 245810 135244
rect 245930 135232 245936 135244
rect 245804 135204 245936 135232
rect 245804 135192 245810 135204
rect 245930 135192 245936 135204
rect 245988 135192 245994 135244
rect 251542 135232 251548 135244
rect 251503 135204 251548 135232
rect 251542 135192 251548 135204
rect 251600 135192 251606 135244
rect 267090 135232 267096 135244
rect 267051 135204 267096 135232
rect 267090 135192 267096 135204
rect 267148 135192 267154 135244
rect 327350 135232 327356 135244
rect 327311 135204 327356 135232
rect 327350 135192 327356 135204
rect 327408 135192 327414 135244
rect 328546 135192 328552 135244
rect 328604 135232 328610 135244
rect 328730 135232 328736 135244
rect 328604 135204 328736 135232
rect 328604 135192 328610 135204
rect 328730 135192 328736 135204
rect 328788 135192 328794 135244
rect 347958 135192 347964 135244
rect 348016 135232 348022 135244
rect 348142 135232 348148 135244
rect 348016 135204 348148 135232
rect 348016 135192 348022 135204
rect 348142 135192 348148 135204
rect 348200 135192 348206 135244
rect 234801 134623 234859 134629
rect 234801 134589 234813 134623
rect 234847 134620 234859 134623
rect 234982 134620 234988 134632
rect 234847 134592 234988 134620
rect 234847 134589 234859 134592
rect 234801 134583 234859 134589
rect 234982 134580 234988 134592
rect 235040 134580 235046 134632
rect 309502 134512 309508 134564
rect 309560 134552 309566 134564
rect 309686 134552 309692 134564
rect 309560 134524 309692 134552
rect 309560 134512 309566 134524
rect 309686 134512 309692 134524
rect 309744 134512 309750 134564
rect 269114 134104 269120 134156
rect 269172 134144 269178 134156
rect 275370 134144 275376 134156
rect 269172 134116 275376 134144
rect 269172 134104 269178 134116
rect 275370 134104 275376 134116
rect 275428 134104 275434 134156
rect 357434 134036 357440 134088
rect 357492 134076 357498 134088
rect 361114 134076 361120 134088
rect 357492 134048 361120 134076
rect 357492 134036 357498 134048
rect 361114 134036 361120 134048
rect 361172 134036 361178 134088
rect 398466 134036 398472 134088
rect 398524 134076 398530 134088
rect 399018 134076 399024 134088
rect 398524 134048 399024 134076
rect 398524 134036 398530 134048
rect 399018 134036 399024 134048
rect 399076 134036 399082 134088
rect 417878 134036 417884 134088
rect 417936 134076 417942 134088
rect 418338 134076 418344 134088
rect 417936 134048 418344 134076
rect 417936 134036 417942 134048
rect 418338 134036 418344 134048
rect 418396 134036 418402 134088
rect 317506 133968 317512 134020
rect 317564 134008 317570 134020
rect 326890 134008 326896 134020
rect 317564 133980 326896 134008
rect 317564 133968 317570 133980
rect 326890 133968 326896 133980
rect 326948 133968 326954 134020
rect 251174 133900 251180 133952
rect 251232 133940 251238 133952
rect 260742 133940 260748 133952
rect 251232 133912 260748 133940
rect 251232 133900 251238 133912
rect 260742 133900 260748 133912
rect 260800 133900 260806 133952
rect 308122 133900 308128 133952
rect 308180 133940 308186 133952
rect 308214 133940 308220 133952
rect 308180 133912 308220 133940
rect 308180 133900 308186 133912
rect 308214 133900 308220 133912
rect 308272 133900 308278 133952
rect 327258 133900 327264 133952
rect 327316 133940 327322 133952
rect 336642 133940 336648 133952
rect 327316 133912 336648 133940
rect 327316 133900 327322 133912
rect 336642 133900 336648 133912
rect 336700 133900 336706 133952
rect 251453 133875 251511 133881
rect 251453 133841 251465 133875
rect 251499 133872 251511 133875
rect 251542 133872 251548 133884
rect 251499 133844 251548 133872
rect 251499 133841 251511 133844
rect 251453 133835 251511 133841
rect 251542 133832 251548 133844
rect 251600 133832 251606 133884
rect 287330 133832 287336 133884
rect 287388 133872 287394 133884
rect 287514 133872 287520 133884
rect 287388 133844 287520 133872
rect 287388 133832 287394 133844
rect 287514 133832 287520 133844
rect 287572 133832 287578 133884
rect 310790 133872 310796 133884
rect 310751 133844 310796 133872
rect 310790 133832 310796 133844
rect 310848 133832 310854 133884
rect 233418 132512 233424 132524
rect 233379 132484 233424 132512
rect 233418 132472 233424 132484
rect 233476 132472 233482 132524
rect 239122 132512 239128 132524
rect 239083 132484 239128 132512
rect 239122 132472 239128 132484
rect 239180 132472 239186 132524
rect 240321 132515 240379 132521
rect 240321 132481 240333 132515
rect 240367 132512 240379 132515
rect 240410 132512 240416 132524
rect 240367 132484 240416 132512
rect 240367 132481 240379 132484
rect 240321 132475 240379 132481
rect 240410 132472 240416 132484
rect 240468 132472 240474 132524
rect 316310 132512 316316 132524
rect 316271 132484 316316 132512
rect 316310 132472 316316 132484
rect 316368 132472 316374 132524
rect 305362 132444 305368 132456
rect 305323 132416 305368 132444
rect 305362 132404 305368 132416
rect 305420 132404 305426 132456
rect 233418 131152 233424 131164
rect 233379 131124 233424 131152
rect 233418 131112 233424 131124
rect 233476 131112 233482 131164
rect 324590 131044 324596 131096
rect 324648 131084 324654 131096
rect 324866 131084 324872 131096
rect 324648 131056 324872 131084
rect 324648 131044 324654 131056
rect 324866 131044 324872 131056
rect 324924 131044 324930 131096
rect 255498 130432 255504 130484
rect 255556 130472 255562 130484
rect 255774 130472 255780 130484
rect 255556 130444 255780 130472
rect 255556 130432 255562 130444
rect 255774 130432 255780 130444
rect 255832 130432 255838 130484
rect 262677 129795 262735 129801
rect 262677 129761 262689 129795
rect 262723 129792 262735 129795
rect 262858 129792 262864 129804
rect 262723 129764 262864 129792
rect 262723 129761 262735 129764
rect 262677 129755 262735 129761
rect 262858 129752 262864 129764
rect 262916 129752 262922 129804
rect 235074 128364 235080 128376
rect 235035 128336 235080 128364
rect 235074 128324 235080 128336
rect 235132 128324 235138 128376
rect 238754 128256 238760 128308
rect 238812 128296 238818 128308
rect 238938 128296 238944 128308
rect 238812 128268 238944 128296
rect 238812 128256 238818 128268
rect 238938 128256 238944 128268
rect 238996 128256 239002 128308
rect 267090 128296 267096 128308
rect 267051 128268 267096 128296
rect 267090 128256 267096 128268
rect 267148 128256 267154 128308
rect 327350 128296 327356 128308
rect 327311 128268 327356 128296
rect 327350 128256 327356 128268
rect 327408 128256 327414 128308
rect 444098 128296 444104 128308
rect 444059 128268 444104 128296
rect 444098 128256 444104 128268
rect 444156 128256 444162 128308
rect 241882 125644 241888 125656
rect 241843 125616 241888 125644
rect 241882 125604 241888 125616
rect 241940 125604 241946 125656
rect 345198 125604 345204 125656
rect 345256 125644 345262 125656
rect 345382 125644 345388 125656
rect 345256 125616 345388 125644
rect 345256 125604 345262 125616
rect 345382 125604 345388 125616
rect 345440 125604 345446 125656
rect 254210 125576 254216 125588
rect 254171 125548 254216 125576
rect 254210 125536 254216 125548
rect 254268 125536 254274 125588
rect 328454 125536 328460 125588
rect 328512 125576 328518 125588
rect 347958 125576 347964 125588
rect 328512 125548 328557 125576
rect 347919 125548 347964 125576
rect 328512 125536 328518 125548
rect 347958 125536 347964 125548
rect 348016 125536 348022 125588
rect 435358 125536 435364 125588
rect 435416 125576 435422 125588
rect 435542 125576 435548 125588
rect 435416 125548 435548 125576
rect 435416 125536 435422 125548
rect 435542 125536 435548 125548
rect 435600 125536 435606 125588
rect 444098 125536 444104 125588
rect 444156 125576 444162 125588
rect 444193 125579 444251 125585
rect 444193 125576 444205 125579
rect 444156 125548 444205 125576
rect 444156 125536 444162 125548
rect 444193 125545 444205 125548
rect 444239 125545 444251 125579
rect 444193 125539 444251 125545
rect 233418 125508 233424 125520
rect 233379 125480 233424 125508
rect 233418 125468 233424 125480
rect 233476 125468 233482 125520
rect 316310 124284 316316 124296
rect 316236 124256 316316 124284
rect 316236 124228 316264 124256
rect 316310 124244 316316 124256
rect 316368 124244 316374 124296
rect 251450 124216 251456 124228
rect 251411 124188 251456 124216
rect 251450 124176 251456 124188
rect 251508 124176 251514 124228
rect 291562 124216 291568 124228
rect 291523 124188 291568 124216
rect 291562 124176 291568 124188
rect 291620 124176 291626 124228
rect 310790 124216 310796 124228
rect 310751 124188 310796 124216
rect 310790 124176 310796 124188
rect 310848 124176 310854 124228
rect 316218 124176 316224 124228
rect 316276 124176 316282 124228
rect 241882 124148 241888 124160
rect 241843 124120 241888 124148
rect 241882 124108 241888 124120
rect 241940 124108 241946 124160
rect 261205 124151 261263 124157
rect 261205 124117 261217 124151
rect 261251 124148 261263 124151
rect 261294 124148 261300 124160
rect 261251 124120 261300 124148
rect 261251 124117 261263 124120
rect 261205 124111 261263 124117
rect 261294 124108 261300 124120
rect 261352 124108 261358 124160
rect 287238 124108 287244 124160
rect 287296 124108 287302 124160
rect 345198 124148 345204 124160
rect 345159 124120 345204 124148
rect 345198 124108 345204 124120
rect 345256 124108 345262 124160
rect 287256 124080 287284 124108
rect 287422 124080 287428 124092
rect 287256 124052 287428 124080
rect 287422 124040 287428 124052
rect 287480 124040 287486 124092
rect 252830 123604 252836 123616
rect 252756 123576 252836 123604
rect 252756 123548 252784 123576
rect 252830 123564 252836 123576
rect 252888 123564 252894 123616
rect 252738 123496 252744 123548
rect 252796 123496 252802 123548
rect 235074 122856 235080 122868
rect 235035 122828 235080 122856
rect 235074 122816 235080 122828
rect 235132 122816 235138 122868
rect 305362 122856 305368 122868
rect 305323 122828 305368 122856
rect 305362 122816 305368 122828
rect 305420 122816 305426 122868
rect 240321 122791 240379 122797
rect 240321 122757 240333 122791
rect 240367 122788 240379 122791
rect 240410 122788 240416 122800
rect 240367 122760 240416 122788
rect 240367 122757 240379 122760
rect 240321 122751 240379 122757
rect 240410 122748 240416 122760
rect 240468 122748 240474 122800
rect 2774 122068 2780 122120
rect 2832 122108 2838 122120
rect 4798 122108 4804 122120
rect 2832 122080 4804 122108
rect 2832 122068 2838 122080
rect 4798 122068 4804 122080
rect 4856 122068 4862 122120
rect 233418 121496 233424 121508
rect 233379 121468 233424 121496
rect 233418 121456 233424 121468
rect 233476 121456 233482 121508
rect 291562 121496 291568 121508
rect 291523 121468 291568 121496
rect 291562 121456 291568 121468
rect 291620 121456 291626 121508
rect 309410 120096 309416 120148
rect 309468 120136 309474 120148
rect 309686 120136 309692 120148
rect 309468 120108 309692 120136
rect 309468 120096 309474 120108
rect 309686 120096 309692 120108
rect 309744 120096 309750 120148
rect 234890 120068 234896 120080
rect 234851 120040 234896 120068
rect 234890 120028 234896 120040
rect 234948 120028 234954 120080
rect 262677 120071 262735 120077
rect 262677 120037 262689 120071
rect 262723 120068 262735 120071
rect 262858 120068 262864 120080
rect 262723 120040 262864 120068
rect 262723 120037 262735 120040
rect 262677 120031 262735 120037
rect 262858 120028 262864 120040
rect 262916 120028 262922 120080
rect 292850 118736 292856 118788
rect 292908 118736 292914 118788
rect 304994 118736 305000 118788
rect 305052 118776 305058 118788
rect 305362 118776 305368 118788
rect 305052 118748 305368 118776
rect 305052 118736 305058 118748
rect 305362 118736 305368 118748
rect 305420 118736 305426 118788
rect 229278 118668 229284 118720
rect 229336 118668 229342 118720
rect 266998 118668 267004 118720
rect 267056 118708 267062 118720
rect 267182 118708 267188 118720
rect 267056 118680 267188 118708
rect 267056 118668 267062 118680
rect 267182 118668 267188 118680
rect 267240 118668 267246 118720
rect 280522 118668 280528 118720
rect 280580 118668 280586 118720
rect 229296 118640 229324 118668
rect 229370 118640 229376 118652
rect 229296 118612 229376 118640
rect 229370 118600 229376 118612
rect 229428 118600 229434 118652
rect 261202 118640 261208 118652
rect 261163 118612 261208 118640
rect 261202 118600 261208 118612
rect 261260 118600 261266 118652
rect 280540 118640 280568 118668
rect 292868 118652 292896 118736
rect 280614 118640 280620 118652
rect 280540 118612 280620 118640
rect 280614 118600 280620 118612
rect 280672 118600 280678 118652
rect 292850 118600 292856 118652
rect 292908 118600 292914 118652
rect 328457 118643 328515 118649
rect 328457 118609 328469 118643
rect 328503 118640 328515 118643
rect 328546 118640 328552 118652
rect 328503 118612 328552 118640
rect 328503 118609 328515 118612
rect 328457 118603 328515 118609
rect 328546 118600 328552 118612
rect 328604 118600 328610 118652
rect 444190 118640 444196 118652
rect 444151 118612 444196 118640
rect 444190 118600 444196 118612
rect 444248 118600 444254 118652
rect 347958 116056 347964 116068
rect 347919 116028 347964 116056
rect 347958 116016 347964 116028
rect 348016 116016 348022 116068
rect 254210 115988 254216 116000
rect 254171 115960 254216 115988
rect 254210 115948 254216 115960
rect 254268 115948 254274 116000
rect 229281 115923 229339 115929
rect 229281 115889 229293 115923
rect 229327 115920 229339 115923
rect 229370 115920 229376 115932
rect 229327 115892 229376 115920
rect 229327 115889 229339 115892
rect 229281 115883 229339 115889
rect 229370 115880 229376 115892
rect 229428 115880 229434 115932
rect 245930 115920 245936 115932
rect 245891 115892 245936 115920
rect 245930 115880 245936 115892
rect 245988 115880 245994 115932
rect 266998 115880 267004 115932
rect 267056 115920 267062 115932
rect 267182 115920 267188 115932
rect 267056 115892 267188 115920
rect 267056 115880 267062 115892
rect 267182 115880 267188 115892
rect 267240 115880 267246 115932
rect 298462 115920 298468 115932
rect 298423 115892 298468 115920
rect 298462 115880 298468 115892
rect 298520 115880 298526 115932
rect 347958 115880 347964 115932
rect 348016 115920 348022 115932
rect 348142 115920 348148 115932
rect 348016 115892 348148 115920
rect 348016 115880 348022 115892
rect 348142 115880 348148 115892
rect 348200 115880 348206 115932
rect 309318 115240 309324 115252
rect 309279 115212 309324 115240
rect 309318 115200 309324 115212
rect 309376 115200 309382 115252
rect 310790 114588 310796 114640
rect 310848 114588 310854 114640
rect 241882 114560 241888 114572
rect 241843 114532 241888 114560
rect 241882 114520 241888 114532
rect 241940 114520 241946 114572
rect 234982 114452 234988 114504
rect 235040 114492 235046 114504
rect 235074 114492 235080 114504
rect 235040 114464 235080 114492
rect 235040 114452 235046 114464
rect 235074 114452 235080 114464
rect 235132 114452 235138 114504
rect 255590 114492 255596 114504
rect 255551 114464 255596 114492
rect 255590 114452 255596 114464
rect 255648 114452 255654 114504
rect 287330 114492 287336 114504
rect 287291 114464 287336 114492
rect 287330 114452 287336 114464
rect 287388 114452 287394 114504
rect 288710 114492 288716 114504
rect 288671 114464 288716 114492
rect 288710 114452 288716 114464
rect 288768 114452 288774 114504
rect 310808 114492 310836 114588
rect 316218 114520 316224 114572
rect 316276 114560 316282 114572
rect 316310 114560 316316 114572
rect 316276 114532 316316 114560
rect 316276 114520 316282 114532
rect 316310 114520 316316 114532
rect 316368 114520 316374 114572
rect 345198 114560 345204 114572
rect 345159 114532 345204 114560
rect 345198 114520 345204 114532
rect 345256 114520 345262 114572
rect 310882 114492 310888 114504
rect 310808 114464 310888 114492
rect 310882 114452 310888 114464
rect 310940 114452 310946 114504
rect 342530 114492 342536 114504
rect 342491 114464 342536 114492
rect 342530 114452 342536 114464
rect 342588 114452 342594 114504
rect 313642 113132 313648 113144
rect 313603 113104 313648 113132
rect 313642 113092 313648 113104
rect 313700 113092 313706 113144
rect 241606 111052 241612 111104
rect 241664 111092 241670 111104
rect 241882 111092 241888 111104
rect 241664 111064 241888 111092
rect 241664 111052 241670 111064
rect 241882 111052 241888 111064
rect 241940 111052 241946 111104
rect 239122 109080 239128 109132
rect 239180 109080 239186 109132
rect 238754 109012 238760 109064
rect 238812 109052 238818 109064
rect 238938 109052 238944 109064
rect 238812 109024 238944 109052
rect 238812 109012 238818 109024
rect 238938 109012 238944 109024
rect 238996 109012 239002 109064
rect 238938 108876 238944 108928
rect 238996 108916 239002 108928
rect 239140 108916 239168 109080
rect 280430 109012 280436 109064
rect 280488 109052 280494 109064
rect 280614 109052 280620 109064
rect 280488 109024 280620 109052
rect 280488 109012 280494 109024
rect 280614 109012 280620 109024
rect 280672 109012 280678 109064
rect 434346 109012 434352 109064
rect 434404 109012 434410 109064
rect 435358 109012 435364 109064
rect 435416 109052 435422 109064
rect 435542 109052 435548 109064
rect 435416 109024 435548 109052
rect 435416 109012 435422 109024
rect 435542 109012 435548 109024
rect 435600 109012 435606 109064
rect 444006 109012 444012 109064
rect 444064 109052 444070 109064
rect 444190 109052 444196 109064
rect 444064 109024 444196 109052
rect 444064 109012 444070 109024
rect 444190 109012 444196 109024
rect 444248 109012 444254 109064
rect 434364 108984 434392 109012
rect 434438 108984 434444 108996
rect 434364 108956 434444 108984
rect 434438 108944 434444 108956
rect 434496 108944 434502 108996
rect 238996 108888 239168 108916
rect 238996 108876 239002 108888
rect 298465 108851 298523 108857
rect 298465 108817 298477 108851
rect 298511 108848 298523 108851
rect 298554 108848 298560 108860
rect 298511 108820 298560 108848
rect 298511 108817 298523 108820
rect 298465 108811 298523 108817
rect 298554 108808 298560 108820
rect 298612 108808 298618 108860
rect 229278 106332 229284 106344
rect 229239 106304 229284 106332
rect 229278 106292 229284 106304
rect 229336 106292 229342 106344
rect 245930 106332 245936 106344
rect 245891 106304 245936 106332
rect 245930 106292 245936 106304
rect 245988 106292 245994 106344
rect 324682 106332 324688 106344
rect 324643 106304 324688 106332
rect 324682 106292 324688 106304
rect 324740 106292 324746 106344
rect 305270 106264 305276 106276
rect 305231 106236 305276 106264
rect 305270 106224 305276 106236
rect 305328 106224 305334 106276
rect 347958 106264 347964 106276
rect 347919 106236 347964 106264
rect 347958 106224 347964 106236
rect 348016 106224 348022 106276
rect 444098 106264 444104 106276
rect 444059 106236 444104 106264
rect 444098 106224 444104 106236
rect 444156 106224 444162 106276
rect 342530 104972 342536 104984
rect 342491 104944 342536 104972
rect 342530 104932 342536 104944
rect 342588 104932 342594 104984
rect 240318 104904 240324 104916
rect 240279 104876 240324 104904
rect 240318 104864 240324 104876
rect 240376 104864 240382 104916
rect 255590 104904 255596 104916
rect 255551 104876 255596 104904
rect 255590 104864 255596 104876
rect 255648 104864 255654 104916
rect 287330 104904 287336 104916
rect 287291 104876 287336 104904
rect 287330 104864 287336 104876
rect 287388 104864 287394 104916
rect 288713 104907 288771 104913
rect 288713 104873 288725 104907
rect 288759 104904 288771 104907
rect 288802 104904 288808 104916
rect 288759 104876 288808 104904
rect 288759 104873 288771 104876
rect 288713 104867 288771 104873
rect 288802 104864 288808 104876
rect 288860 104864 288866 104916
rect 324682 104904 324688 104916
rect 324643 104876 324688 104904
rect 324682 104864 324688 104876
rect 324740 104864 324746 104916
rect 234982 104796 234988 104848
rect 235040 104836 235046 104848
rect 235074 104836 235080 104848
rect 235040 104808 235080 104836
rect 235040 104796 235046 104808
rect 235074 104796 235080 104808
rect 235132 104796 235138 104848
rect 241790 104836 241796 104848
rect 241751 104808 241796 104836
rect 241790 104796 241796 104808
rect 241848 104796 241854 104848
rect 251450 104836 251456 104848
rect 251411 104808 251456 104836
rect 251450 104796 251456 104808
rect 251508 104796 251514 104848
rect 280522 104836 280528 104848
rect 280483 104808 280528 104836
rect 280522 104796 280528 104808
rect 280580 104796 280586 104848
rect 327353 104839 327411 104845
rect 327353 104805 327365 104839
rect 327399 104836 327411 104839
rect 327442 104836 327448 104848
rect 327399 104808 327448 104836
rect 327399 104805 327411 104808
rect 327353 104799 327411 104805
rect 327442 104796 327448 104808
rect 327500 104796 327506 104848
rect 342530 104836 342536 104848
rect 342491 104808 342536 104836
rect 342530 104796 342536 104808
rect 342588 104796 342594 104848
rect 345198 104836 345204 104848
rect 345159 104808 345204 104836
rect 345198 104796 345204 104808
rect 345256 104796 345262 104848
rect 434349 104839 434407 104845
rect 434349 104805 434361 104839
rect 434395 104836 434407 104839
rect 434438 104836 434444 104848
rect 434395 104808 434444 104836
rect 434395 104805 434407 104808
rect 434349 104799 434407 104805
rect 434438 104796 434444 104808
rect 434496 104796 434502 104848
rect 305086 103572 305092 103624
rect 305144 103572 305150 103624
rect 305104 103488 305132 103572
rect 305086 103436 305092 103488
rect 305144 103436 305150 103488
rect 308030 103436 308036 103488
rect 308088 103476 308094 103488
rect 308122 103476 308128 103488
rect 308088 103448 308128 103476
rect 308088 103436 308094 103448
rect 308122 103436 308128 103448
rect 308180 103436 308186 103488
rect 310882 103436 310888 103488
rect 310940 103476 310946 103488
rect 311066 103476 311072 103488
rect 310940 103448 311072 103476
rect 310940 103436 310946 103448
rect 311066 103436 311072 103448
rect 311124 103436 311130 103488
rect 309318 102456 309324 102468
rect 309279 102428 309324 102456
rect 309318 102416 309324 102428
rect 309376 102416 309382 102468
rect 313458 102416 313464 102468
rect 313516 102456 313522 102468
rect 313645 102459 313703 102465
rect 313645 102456 313657 102459
rect 313516 102428 313657 102456
rect 313516 102416 313522 102428
rect 313645 102425 313657 102428
rect 313691 102425 313703 102459
rect 313645 102419 313703 102425
rect 262674 102184 262680 102196
rect 262635 102156 262680 102184
rect 262674 102144 262680 102156
rect 262732 102144 262738 102196
rect 305270 102184 305276 102196
rect 305231 102156 305276 102184
rect 305270 102144 305276 102156
rect 305328 102144 305334 102196
rect 267001 102119 267059 102125
rect 267001 102085 267013 102119
rect 267047 102116 267059 102119
rect 267090 102116 267096 102128
rect 267047 102088 267096 102116
rect 267047 102085 267059 102088
rect 267001 102079 267059 102085
rect 267090 102076 267096 102088
rect 267148 102076 267154 102128
rect 234801 100759 234859 100765
rect 234801 100725 234813 100759
rect 234847 100756 234859 100759
rect 234893 100759 234951 100765
rect 234893 100756 234905 100759
rect 234847 100728 234905 100756
rect 234847 100725 234859 100728
rect 234801 100719 234859 100725
rect 234893 100725 234905 100728
rect 234939 100725 234951 100759
rect 234893 100719 234951 100725
rect 238938 100036 238944 100088
rect 238996 100076 239002 100088
rect 239122 100076 239128 100088
rect 238996 100048 239128 100076
rect 238996 100036 239002 100048
rect 239122 100036 239128 100048
rect 239180 100036 239186 100088
rect 262493 99467 262551 99473
rect 262493 99433 262505 99467
rect 262539 99464 262551 99467
rect 262674 99464 262680 99476
rect 262539 99436 262680 99464
rect 262539 99433 262551 99436
rect 262493 99427 262551 99433
rect 262674 99424 262680 99436
rect 262732 99424 262738 99476
rect 288621 99467 288679 99473
rect 288621 99433 288633 99467
rect 288667 99464 288679 99467
rect 288802 99464 288808 99476
rect 288667 99436 288808 99464
rect 288667 99433 288679 99436
rect 288621 99427 288679 99433
rect 288802 99424 288808 99436
rect 288860 99424 288866 99476
rect 290090 99424 290096 99476
rect 290148 99424 290154 99476
rect 298554 99464 298560 99476
rect 298480 99436 298560 99464
rect 229278 99356 229284 99408
rect 229336 99356 229342 99408
rect 229296 99328 229324 99356
rect 290108 99340 290136 99424
rect 298480 99340 298508 99436
rect 298554 99424 298560 99436
rect 298612 99424 298618 99476
rect 324682 99464 324688 99476
rect 324608 99436 324688 99464
rect 324608 99340 324636 99436
rect 324682 99424 324688 99436
rect 324740 99424 324746 99476
rect 229370 99328 229376 99340
rect 229296 99300 229376 99328
rect 229370 99288 229376 99300
rect 229428 99288 229434 99340
rect 290090 99288 290096 99340
rect 290148 99288 290154 99340
rect 298462 99288 298468 99340
rect 298520 99288 298526 99340
rect 324590 99288 324596 99340
rect 324648 99288 324654 99340
rect 444098 99328 444104 99340
rect 444059 99300 444104 99328
rect 444098 99288 444104 99300
rect 444156 99288 444162 99340
rect 255590 98676 255596 98728
rect 255648 98716 255654 98728
rect 255685 98719 255743 98725
rect 255685 98716 255697 98719
rect 255648 98688 255697 98716
rect 255648 98676 255654 98688
rect 255685 98685 255697 98688
rect 255731 98685 255743 98719
rect 255685 98679 255743 98685
rect 345201 98719 345259 98725
rect 345201 98685 345213 98719
rect 345247 98716 345259 98719
rect 345382 98716 345388 98728
rect 345247 98688 345388 98716
rect 345247 98685 345259 98688
rect 345201 98679 345259 98685
rect 345382 98676 345388 98688
rect 345440 98676 345446 98728
rect 347958 96744 347964 96756
rect 347919 96716 347964 96744
rect 347958 96704 347964 96716
rect 348016 96704 348022 96756
rect 229281 96611 229339 96617
rect 229281 96577 229293 96611
rect 229327 96608 229339 96611
rect 229370 96608 229376 96620
rect 229327 96580 229376 96608
rect 229327 96577 229339 96580
rect 229281 96571 229339 96577
rect 229370 96568 229376 96580
rect 229428 96568 229434 96620
rect 347958 96568 347964 96620
rect 348016 96608 348022 96620
rect 348050 96608 348056 96620
rect 348016 96580 348056 96608
rect 348016 96568 348022 96580
rect 348050 96568 348056 96580
rect 348108 96568 348114 96620
rect 251450 95316 251456 95328
rect 251411 95288 251456 95316
rect 251450 95276 251456 95288
rect 251508 95276 251514 95328
rect 241793 95251 241851 95257
rect 241793 95217 241805 95251
rect 241839 95248 241851 95251
rect 241882 95248 241888 95260
rect 241839 95220 241888 95248
rect 241839 95217 241851 95220
rect 241793 95211 241851 95217
rect 241882 95208 241888 95220
rect 241940 95208 241946 95260
rect 280525 95251 280583 95257
rect 280525 95217 280537 95251
rect 280571 95248 280583 95251
rect 280614 95248 280620 95260
rect 280571 95220 280620 95248
rect 280571 95217 280583 95220
rect 280525 95211 280583 95217
rect 280614 95208 280620 95220
rect 280672 95208 280678 95260
rect 327350 95248 327356 95260
rect 327311 95220 327356 95248
rect 327350 95208 327356 95220
rect 327408 95208 327414 95260
rect 342530 95248 342536 95260
rect 342491 95220 342536 95248
rect 342530 95208 342536 95220
rect 342588 95208 342594 95260
rect 434346 95248 434352 95260
rect 434307 95220 434352 95248
rect 434346 95208 434352 95220
rect 434404 95208 434410 95260
rect 240410 95140 240416 95192
rect 240468 95180 240474 95192
rect 240502 95180 240508 95192
rect 240468 95152 240508 95180
rect 240468 95140 240474 95152
rect 240502 95140 240508 95152
rect 240560 95140 240566 95192
rect 251174 95140 251180 95192
rect 251232 95180 251238 95192
rect 251450 95180 251456 95192
rect 251232 95152 251456 95180
rect 251232 95140 251238 95152
rect 251450 95140 251456 95152
rect 251508 95140 251514 95192
rect 244458 94636 244464 94648
rect 244419 94608 244464 94636
rect 244458 94596 244464 94608
rect 244516 94596 244522 94648
rect 248690 94636 248696 94648
rect 248651 94608 248696 94636
rect 248690 94596 248696 94608
rect 248748 94596 248754 94648
rect 255682 93848 255688 93900
rect 255740 93888 255746 93900
rect 255740 93860 255785 93888
rect 255740 93848 255746 93860
rect 240502 93820 240508 93832
rect 240463 93792 240508 93820
rect 240502 93780 240508 93792
rect 240560 93780 240566 93832
rect 345201 93823 345259 93829
rect 345201 93789 345213 93823
rect 345247 93820 345259 93823
rect 345382 93820 345388 93832
rect 345247 93792 345388 93820
rect 345247 93789 345259 93792
rect 345201 93783 345259 93789
rect 345382 93780 345388 93792
rect 345440 93780 345446 93832
rect 255682 93752 255688 93764
rect 255643 93724 255688 93752
rect 255682 93712 255688 93724
rect 255740 93712 255746 93764
rect 234798 92052 234804 92064
rect 234759 92024 234804 92052
rect 234798 92012 234804 92024
rect 234856 92012 234862 92064
rect 434346 91780 434352 91792
rect 434307 91752 434352 91780
rect 434346 91740 434352 91752
rect 434404 91740 434410 91792
rect 309410 89808 309416 89820
rect 309371 89780 309416 89808
rect 309410 89768 309416 89780
rect 309468 89768 309474 89820
rect 233326 89700 233332 89752
rect 233384 89740 233390 89752
rect 233510 89740 233516 89752
rect 233384 89712 233516 89740
rect 233384 89700 233390 89712
rect 233510 89700 233516 89712
rect 233568 89700 233574 89752
rect 280430 89700 280436 89752
rect 280488 89740 280494 89752
rect 280614 89740 280620 89752
rect 280488 89712 280620 89740
rect 280488 89700 280494 89712
rect 280614 89700 280620 89712
rect 280672 89700 280678 89752
rect 444006 89700 444012 89752
rect 444064 89740 444070 89752
rect 444190 89740 444196 89752
rect 444064 89712 444196 89740
rect 444064 89700 444070 89712
rect 444190 89700 444196 89712
rect 444248 89700 444254 89752
rect 434622 87320 434628 87372
rect 434680 87320 434686 87372
rect 282822 87184 282828 87236
rect 282880 87224 282886 87236
rect 292758 87224 292764 87236
rect 282880 87196 292764 87224
rect 282880 87184 282886 87196
rect 292758 87184 292764 87196
rect 292816 87184 292822 87236
rect 434640 87168 434668 87320
rect 356054 87116 356060 87168
rect 356112 87156 356118 87168
rect 365622 87156 365628 87168
rect 356112 87128 365628 87156
rect 356112 87116 356118 87128
rect 365622 87116 365628 87128
rect 365680 87116 365686 87168
rect 417878 87116 417884 87168
rect 417936 87156 417942 87168
rect 418338 87156 418344 87168
rect 417936 87128 418344 87156
rect 417936 87116 417942 87128
rect 418338 87116 418344 87128
rect 418396 87116 418402 87168
rect 434349 87159 434407 87165
rect 434349 87125 434361 87159
rect 434395 87156 434407 87159
rect 434530 87156 434536 87168
rect 434395 87128 434536 87156
rect 434395 87125 434407 87128
rect 434349 87119 434407 87125
rect 434530 87116 434536 87128
rect 434588 87116 434594 87168
rect 434622 87116 434628 87168
rect 434680 87116 434686 87168
rect 398466 87048 398472 87100
rect 398524 87088 398530 87100
rect 398834 87088 398840 87100
rect 398524 87060 398840 87088
rect 398524 87048 398530 87060
rect 398834 87048 398840 87060
rect 398892 87048 398898 87100
rect 229278 87020 229284 87032
rect 229239 86992 229284 87020
rect 229278 86980 229284 86992
rect 229336 86980 229342 87032
rect 305546 87020 305552 87032
rect 305472 86992 305552 87020
rect 305472 86964 305500 86992
rect 305546 86980 305552 86992
rect 305604 86980 305610 87032
rect 444374 86980 444380 87032
rect 444432 87020 444438 87032
rect 449250 87020 449256 87032
rect 444432 86992 449256 87020
rect 444432 86980 444438 86992
rect 449250 86980 449256 86992
rect 449308 86980 449314 87032
rect 463786 86980 463792 87032
rect 463844 87020 463850 87032
rect 466546 87020 466552 87032
rect 463844 86992 466552 87020
rect 463844 86980 463850 86992
rect 466546 86980 466552 86992
rect 466604 86980 466610 87032
rect 262490 86952 262496 86964
rect 262451 86924 262496 86952
rect 262490 86912 262496 86924
rect 262548 86912 262554 86964
rect 298462 86912 298468 86964
rect 298520 86952 298526 86964
rect 298554 86952 298560 86964
rect 298520 86924 298560 86952
rect 298520 86912 298526 86924
rect 298554 86912 298560 86924
rect 298612 86912 298618 86964
rect 305454 86912 305460 86964
rect 305512 86912 305518 86964
rect 343726 86912 343732 86964
rect 343784 86952 343790 86964
rect 343818 86952 343824 86964
rect 343784 86924 343824 86952
rect 343784 86912 343790 86924
rect 343818 86912 343824 86924
rect 343876 86912 343882 86964
rect 362957 86955 363015 86961
rect 362957 86921 362969 86955
rect 363003 86952 363015 86955
rect 363046 86952 363052 86964
rect 363003 86924 363052 86952
rect 363003 86921 363015 86924
rect 362957 86915 363015 86921
rect 363046 86912 363052 86924
rect 363104 86912 363110 86964
rect 444098 86952 444104 86964
rect 444059 86924 444104 86952
rect 444098 86912 444104 86924
rect 444156 86912 444162 86964
rect 327350 86884 327356 86896
rect 327311 86856 327356 86884
rect 327350 86844 327356 86856
rect 327408 86844 327414 86896
rect 288618 86136 288624 86148
rect 288579 86108 288624 86136
rect 288618 86096 288624 86108
rect 288676 86096 288682 86148
rect 244458 85592 244464 85604
rect 244419 85564 244464 85592
rect 244458 85552 244464 85564
rect 244516 85552 244522 85604
rect 248693 85595 248751 85601
rect 248693 85561 248705 85595
rect 248739 85592 248751 85595
rect 248782 85592 248788 85604
rect 248739 85564 248788 85592
rect 248739 85561 248751 85564
rect 248693 85555 248751 85561
rect 248782 85552 248788 85564
rect 248840 85552 248846 85604
rect 287330 85552 287336 85604
rect 287388 85592 287394 85604
rect 287422 85592 287428 85604
rect 287388 85564 287428 85592
rect 287388 85552 287394 85564
rect 287422 85552 287428 85564
rect 287480 85552 287486 85604
rect 309410 85592 309416 85604
rect 309371 85564 309416 85592
rect 309410 85552 309416 85564
rect 309468 85552 309474 85604
rect 313458 85552 313464 85604
rect 313516 85592 313522 85604
rect 313642 85592 313648 85604
rect 313516 85564 313648 85592
rect 313516 85552 313522 85564
rect 313642 85552 313648 85564
rect 313700 85552 313706 85604
rect 343726 85524 343732 85536
rect 343687 85496 343732 85524
rect 343726 85484 343732 85496
rect 343784 85484 343790 85536
rect 435174 85524 435180 85536
rect 435135 85496 435180 85524
rect 435174 85484 435180 85496
rect 435232 85484 435238 85536
rect 240410 84192 240416 84244
rect 240468 84232 240474 84244
rect 240505 84235 240563 84241
rect 240505 84232 240517 84235
rect 240468 84204 240517 84232
rect 240468 84192 240474 84204
rect 240505 84201 240517 84204
rect 240551 84201 240563 84235
rect 240505 84195 240563 84201
rect 255685 84235 255743 84241
rect 255685 84201 255697 84235
rect 255731 84232 255743 84235
rect 255774 84232 255780 84244
rect 255731 84204 255780 84232
rect 255731 84201 255743 84204
rect 255685 84195 255743 84201
rect 255774 84192 255780 84204
rect 255832 84192 255838 84244
rect 291470 84192 291476 84244
rect 291528 84232 291534 84244
rect 291562 84232 291568 84244
rect 291528 84204 291568 84232
rect 291528 84192 291534 84204
rect 291562 84192 291568 84204
rect 291620 84192 291626 84244
rect 234798 84164 234804 84176
rect 234759 84136 234804 84164
rect 234798 84124 234804 84136
rect 234856 84124 234862 84176
rect 307938 84164 307944 84176
rect 307899 84136 307944 84164
rect 307938 84124 307944 84136
rect 307996 84124 308002 84176
rect 313642 84164 313648 84176
rect 313603 84136 313648 84164
rect 313642 84124 313648 84136
rect 313700 84124 313706 84176
rect 267001 82875 267059 82881
rect 267001 82841 267013 82875
rect 267047 82872 267059 82875
rect 267090 82872 267096 82884
rect 267047 82844 267096 82872
rect 267047 82841 267059 82844
rect 267001 82835 267059 82841
rect 267090 82832 267096 82844
rect 267148 82832 267154 82884
rect 324590 82356 324596 82408
rect 324648 82356 324654 82408
rect 324608 82272 324636 82356
rect 324590 82220 324596 82272
rect 324648 82220 324654 82272
rect 287330 80112 287336 80164
rect 287388 80112 287394 80164
rect 342530 80112 342536 80164
rect 342588 80112 342594 80164
rect 229278 80044 229284 80096
rect 229336 80044 229342 80096
rect 254210 80044 254216 80096
rect 254268 80044 254274 80096
rect 229296 79948 229324 80044
rect 254228 79960 254256 80044
rect 287348 80028 287376 80112
rect 299842 80044 299848 80096
rect 299900 80044 299906 80096
rect 325970 80044 325976 80096
rect 326028 80044 326034 80096
rect 287330 79976 287336 80028
rect 287388 79976 287394 80028
rect 299860 79960 299888 80044
rect 325988 79960 326016 80044
rect 342548 80028 342576 80112
rect 342530 79976 342536 80028
rect 342588 79976 342594 80028
rect 229370 79948 229376 79960
rect 229296 79920 229376 79948
rect 229370 79908 229376 79920
rect 229428 79908 229434 79960
rect 254210 79908 254216 79960
rect 254268 79908 254274 79960
rect 299842 79908 299848 79960
rect 299900 79908 299906 79960
rect 325970 79908 325976 79960
rect 326028 79908 326034 79960
rect 2774 79432 2780 79484
rect 2832 79472 2838 79484
rect 6178 79472 6184 79484
rect 2832 79444 6184 79472
rect 2832 79432 2838 79444
rect 6178 79432 6184 79444
rect 6236 79432 6242 79484
rect 291473 79339 291531 79345
rect 291473 79305 291485 79339
rect 291519 79336 291531 79339
rect 291562 79336 291568 79348
rect 291519 79308 291568 79336
rect 291519 79305 291531 79308
rect 291473 79299 291531 79305
rect 291562 79296 291568 79308
rect 291620 79296 291626 79348
rect 267090 77976 267096 77988
rect 267051 77948 267096 77976
rect 267090 77936 267096 77948
rect 267148 77936 267154 77988
rect 255590 77528 255596 77580
rect 255648 77568 255654 77580
rect 255774 77568 255780 77580
rect 255648 77540 255780 77568
rect 255648 77528 255654 77540
rect 255774 77528 255780 77540
rect 255832 77528 255838 77580
rect 233418 77256 233424 77308
rect 233476 77296 233482 77308
rect 233510 77296 233516 77308
rect 233476 77268 233516 77296
rect 233476 77256 233482 77268
rect 233510 77256 233516 77268
rect 233568 77256 233574 77308
rect 234982 77256 234988 77308
rect 235040 77296 235046 77308
rect 235074 77296 235080 77308
rect 235040 77268 235080 77296
rect 235040 77256 235046 77268
rect 235074 77256 235080 77268
rect 235132 77256 235138 77308
rect 244458 77256 244464 77308
rect 244516 77296 244522 77308
rect 244550 77296 244556 77308
rect 244516 77268 244556 77296
rect 244516 77256 244522 77268
rect 244550 77256 244556 77268
rect 244608 77256 244614 77308
rect 327350 77296 327356 77308
rect 327311 77268 327356 77296
rect 327350 77256 327356 77268
rect 327408 77256 327414 77308
rect 362954 77296 362960 77308
rect 362915 77268 362960 77296
rect 362954 77256 362960 77268
rect 363012 77256 363018 77308
rect 444101 77299 444159 77305
rect 444101 77265 444113 77299
rect 444147 77296 444159 77299
rect 444190 77296 444196 77308
rect 444147 77268 444196 77296
rect 444147 77265 444159 77268
rect 444101 77259 444159 77265
rect 444190 77256 444196 77268
rect 444248 77256 444254 77308
rect 261110 77188 261116 77240
rect 261168 77188 261174 77240
rect 262490 77188 262496 77240
rect 262548 77228 262554 77240
rect 262858 77228 262864 77240
rect 262548 77200 262864 77228
rect 262548 77188 262554 77200
rect 262858 77188 262864 77200
rect 262916 77188 262922 77240
rect 261128 77160 261156 77188
rect 261294 77160 261300 77172
rect 261128 77132 261300 77160
rect 261294 77120 261300 77132
rect 261352 77120 261358 77172
rect 362954 77160 362960 77172
rect 362915 77132 362960 77160
rect 362954 77120 362960 77132
rect 363012 77120 363018 77172
rect 343726 76004 343732 76016
rect 343687 75976 343732 76004
rect 343726 75964 343732 75976
rect 343784 75964 343790 76016
rect 290090 75896 290096 75948
rect 290148 75896 290154 75948
rect 345198 75936 345204 75948
rect 345159 75908 345204 75936
rect 345198 75896 345204 75908
rect 345256 75896 345262 75948
rect 435174 75936 435180 75948
rect 435135 75908 435180 75936
rect 435174 75896 435180 75908
rect 435232 75896 435238 75948
rect 240410 75828 240416 75880
rect 240468 75868 240474 75880
rect 240505 75871 240563 75877
rect 240505 75868 240517 75871
rect 240468 75840 240517 75868
rect 240468 75828 240474 75840
rect 240505 75837 240517 75840
rect 240551 75837 240563 75871
rect 240505 75831 240563 75837
rect 244458 75828 244464 75880
rect 244516 75868 244522 75880
rect 244550 75868 244556 75880
rect 244516 75840 244556 75868
rect 244516 75828 244522 75840
rect 244550 75828 244556 75840
rect 244608 75828 244614 75880
rect 248782 75868 248788 75880
rect 248743 75840 248788 75868
rect 248782 75828 248788 75840
rect 248840 75828 248846 75880
rect 262769 75871 262827 75877
rect 262769 75837 262781 75871
rect 262815 75868 262827 75871
rect 262858 75868 262864 75880
rect 262815 75840 262864 75868
rect 262815 75837 262827 75840
rect 262769 75831 262827 75837
rect 262858 75828 262864 75840
rect 262916 75828 262922 75880
rect 290108 75800 290136 75896
rect 343726 75868 343732 75880
rect 343687 75840 343732 75868
rect 343726 75828 343732 75840
rect 343784 75828 343790 75880
rect 434257 75871 434315 75877
rect 434257 75837 434269 75871
rect 434303 75868 434315 75871
rect 434346 75868 434352 75880
rect 434303 75840 434352 75868
rect 434303 75837 434315 75840
rect 434257 75831 434315 75837
rect 434346 75828 434352 75840
rect 434404 75828 434410 75880
rect 290182 75800 290188 75812
rect 290108 75772 290188 75800
rect 290182 75760 290188 75772
rect 290240 75760 290246 75812
rect 234798 74576 234804 74588
rect 234759 74548 234804 74576
rect 234798 74536 234804 74548
rect 234856 74536 234862 74588
rect 305270 74536 305276 74588
rect 305328 74576 305334 74588
rect 305454 74576 305460 74588
rect 305328 74548 305460 74576
rect 305328 74536 305334 74548
rect 305454 74536 305460 74548
rect 305512 74536 305518 74588
rect 307941 74579 307999 74585
rect 307941 74545 307953 74579
rect 307987 74576 307999 74579
rect 308122 74576 308128 74588
rect 307987 74548 308128 74576
rect 307987 74545 307999 74548
rect 307941 74539 307999 74545
rect 308122 74536 308128 74548
rect 308180 74536 308186 74588
rect 313645 74579 313703 74585
rect 313645 74545 313657 74579
rect 313691 74576 313703 74579
rect 313734 74576 313740 74588
rect 313691 74548 313740 74576
rect 313691 74545 313703 74548
rect 313645 74539 313703 74545
rect 313734 74536 313740 74548
rect 313792 74536 313798 74588
rect 229281 74511 229339 74517
rect 229281 74477 229293 74511
rect 229327 74508 229339 74511
rect 229370 74508 229376 74520
rect 229327 74480 229376 74508
rect 229327 74477 229339 74480
rect 229281 74471 229339 74477
rect 229370 74468 229376 74480
rect 229428 74468 229434 74520
rect 347961 74511 348019 74517
rect 347961 74477 347973 74511
rect 348007 74508 348019 74511
rect 348050 74508 348056 74520
rect 348007 74480 348056 74508
rect 348007 74477 348019 74480
rect 347961 74471 348019 74477
rect 348050 74468 348056 74480
rect 348108 74468 348114 74520
rect 305270 74440 305276 74452
rect 305231 74412 305276 74440
rect 305270 74400 305276 74412
rect 305328 74400 305334 74452
rect 288618 73788 288624 73840
rect 288676 73828 288682 73840
rect 288713 73831 288771 73837
rect 288713 73828 288725 73831
rect 288676 73800 288725 73828
rect 288676 73788 288682 73800
rect 288713 73797 288725 73800
rect 288759 73797 288771 73831
rect 288713 73791 288771 73797
rect 280522 73176 280528 73228
rect 280580 73216 280586 73228
rect 280614 73216 280620 73228
rect 280580 73188 280620 73216
rect 280580 73176 280586 73188
rect 280614 73176 280620 73188
rect 280672 73176 280678 73228
rect 289998 70864 290004 70916
rect 290056 70904 290062 70916
rect 290182 70904 290188 70916
rect 290056 70876 290188 70904
rect 290056 70864 290062 70876
rect 290182 70864 290188 70876
rect 290240 70864 290246 70916
rect 276290 70496 276296 70508
rect 276124 70468 276296 70496
rect 276124 70440 276152 70468
rect 276290 70456 276296 70468
rect 276348 70456 276354 70508
rect 287330 70456 287336 70508
rect 287388 70456 287394 70508
rect 328546 70456 328552 70508
rect 328604 70456 328610 70508
rect 346578 70456 346584 70508
rect 346636 70456 346642 70508
rect 276106 70388 276112 70440
rect 276164 70388 276170 70440
rect 287348 70372 287376 70456
rect 328564 70372 328592 70456
rect 346596 70372 346624 70456
rect 287330 70320 287336 70372
rect 287388 70320 287394 70372
rect 328546 70320 328552 70372
rect 328604 70320 328610 70372
rect 346578 70320 346584 70372
rect 346636 70320 346642 70372
rect 362957 70295 363015 70301
rect 362957 70261 362969 70295
rect 363003 70292 363015 70295
rect 363046 70292 363052 70304
rect 363003 70264 363052 70292
rect 363003 70261 363015 70264
rect 362957 70255 363015 70261
rect 363046 70252 363052 70264
rect 363104 70252 363110 70304
rect 324590 67736 324596 67788
rect 324648 67736 324654 67788
rect 435174 67736 435180 67788
rect 435232 67736 435238 67788
rect 324608 67652 324636 67736
rect 325970 67708 325976 67720
rect 325896 67680 325976 67708
rect 325896 67652 325924 67680
rect 325970 67668 325976 67680
rect 326028 67668 326034 67720
rect 435192 67652 435220 67736
rect 267090 67640 267096 67652
rect 267051 67612 267096 67640
rect 267090 67600 267096 67612
rect 267148 67600 267154 67652
rect 324590 67600 324596 67652
rect 324648 67600 324654 67652
rect 325878 67600 325884 67652
rect 325936 67600 325942 67652
rect 327350 67640 327356 67652
rect 327311 67612 327356 67640
rect 327350 67600 327356 67612
rect 327408 67600 327414 67652
rect 435174 67600 435180 67652
rect 435232 67600 435238 67652
rect 444098 67600 444104 67652
rect 444156 67640 444162 67652
rect 444190 67640 444196 67652
rect 444156 67612 444196 67640
rect 444156 67600 444162 67612
rect 444190 67600 444196 67612
rect 444248 67600 444254 67652
rect 244274 67572 244280 67584
rect 244235 67544 244280 67572
rect 244274 67532 244280 67544
rect 244332 67532 244338 67584
rect 252738 67532 252744 67584
rect 252796 67572 252802 67584
rect 252830 67572 252836 67584
rect 252796 67544 252836 67572
rect 252796 67532 252802 67544
rect 252830 67532 252836 67544
rect 252888 67532 252894 67584
rect 240410 66308 240416 66360
rect 240468 66348 240474 66360
rect 240505 66351 240563 66357
rect 240505 66348 240517 66351
rect 240468 66320 240517 66348
rect 240468 66308 240474 66320
rect 240505 66317 240517 66320
rect 240551 66317 240563 66351
rect 434254 66348 434260 66360
rect 434215 66320 434260 66348
rect 240505 66311 240563 66317
rect 434254 66308 434260 66320
rect 434312 66308 434318 66360
rect 248782 66280 248788 66292
rect 248743 66252 248788 66280
rect 248782 66240 248788 66252
rect 248840 66240 248846 66292
rect 262766 66280 262772 66292
rect 262727 66252 262772 66280
rect 262766 66240 262772 66252
rect 262824 66240 262830 66292
rect 291473 66283 291531 66289
rect 291473 66249 291485 66283
rect 291519 66280 291531 66283
rect 308030 66280 308036 66292
rect 291519 66252 291608 66280
rect 307991 66252 308036 66280
rect 291519 66249 291531 66252
rect 291473 66243 291531 66249
rect 255590 66212 255596 66224
rect 255551 66184 255596 66212
rect 255590 66172 255596 66184
rect 255648 66172 255654 66224
rect 291470 66104 291476 66156
rect 291528 66144 291534 66156
rect 291580 66144 291608 66252
rect 308030 66240 308036 66252
rect 308088 66240 308094 66292
rect 327350 66280 327356 66292
rect 327311 66252 327356 66280
rect 327350 66240 327356 66252
rect 327408 66240 327414 66292
rect 343729 66283 343787 66289
rect 343729 66249 343741 66283
rect 343775 66280 343787 66283
rect 343910 66280 343916 66292
rect 343775 66252 343916 66280
rect 343775 66249 343787 66252
rect 343729 66243 343787 66249
rect 343910 66240 343916 66252
rect 343968 66240 343974 66292
rect 309318 66172 309324 66224
rect 309376 66212 309382 66224
rect 309410 66212 309416 66224
rect 309376 66184 309416 66212
rect 309376 66172 309382 66184
rect 309410 66172 309416 66184
rect 309468 66172 309474 66224
rect 324590 66212 324596 66224
rect 324551 66184 324596 66212
rect 324590 66172 324596 66184
rect 324648 66172 324654 66224
rect 345198 66212 345204 66224
rect 345159 66184 345204 66212
rect 345198 66172 345204 66184
rect 345256 66172 345262 66224
rect 434254 66172 434260 66224
rect 434312 66172 434318 66224
rect 435174 66212 435180 66224
rect 435135 66184 435180 66212
rect 435174 66172 435180 66184
rect 435232 66172 435238 66224
rect 291528 66116 291608 66144
rect 434272 66144 434300 66172
rect 434438 66144 434444 66156
rect 434272 66116 434444 66144
rect 291528 66104 291534 66116
rect 434438 66104 434444 66116
rect 434496 66104 434502 66156
rect 229278 64988 229284 65000
rect 229239 64960 229284 64988
rect 229278 64948 229284 64960
rect 229336 64948 229342 65000
rect 233418 64880 233424 64932
rect 233476 64920 233482 64932
rect 233510 64920 233516 64932
rect 233476 64892 233516 64920
rect 233476 64880 233482 64892
rect 233510 64880 233516 64892
rect 233568 64880 233574 64932
rect 305273 64923 305331 64929
rect 305273 64889 305285 64923
rect 305319 64920 305331 64923
rect 305362 64920 305368 64932
rect 305319 64892 305368 64920
rect 305319 64889 305331 64892
rect 305273 64883 305331 64889
rect 305362 64880 305368 64892
rect 305420 64880 305426 64932
rect 308030 64920 308036 64932
rect 307991 64892 308036 64920
rect 308030 64880 308036 64892
rect 308088 64880 308094 64932
rect 310882 64880 310888 64932
rect 310940 64920 310946 64932
rect 310974 64920 310980 64932
rect 310940 64892 310980 64920
rect 310940 64880 310946 64892
rect 310974 64880 310980 64892
rect 311032 64880 311038 64932
rect 347958 64920 347964 64932
rect 347919 64892 347964 64920
rect 347958 64880 347964 64892
rect 348016 64880 348022 64932
rect 229278 64812 229284 64864
rect 229336 64852 229342 64864
rect 229462 64852 229468 64864
rect 229336 64824 229468 64852
rect 229336 64812 229342 64824
rect 229462 64812 229468 64824
rect 229520 64812 229526 64864
rect 234798 64852 234804 64864
rect 234759 64824 234804 64852
rect 234798 64812 234804 64824
rect 234856 64812 234862 64864
rect 240321 64855 240379 64861
rect 240321 64821 240333 64855
rect 240367 64852 240379 64855
rect 240410 64852 240416 64864
rect 240367 64824 240416 64852
rect 240367 64821 240379 64824
rect 240321 64815 240379 64821
rect 240410 64812 240416 64824
rect 240468 64812 240474 64864
rect 292758 64812 292764 64864
rect 292816 64852 292822 64864
rect 292850 64852 292856 64864
rect 292816 64824 292856 64852
rect 292816 64812 292822 64824
rect 292850 64812 292856 64824
rect 292908 64812 292914 64864
rect 255593 64719 255651 64725
rect 255593 64685 255605 64719
rect 255639 64716 255651 64719
rect 255774 64716 255780 64728
rect 255639 64688 255780 64716
rect 255639 64685 255651 64688
rect 255593 64679 255651 64685
rect 255774 64676 255780 64688
rect 255832 64676 255838 64728
rect 326798 63724 326804 63776
rect 326856 63764 326862 63776
rect 335262 63764 335268 63776
rect 326856 63736 335268 63764
rect 326856 63724 326862 63736
rect 335262 63724 335268 63736
rect 335320 63724 335326 63776
rect 398466 63724 398472 63776
rect 398524 63764 398530 63776
rect 399018 63764 399024 63776
rect 398524 63736 399024 63764
rect 398524 63724 398530 63736
rect 399018 63724 399024 63736
rect 399076 63724 399082 63776
rect 359550 63656 359556 63708
rect 359608 63696 359614 63708
rect 365622 63696 365628 63708
rect 359608 63668 365628 63696
rect 359608 63656 359614 63668
rect 365622 63656 365628 63668
rect 365680 63656 365686 63708
rect 417878 63656 417884 63708
rect 417936 63696 417942 63708
rect 419626 63696 419632 63708
rect 417936 63668 419632 63696
rect 417936 63656 417942 63668
rect 419626 63656 419632 63668
rect 419684 63656 419690 63708
rect 280246 63452 280252 63504
rect 280304 63492 280310 63504
rect 280522 63492 280528 63504
rect 280304 63464 280528 63492
rect 280304 63452 280310 63464
rect 280522 63452 280528 63464
rect 280580 63452 280586 63504
rect 267001 61115 267059 61121
rect 267001 61081 267013 61115
rect 267047 61112 267059 61115
rect 267090 61112 267096 61124
rect 267047 61084 267096 61112
rect 267047 61081 267059 61084
rect 267001 61075 267059 61081
rect 267090 61072 267096 61084
rect 267148 61072 267154 61124
rect 261294 60840 261300 60852
rect 261220 60812 261300 60840
rect 261220 60716 261248 60812
rect 261294 60800 261300 60812
rect 261352 60800 261358 60852
rect 444098 60840 444104 60852
rect 444024 60812 444104 60840
rect 444024 60716 444052 60812
rect 444098 60800 444104 60812
rect 444156 60800 444162 60852
rect 261202 60664 261208 60716
rect 261260 60664 261266 60716
rect 273346 60664 273352 60716
rect 273404 60664 273410 60716
rect 336918 60664 336924 60716
rect 336976 60704 336982 60716
rect 337102 60704 337108 60716
rect 336976 60676 337108 60704
rect 336976 60664 336982 60676
rect 337102 60664 337108 60676
rect 337160 60664 337166 60716
rect 363046 60664 363052 60716
rect 363104 60704 363110 60716
rect 363230 60704 363236 60716
rect 363104 60676 363236 60704
rect 363104 60664 363110 60676
rect 363230 60664 363236 60676
rect 363288 60664 363294 60716
rect 444006 60664 444012 60716
rect 444064 60664 444070 60716
rect 273364 60636 273392 60664
rect 273530 60636 273536 60648
rect 273364 60608 273536 60636
rect 273530 60596 273536 60608
rect 273588 60596 273594 60648
rect 310790 58760 310796 58812
rect 310848 58800 310854 58812
rect 310974 58800 310980 58812
rect 310848 58772 310980 58800
rect 310848 58760 310854 58772
rect 310974 58760 310980 58772
rect 311032 58760 311038 58812
rect 325878 58012 325884 58064
rect 325936 58012 325942 58064
rect 244274 57984 244280 57996
rect 244235 57956 244280 57984
rect 244274 57944 244280 57956
rect 244332 57944 244338 57996
rect 287330 57944 287336 57996
rect 287388 57984 287394 57996
rect 287422 57984 287428 57996
rect 287388 57956 287428 57984
rect 287388 57944 287394 57956
rect 287422 57944 287428 57956
rect 287480 57944 287486 57996
rect 288710 57984 288716 57996
rect 288671 57956 288716 57984
rect 288710 57944 288716 57956
rect 288768 57944 288774 57996
rect 325896 57928 325924 58012
rect 239033 57919 239091 57925
rect 239033 57885 239045 57919
rect 239079 57916 239091 57919
rect 239122 57916 239128 57928
rect 239079 57888 239128 57916
rect 239079 57885 239091 57888
rect 239033 57879 239091 57885
rect 239122 57876 239128 57888
rect 239180 57876 239186 57928
rect 245930 57916 245936 57928
rect 245891 57888 245936 57916
rect 245930 57876 245936 57888
rect 245988 57876 245994 57928
rect 325878 57876 325884 57928
rect 325936 57876 325942 57928
rect 336921 57919 336979 57925
rect 336921 57885 336933 57919
rect 336967 57916 336979 57919
rect 337102 57916 337108 57928
rect 336967 57888 337108 57916
rect 336967 57885 336979 57888
rect 336921 57879 336979 57885
rect 337102 57876 337108 57888
rect 337160 57876 337166 57928
rect 363141 57919 363199 57925
rect 363141 57885 363153 57919
rect 363187 57916 363199 57919
rect 363230 57916 363236 57928
rect 363187 57888 363236 57916
rect 363187 57885 363199 57888
rect 363141 57879 363199 57885
rect 363230 57876 363236 57888
rect 363288 57876 363294 57928
rect 313734 56652 313740 56704
rect 313792 56652 313798 56704
rect 249978 56584 249984 56636
rect 250036 56624 250042 56636
rect 250070 56624 250076 56636
rect 250036 56596 250076 56624
rect 250036 56584 250042 56596
rect 250070 56584 250076 56596
rect 250128 56584 250134 56636
rect 262674 56584 262680 56636
rect 262732 56624 262738 56636
rect 262858 56624 262864 56636
rect 262732 56596 262864 56624
rect 262732 56584 262738 56596
rect 262858 56584 262864 56596
rect 262916 56584 262922 56636
rect 266998 56624 267004 56636
rect 266959 56596 267004 56624
rect 266998 56584 267004 56596
rect 267056 56584 267062 56636
rect 309410 56584 309416 56636
rect 309468 56584 309474 56636
rect 254118 56556 254124 56568
rect 254079 56528 254124 56556
rect 254118 56516 254124 56528
rect 254176 56516 254182 56568
rect 262674 56448 262680 56500
rect 262732 56488 262738 56500
rect 262858 56488 262864 56500
rect 262732 56460 262864 56488
rect 262732 56448 262738 56460
rect 262858 56448 262864 56460
rect 262916 56448 262922 56500
rect 309428 56488 309456 56584
rect 313752 56568 313780 56652
rect 345198 56624 345204 56636
rect 345159 56596 345204 56624
rect 345198 56584 345204 56596
rect 345256 56584 345262 56636
rect 313734 56516 313740 56568
rect 313792 56516 313798 56568
rect 309502 56488 309508 56500
rect 309428 56460 309508 56488
rect 309502 56448 309508 56460
rect 309560 56448 309566 56500
rect 290090 55332 290096 55344
rect 290016 55304 290096 55332
rect 290016 55276 290044 55304
rect 290090 55292 290096 55304
rect 290148 55292 290154 55344
rect 234798 55264 234804 55276
rect 234759 55236 234804 55264
rect 234798 55224 234804 55236
rect 234856 55224 234862 55276
rect 240318 55264 240324 55276
rect 240279 55236 240324 55264
rect 240318 55224 240324 55236
rect 240376 55224 240382 55276
rect 289998 55224 290004 55276
rect 290056 55224 290062 55276
rect 255593 55199 255651 55205
rect 255593 55165 255605 55199
rect 255639 55196 255651 55199
rect 255774 55196 255780 55208
rect 255639 55168 255780 55196
rect 255639 55165 255651 55168
rect 255593 55159 255651 55165
rect 255774 55156 255780 55168
rect 255832 55156 255838 55208
rect 347869 55199 347927 55205
rect 347869 55165 347881 55199
rect 347915 55196 347927 55199
rect 347958 55196 347964 55208
rect 347915 55168 347964 55196
rect 347915 55165 347927 55168
rect 347869 55159 347927 55165
rect 347958 55156 347964 55168
rect 348016 55156 348022 55208
rect 289998 55128 290004 55140
rect 289959 55100 290004 55128
rect 289998 55088 290004 55100
rect 290056 55088 290062 55140
rect 252738 53116 252744 53168
rect 252796 53116 252802 53168
rect 261202 53156 261208 53168
rect 261163 53128 261208 53156
rect 261202 53116 261208 53128
rect 261260 53116 261266 53168
rect 327350 53156 327356 53168
rect 327276 53128 327356 53156
rect 252756 53088 252784 53116
rect 327276 53100 327304 53128
rect 327350 53116 327356 53128
rect 327408 53116 327414 53168
rect 252830 53088 252836 53100
rect 252756 53060 252836 53088
rect 252830 53048 252836 53060
rect 252888 53048 252894 53100
rect 324593 53091 324651 53097
rect 324593 53057 324605 53091
rect 324639 53088 324651 53091
rect 324774 53088 324780 53100
rect 324639 53060 324780 53088
rect 324639 53057 324651 53060
rect 324593 53051 324651 53057
rect 324774 53048 324780 53060
rect 324832 53048 324838 53100
rect 327258 53048 327264 53100
rect 327316 53048 327322 53100
rect 287330 51252 287336 51264
rect 287256 51224 287336 51252
rect 229370 51116 229376 51128
rect 229296 51088 229376 51116
rect 229296 51060 229324 51088
rect 229370 51076 229376 51088
rect 229428 51076 229434 51128
rect 287256 51060 287284 51224
rect 287330 51212 287336 51224
rect 287388 51212 287394 51264
rect 299842 51184 299848 51196
rect 299803 51156 299848 51184
rect 299842 51144 299848 51156
rect 299900 51144 299906 51196
rect 342530 51184 342536 51196
rect 342491 51156 342536 51184
rect 342530 51144 342536 51156
rect 342588 51144 342594 51196
rect 346578 51184 346584 51196
rect 346539 51156 346584 51184
rect 346578 51144 346584 51156
rect 346636 51144 346642 51196
rect 434346 51116 434352 51128
rect 434272 51088 434352 51116
rect 434272 51060 434300 51088
rect 434346 51076 434352 51088
rect 434404 51076 434410 51128
rect 229278 51008 229284 51060
rect 229336 51008 229342 51060
rect 239030 51048 239036 51060
rect 238991 51020 239036 51048
rect 239030 51008 239036 51020
rect 239088 51008 239094 51060
rect 287238 51008 287244 51060
rect 287296 51008 287302 51060
rect 434254 51008 434260 51060
rect 434312 51008 434318 51060
rect 435174 51048 435180 51060
rect 435135 51020 435180 51048
rect 435174 51008 435180 51020
rect 435232 51008 435238 51060
rect 444006 51008 444012 51060
rect 444064 51048 444070 51060
rect 444190 51048 444196 51060
rect 444064 51020 444196 51048
rect 444064 51008 444070 51020
rect 444190 51008 444196 51020
rect 444248 51008 444254 51060
rect 240318 48288 240324 48340
rect 240376 48328 240382 48340
rect 240410 48328 240416 48340
rect 240376 48300 240416 48328
rect 240376 48288 240382 48300
rect 240410 48288 240416 48300
rect 240468 48288 240474 48340
rect 245930 48328 245936 48340
rect 245891 48300 245936 48328
rect 245930 48288 245936 48300
rect 245988 48288 245994 48340
rect 261205 48331 261263 48337
rect 261205 48297 261217 48331
rect 261251 48328 261263 48331
rect 261294 48328 261300 48340
rect 261251 48300 261300 48328
rect 261251 48297 261263 48300
rect 261205 48291 261263 48297
rect 261294 48288 261300 48300
rect 261352 48288 261358 48340
rect 299842 48328 299848 48340
rect 299803 48300 299848 48328
rect 299842 48288 299848 48300
rect 299900 48288 299906 48340
rect 336918 48328 336924 48340
rect 336879 48300 336924 48328
rect 336918 48288 336924 48300
rect 336976 48288 336982 48340
rect 363138 48328 363144 48340
rect 363099 48300 363144 48328
rect 363138 48288 363144 48300
rect 363196 48288 363202 48340
rect 239030 48220 239036 48272
rect 239088 48260 239094 48272
rect 239122 48260 239128 48272
rect 239088 48232 239128 48260
rect 239088 48220 239094 48232
rect 239122 48220 239128 48232
rect 239180 48220 239186 48272
rect 267093 48263 267151 48269
rect 267093 48229 267105 48263
rect 267139 48260 267151 48263
rect 267182 48260 267188 48272
rect 267139 48232 267188 48260
rect 267139 48229 267151 48232
rect 267093 48223 267151 48229
rect 267182 48220 267188 48232
rect 267240 48220 267246 48272
rect 288618 48220 288624 48272
rect 288676 48260 288682 48272
rect 288802 48260 288808 48272
rect 288676 48232 288808 48260
rect 288676 48220 288682 48232
rect 288802 48220 288808 48232
rect 288860 48220 288866 48272
rect 435266 48260 435272 48272
rect 435227 48232 435272 48260
rect 435266 48220 435272 48232
rect 435324 48220 435330 48272
rect 444101 48263 444159 48269
rect 444101 48229 444113 48263
rect 444147 48260 444159 48263
rect 444190 48260 444196 48272
rect 444147 48232 444196 48260
rect 444147 48229 444159 48232
rect 444101 48223 444159 48229
rect 444190 48220 444196 48232
rect 444248 48220 444254 48272
rect 254118 46968 254124 46980
rect 254079 46940 254124 46968
rect 254118 46928 254124 46940
rect 254176 46928 254182 46980
rect 291470 46928 291476 46980
rect 291528 46968 291534 46980
rect 291562 46968 291568 46980
rect 291528 46940 291568 46968
rect 291528 46928 291534 46940
rect 291562 46928 291568 46940
rect 291620 46928 291626 46980
rect 342530 46968 342536 46980
rect 342491 46940 342536 46968
rect 342530 46928 342536 46940
rect 342588 46928 342594 46980
rect 251358 46860 251364 46912
rect 251416 46900 251422 46912
rect 251450 46900 251456 46912
rect 251416 46872 251456 46900
rect 251416 46860 251422 46872
rect 251450 46860 251456 46872
rect 251508 46860 251514 46912
rect 262858 46860 262864 46912
rect 262916 46900 262922 46912
rect 345198 46900 345204 46912
rect 262916 46872 262961 46900
rect 345159 46872 345204 46900
rect 262916 46860 262922 46872
rect 345198 46860 345204 46872
rect 345256 46860 345262 46912
rect 325878 46792 325884 46844
rect 325936 46832 325942 46844
rect 326154 46832 326160 46844
rect 325936 46804 326160 46832
rect 325936 46792 325942 46804
rect 326154 46792 326160 46804
rect 326212 46792 326218 46844
rect 255590 45676 255596 45688
rect 255551 45648 255596 45676
rect 255590 45636 255596 45648
rect 255648 45636 255654 45688
rect 347869 45679 347927 45685
rect 347869 45645 347881 45679
rect 347915 45676 347927 45679
rect 347958 45676 347964 45688
rect 347915 45648 347964 45676
rect 347915 45645 347927 45648
rect 347869 45639 347927 45645
rect 347958 45636 347964 45648
rect 348016 45636 348022 45688
rect 289998 45608 290004 45620
rect 289959 45580 290004 45608
rect 289998 45568 290004 45580
rect 290056 45568 290062 45620
rect 346578 45608 346584 45620
rect 346539 45580 346584 45608
rect 346578 45568 346584 45580
rect 346636 45568 346642 45620
rect 234798 45540 234804 45552
rect 234759 45512 234804 45540
rect 234798 45500 234804 45512
rect 234856 45500 234862 45552
rect 234982 45500 234988 45552
rect 235040 45540 235046 45552
rect 235166 45540 235172 45552
rect 235040 45512 235172 45540
rect 235040 45500 235046 45512
rect 235166 45500 235172 45512
rect 235224 45500 235230 45552
rect 255590 45500 255596 45552
rect 255648 45540 255654 45552
rect 255682 45540 255688 45552
rect 255648 45512 255688 45540
rect 255648 45500 255654 45512
rect 255682 45500 255688 45512
rect 255740 45500 255746 45552
rect 299842 45500 299848 45552
rect 299900 45540 299906 45552
rect 299934 45540 299940 45552
rect 299900 45512 299940 45540
rect 299900 45500 299906 45512
rect 299934 45500 299940 45512
rect 299992 45500 299998 45552
rect 280246 44480 280252 44532
rect 280304 44520 280310 44532
rect 280525 44523 280583 44529
rect 280525 44520 280537 44523
rect 280304 44492 280537 44520
rect 280304 44480 280310 44492
rect 280525 44489 280537 44492
rect 280571 44489 280583 44523
rect 280525 44483 280583 44489
rect 241790 44112 241796 44124
rect 241751 44084 241796 44112
rect 241790 44072 241796 44084
rect 241848 44072 241854 44124
rect 229278 41460 229284 41472
rect 229239 41432 229284 41460
rect 229278 41420 229284 41432
rect 229336 41420 229342 41472
rect 313550 41420 313556 41472
rect 313608 41460 313614 41472
rect 313734 41460 313740 41472
rect 313608 41432 313740 41460
rect 313608 41420 313614 41432
rect 313734 41420 313740 41432
rect 313792 41420 313798 41472
rect 363046 41352 363052 41404
rect 363104 41392 363110 41404
rect 363230 41392 363236 41404
rect 363104 41364 363236 41392
rect 363104 41352 363110 41364
rect 363230 41352 363236 41364
rect 363288 41352 363294 41404
rect 270494 40332 270500 40384
rect 270552 40372 270558 40384
rect 280522 40372 280528 40384
rect 270552 40344 280528 40372
rect 270552 40332 270558 40344
rect 280522 40332 280528 40344
rect 280580 40332 280586 40384
rect 398466 40196 398472 40248
rect 398524 40236 398530 40248
rect 399018 40236 399024 40248
rect 398524 40208 399024 40236
rect 398524 40196 398530 40208
rect 399018 40196 399024 40208
rect 399076 40196 399082 40248
rect 417878 40196 417884 40248
rect 417936 40236 417942 40248
rect 418338 40236 418344 40248
rect 417936 40208 418344 40236
rect 417936 40196 417942 40208
rect 418338 40196 418344 40208
rect 418396 40196 418402 40248
rect 356054 40060 356060 40112
rect 356112 40100 356118 40112
rect 365622 40100 365628 40112
rect 356112 40072 365628 40100
rect 356112 40060 356118 40072
rect 365622 40060 365628 40072
rect 365680 40060 365686 40112
rect 229281 38743 229339 38749
rect 229281 38709 229293 38743
rect 229327 38740 229339 38743
rect 229370 38740 229376 38752
rect 229327 38712 229376 38740
rect 229327 38709 229339 38712
rect 229281 38703 229339 38709
rect 229370 38700 229376 38712
rect 229428 38700 229434 38752
rect 287238 38700 287244 38752
rect 287296 38700 287302 38752
rect 267090 38672 267096 38684
rect 267051 38644 267096 38672
rect 267090 38632 267096 38644
rect 267148 38632 267154 38684
rect 273254 38632 273260 38684
rect 273312 38672 273318 38684
rect 273530 38672 273536 38684
rect 273312 38644 273536 38672
rect 273312 38632 273318 38644
rect 273530 38632 273536 38644
rect 273588 38632 273594 38684
rect 287256 38616 287284 38700
rect 435269 38675 435327 38681
rect 435269 38641 435281 38675
rect 435315 38672 435327 38675
rect 435358 38672 435364 38684
rect 435315 38644 435364 38672
rect 435315 38641 435327 38644
rect 435269 38635 435327 38641
rect 435358 38632 435364 38644
rect 435416 38632 435422 38684
rect 444098 38672 444104 38684
rect 444059 38644 444104 38672
rect 444098 38632 444104 38644
rect 444156 38632 444162 38684
rect 245930 38604 245936 38616
rect 245891 38576 245936 38604
rect 245930 38564 245936 38576
rect 245988 38564 245994 38616
rect 287238 38564 287244 38616
rect 287296 38564 287302 38616
rect 324774 38564 324780 38616
rect 324832 38564 324838 38616
rect 363141 38607 363199 38613
rect 363141 38573 363153 38607
rect 363187 38604 363199 38607
rect 363230 38604 363236 38616
rect 363187 38576 363236 38604
rect 363187 38573 363199 38576
rect 363141 38567 363199 38573
rect 363230 38564 363236 38576
rect 363288 38564 363294 38616
rect 324792 38480 324820 38564
rect 324774 38428 324780 38480
rect 324832 38428 324838 38480
rect 254118 37272 254124 37324
rect 254176 37312 254182 37324
rect 254210 37312 254216 37324
rect 254176 37284 254216 37312
rect 254176 37272 254182 37284
rect 254210 37272 254216 37284
rect 254268 37272 254274 37324
rect 262674 37272 262680 37324
rect 262732 37312 262738 37324
rect 262861 37315 262919 37321
rect 262861 37312 262873 37315
rect 262732 37284 262873 37312
rect 262732 37272 262738 37284
rect 262861 37281 262873 37284
rect 262907 37281 262919 37315
rect 262861 37275 262919 37281
rect 267001 37247 267059 37253
rect 267001 37213 267013 37247
rect 267047 37244 267059 37247
rect 267090 37244 267096 37256
rect 267047 37216 267096 37244
rect 267047 37213 267059 37216
rect 267001 37207 267059 37213
rect 267090 37204 267096 37216
rect 267148 37204 267154 37256
rect 234798 35952 234804 35964
rect 234759 35924 234804 35952
rect 234798 35912 234804 35924
rect 234856 35912 234862 35964
rect 289998 35884 290004 35896
rect 289959 35856 290004 35884
rect 289998 35844 290004 35856
rect 290056 35844 290062 35896
rect 299750 35844 299756 35896
rect 299808 35884 299814 35896
rect 300026 35884 300032 35896
rect 299808 35856 300032 35884
rect 299808 35844 299814 35856
rect 300026 35844 300032 35856
rect 300084 35844 300090 35896
rect 305362 35884 305368 35896
rect 305323 35856 305368 35884
rect 305362 35844 305368 35856
rect 305420 35844 305426 35896
rect 434438 35068 434444 35080
rect 434399 35040 434444 35068
rect 434438 35028 434444 35040
rect 434496 35028 434502 35080
rect 307938 34484 307944 34536
rect 307996 34524 308002 34536
rect 308122 34524 308128 34536
rect 307996 34496 308128 34524
rect 307996 34484 308002 34496
rect 308122 34484 308128 34496
rect 308180 34484 308186 34536
rect 253934 32376 253940 32428
rect 253992 32416 253998 32428
rect 254210 32416 254216 32428
rect 253992 32388 254216 32416
rect 253992 32376 253998 32388
rect 254210 32376 254216 32388
rect 254268 32376 254274 32428
rect 328546 31872 328552 31884
rect 328507 31844 328552 31872
rect 328546 31832 328552 31844
rect 328604 31832 328610 31884
rect 444098 31872 444104 31884
rect 444059 31844 444104 31872
rect 444098 31832 444104 31844
rect 444156 31832 444162 31884
rect 229278 31764 229284 31816
rect 229336 31764 229342 31816
rect 261202 31804 261208 31816
rect 261163 31776 261208 31804
rect 261202 31764 261208 31776
rect 261260 31764 261266 31816
rect 229296 31668 229324 31764
rect 229370 31668 229376 31680
rect 229296 31640 229376 31668
rect 229370 31628 229376 31640
rect 229428 31628 229434 31680
rect 292761 30719 292819 30725
rect 292761 30685 292773 30719
rect 292807 30716 292819 30719
rect 292850 30716 292856 30728
rect 292807 30688 292856 30716
rect 292807 30685 292819 30688
rect 292761 30679 292819 30685
rect 292850 30676 292856 30688
rect 292908 30676 292914 30728
rect 270494 29180 270500 29232
rect 270552 29220 270558 29232
rect 273990 29220 273996 29232
rect 270552 29192 273996 29220
rect 270552 29180 270558 29192
rect 273990 29180 273996 29192
rect 274048 29180 274054 29232
rect 398466 29180 398472 29232
rect 398524 29220 398530 29232
rect 399018 29220 399024 29232
rect 398524 29192 399024 29220
rect 398524 29180 398530 29192
rect 399018 29180 399024 29192
rect 399076 29180 399082 29232
rect 476022 29180 476028 29232
rect 476080 29220 476086 29232
rect 482922 29220 482928 29232
rect 476080 29192 482928 29220
rect 476080 29180 476086 29192
rect 482922 29180 482928 29192
rect 482980 29180 482986 29232
rect 417878 29112 417884 29164
rect 417936 29152 417942 29164
rect 418154 29152 418160 29164
rect 417936 29124 418160 29152
rect 417936 29112 417942 29124
rect 418154 29112 418160 29124
rect 418212 29112 418218 29164
rect 342438 29044 342444 29096
rect 342496 29044 342502 29096
rect 434441 29087 434499 29093
rect 434441 29053 434453 29087
rect 434487 29084 434499 29087
rect 434530 29084 434536 29096
rect 434487 29056 434536 29084
rect 434487 29053 434499 29056
rect 434441 29047 434499 29053
rect 434530 29044 434536 29056
rect 434588 29044 434594 29096
rect 444374 29044 444380 29096
rect 444432 29084 444438 29096
rect 449250 29084 449256 29096
rect 444432 29056 449256 29084
rect 444432 29044 444438 29056
rect 449250 29044 449256 29056
rect 449308 29044 449314 29096
rect 241790 29016 241796 29028
rect 241751 28988 241796 29016
rect 241790 28976 241796 28988
rect 241848 28976 241854 29028
rect 245930 29016 245936 29028
rect 245891 28988 245936 29016
rect 245930 28976 245936 28988
rect 245988 28976 245994 29028
rect 342456 29016 342484 29044
rect 342530 29016 342536 29028
rect 342456 28988 342536 29016
rect 342530 28976 342536 28988
rect 342588 28976 342594 29028
rect 345201 29019 345259 29025
rect 345201 28985 345213 29019
rect 345247 29016 345259 29019
rect 345290 29016 345296 29028
rect 345247 28988 345296 29016
rect 345247 28985 345259 28988
rect 345201 28979 345259 28985
rect 345290 28976 345296 28988
rect 345348 28976 345354 29028
rect 363138 29016 363144 29028
rect 363099 28988 363144 29016
rect 363138 28976 363144 28988
rect 363196 28976 363202 29028
rect 444098 29016 444104 29028
rect 444059 28988 444104 29016
rect 444098 28976 444104 28988
rect 444156 28976 444162 29028
rect 298554 28908 298560 28960
rect 298612 28948 298618 28960
rect 298646 28948 298652 28960
rect 298612 28920 298652 28948
rect 298612 28908 298618 28920
rect 298646 28908 298652 28920
rect 298704 28908 298710 28960
rect 324590 28948 324596 28960
rect 324551 28920 324596 28948
rect 324590 28908 324596 28920
rect 324648 28908 324654 28960
rect 327258 28908 327264 28960
rect 327316 28948 327322 28960
rect 327442 28948 327448 28960
rect 327316 28920 327448 28948
rect 327316 28908 327322 28920
rect 327442 28908 327448 28920
rect 327500 28908 327506 28960
rect 435269 28951 435327 28957
rect 435269 28917 435281 28951
rect 435315 28948 435327 28951
rect 435358 28948 435364 28960
rect 435315 28920 435364 28948
rect 435315 28917 435327 28920
rect 435269 28911 435327 28917
rect 435358 28908 435364 28920
rect 435416 28908 435422 28960
rect 280522 28880 280528 28892
rect 280483 28852 280528 28880
rect 280522 28840 280528 28852
rect 280580 28840 280586 28892
rect 261202 27656 261208 27668
rect 261163 27628 261208 27656
rect 261202 27616 261208 27628
rect 261260 27616 261266 27668
rect 266998 27656 267004 27668
rect 266959 27628 267004 27656
rect 266998 27616 267004 27628
rect 267056 27616 267062 27668
rect 328546 27656 328552 27668
rect 328507 27628 328552 27656
rect 328546 27616 328552 27628
rect 328604 27616 328610 27668
rect 251361 27591 251419 27597
rect 251361 27557 251373 27591
rect 251407 27588 251419 27591
rect 251450 27588 251456 27600
rect 251407 27560 251456 27588
rect 251407 27557 251419 27560
rect 251361 27551 251419 27557
rect 251450 27548 251456 27560
rect 251508 27548 251514 27600
rect 342441 27591 342499 27597
rect 342441 27557 342453 27591
rect 342487 27588 342499 27591
rect 342530 27588 342536 27600
rect 342487 27560 342536 27588
rect 342487 27557 342499 27560
rect 342441 27551 342499 27557
rect 342530 27548 342536 27560
rect 342588 27548 342594 27600
rect 345201 27591 345259 27597
rect 345201 27557 345213 27591
rect 345247 27588 345259 27591
rect 345290 27588 345296 27600
rect 345247 27560 345296 27588
rect 345247 27557 345259 27560
rect 345201 27551 345259 27557
rect 345290 27548 345296 27560
rect 345348 27548 345354 27600
rect 434530 27548 434536 27600
rect 434588 27588 434594 27600
rect 434625 27591 434683 27597
rect 434625 27588 434637 27591
rect 434588 27560 434637 27588
rect 434588 27548 434594 27560
rect 434625 27557 434637 27560
rect 434671 27557 434683 27591
rect 434625 27551 434683 27557
rect 290001 26299 290059 26305
rect 290001 26265 290013 26299
rect 290047 26296 290059 26299
rect 290182 26296 290188 26308
rect 290047 26268 290188 26296
rect 290047 26265 290059 26268
rect 290001 26259 290059 26265
rect 290182 26256 290188 26268
rect 290240 26256 290246 26308
rect 292758 26296 292764 26308
rect 292719 26268 292764 26296
rect 292758 26256 292764 26268
rect 292816 26256 292822 26308
rect 234798 26228 234804 26240
rect 234759 26200 234804 26228
rect 234798 26188 234804 26200
rect 234856 26188 234862 26240
rect 234893 26231 234951 26237
rect 234893 26197 234905 26231
rect 234939 26228 234951 26231
rect 235074 26228 235080 26240
rect 234939 26200 235080 26228
rect 234939 26197 234951 26200
rect 234893 26191 234951 26197
rect 235074 26188 235080 26200
rect 235132 26188 235138 26240
rect 238941 26231 238999 26237
rect 238941 26197 238953 26231
rect 238987 26228 238999 26231
rect 239122 26228 239128 26240
rect 238987 26200 239128 26228
rect 238987 26197 238999 26200
rect 238941 26191 238999 26197
rect 239122 26188 239128 26200
rect 239180 26188 239186 26240
rect 346397 26231 346455 26237
rect 346397 26197 346409 26231
rect 346443 26228 346455 26231
rect 346578 26228 346584 26240
rect 346443 26200 346584 26228
rect 346443 26197 346455 26200
rect 346397 26191 346455 26197
rect 346578 26188 346584 26200
rect 346636 26188 346642 26240
rect 305362 24868 305368 24880
rect 305323 24840 305368 24868
rect 305362 24828 305368 24840
rect 305420 24828 305426 24880
rect 262585 24191 262643 24197
rect 262585 24157 262597 24191
rect 262631 24188 262643 24191
rect 262674 24188 262680 24200
rect 262631 24160 262680 24188
rect 262631 24157 262643 24160
rect 262585 24151 262643 24157
rect 262674 24148 262680 24160
rect 262732 24148 262738 24200
rect 252741 22763 252799 22769
rect 252741 22729 252753 22763
rect 252787 22760 252799 22763
rect 252830 22760 252836 22772
rect 252787 22732 252836 22760
rect 252787 22729 252799 22732
rect 252741 22723 252799 22729
rect 252830 22720 252836 22732
rect 252888 22720 252894 22772
rect 253934 22720 253940 22772
rect 253992 22760 253998 22772
rect 254121 22763 254179 22769
rect 254121 22760 254133 22763
rect 253992 22732 254133 22760
rect 253992 22720 253998 22732
rect 254121 22729 254133 22732
rect 254167 22729 254179 22763
rect 254121 22723 254179 22729
rect 255314 22720 255320 22772
rect 255372 22760 255378 22772
rect 255682 22760 255688 22772
rect 255372 22732 255688 22760
rect 255372 22720 255378 22732
rect 255682 22720 255688 22732
rect 255740 22720 255746 22772
rect 328457 22763 328515 22769
rect 328457 22729 328469 22763
rect 328503 22760 328515 22763
rect 328546 22760 328552 22772
rect 328503 22732 328552 22760
rect 328503 22729 328515 22732
rect 328457 22723 328515 22729
rect 328546 22720 328552 22732
rect 328604 22720 328610 22772
rect 245930 22148 245936 22160
rect 245764 22120 245936 22148
rect 245764 22092 245792 22120
rect 245930 22108 245936 22120
rect 245988 22108 245994 22160
rect 245746 22040 245752 22092
rect 245804 22040 245810 22092
rect 363046 22040 363052 22092
rect 363104 22080 363110 22092
rect 363230 22080 363236 22092
rect 363104 22052 363236 22080
rect 363104 22040 363110 22052
rect 363230 22040 363236 22052
rect 363288 22040 363294 22092
rect 308122 19496 308128 19508
rect 308083 19468 308128 19496
rect 308122 19456 308128 19468
rect 308180 19456 308186 19508
rect 244550 19428 244556 19440
rect 244476 19400 244556 19428
rect 244476 19372 244504 19400
rect 244550 19388 244556 19400
rect 244608 19388 244614 19440
rect 248782 19428 248788 19440
rect 248708 19400 248788 19428
rect 248708 19372 248736 19400
rect 248782 19388 248788 19400
rect 248840 19388 248846 19440
rect 244458 19320 244464 19372
rect 244516 19320 244522 19372
rect 248690 19320 248696 19372
rect 248748 19320 248754 19372
rect 249978 19320 249984 19372
rect 250036 19360 250042 19372
rect 250070 19360 250076 19372
rect 250036 19332 250076 19360
rect 250036 19320 250042 19332
rect 250070 19320 250076 19332
rect 250128 19320 250134 19372
rect 261110 19320 261116 19372
rect 261168 19360 261174 19372
rect 261202 19360 261208 19372
rect 261168 19332 261208 19360
rect 261168 19320 261174 19332
rect 261202 19320 261208 19332
rect 261260 19320 261266 19372
rect 262582 19360 262588 19372
rect 262543 19332 262588 19360
rect 262582 19320 262588 19332
rect 262640 19320 262646 19372
rect 288710 19320 288716 19372
rect 288768 19360 288774 19372
rect 288986 19360 288992 19372
rect 288768 19332 288992 19360
rect 288768 19320 288774 19332
rect 288986 19320 288992 19332
rect 289044 19320 289050 19372
rect 292758 19320 292764 19372
rect 292816 19360 292822 19372
rect 292850 19360 292856 19372
rect 292816 19332 292856 19360
rect 292816 19320 292822 19332
rect 292850 19320 292856 19332
rect 292908 19320 292914 19372
rect 324590 19360 324596 19372
rect 324551 19332 324596 19360
rect 324590 19320 324596 19332
rect 324648 19320 324654 19372
rect 435266 19360 435272 19372
rect 435227 19332 435272 19360
rect 435266 19320 435272 19332
rect 435324 19320 435330 19372
rect 327261 19295 327319 19301
rect 327261 19261 327273 19295
rect 327307 19292 327319 19295
rect 327350 19292 327356 19304
rect 327307 19264 327356 19292
rect 327307 19261 327319 19264
rect 327261 19255 327319 19261
rect 327350 19252 327356 19264
rect 327408 19252 327414 19304
rect 363230 19292 363236 19304
rect 363191 19264 363236 19292
rect 363230 19252 363236 19264
rect 363288 19252 363294 19304
rect 310790 18068 310796 18080
rect 310716 18040 310796 18068
rect 310716 18012 310744 18040
rect 310790 18028 310796 18040
rect 310848 18028 310854 18080
rect 251361 18003 251419 18009
rect 251361 17969 251373 18003
rect 251407 17969 251419 18003
rect 251361 17963 251419 17969
rect 229189 17935 229247 17941
rect 229189 17901 229201 17935
rect 229235 17932 229247 17935
rect 229370 17932 229376 17944
rect 229235 17904 229376 17932
rect 229235 17901 229247 17904
rect 229189 17895 229247 17901
rect 229370 17892 229376 17904
rect 229428 17892 229434 17944
rect 240229 17935 240287 17941
rect 240229 17901 240241 17935
rect 240275 17932 240287 17935
rect 240318 17932 240324 17944
rect 240275 17904 240324 17932
rect 240275 17901 240287 17904
rect 240229 17895 240287 17901
rect 240318 17892 240324 17904
rect 240376 17892 240382 17944
rect 241606 17932 241612 17944
rect 241567 17904 241612 17932
rect 241606 17892 241612 17904
rect 241664 17892 241670 17944
rect 251376 17932 251404 17963
rect 280430 17960 280436 18012
rect 280488 18000 280494 18012
rect 280522 18000 280528 18012
rect 280488 17972 280528 18000
rect 280488 17960 280494 17972
rect 280522 17960 280528 17972
rect 280580 17960 280586 18012
rect 310698 17960 310704 18012
rect 310756 17960 310762 18012
rect 434530 17960 434536 18012
rect 434588 18000 434594 18012
rect 434625 18003 434683 18009
rect 434625 18000 434637 18003
rect 434588 17972 434637 18000
rect 434588 17960 434594 17972
rect 434625 17969 434637 17972
rect 434671 17969 434683 18003
rect 434625 17963 434683 17969
rect 251542 17932 251548 17944
rect 251376 17904 251548 17932
rect 251542 17892 251548 17904
rect 251600 17892 251606 17944
rect 434530 17008 434536 17060
rect 434588 17008 434594 17060
rect 434622 17008 434628 17060
rect 434680 17008 434686 17060
rect 434548 16856 434576 17008
rect 434640 16856 434668 17008
rect 398466 16804 398472 16856
rect 398524 16844 398530 16856
rect 399018 16844 399024 16856
rect 398524 16816 399024 16844
rect 398524 16804 398530 16816
rect 399018 16804 399024 16816
rect 399076 16804 399082 16856
rect 434530 16804 434536 16856
rect 434588 16804 434594 16856
rect 434622 16804 434628 16856
rect 434680 16804 434686 16856
rect 476022 16804 476028 16856
rect 476080 16844 476086 16856
rect 482922 16844 482928 16856
rect 476080 16816 482928 16844
rect 476080 16804 476086 16816
rect 482922 16804 482928 16816
rect 482980 16804 482986 16856
rect 360010 16736 360016 16788
rect 360068 16776 360074 16788
rect 361114 16776 361120 16788
rect 360068 16748 361120 16776
rect 360068 16736 360074 16748
rect 361114 16736 361120 16748
rect 361172 16736 361178 16788
rect 299845 16711 299903 16717
rect 299845 16677 299857 16711
rect 299891 16708 299903 16711
rect 300026 16708 300032 16720
rect 299891 16680 300032 16708
rect 299891 16677 299903 16680
rect 299845 16671 299903 16677
rect 300026 16668 300032 16680
rect 300084 16668 300090 16720
rect 425054 16668 425060 16720
rect 425112 16708 425118 16720
rect 434438 16708 434444 16720
rect 425112 16680 434444 16708
rect 425112 16668 425118 16680
rect 434438 16668 434444 16680
rect 434496 16668 434502 16720
rect 444374 16668 444380 16720
rect 444432 16708 444438 16720
rect 447226 16708 447232 16720
rect 444432 16680 447232 16708
rect 444432 16668 444438 16680
rect 447226 16668 447232 16680
rect 447284 16668 447290 16720
rect 234890 16640 234896 16652
rect 234851 16612 234896 16640
rect 234890 16600 234896 16612
rect 234948 16600 234954 16652
rect 346394 16640 346400 16652
rect 346355 16612 346400 16640
rect 346394 16600 346400 16612
rect 346452 16600 346458 16652
rect 299842 15212 299848 15224
rect 299803 15184 299848 15212
rect 299842 15172 299848 15184
rect 299900 15172 299906 15224
rect 107470 15104 107476 15156
rect 107528 15144 107534 15156
rect 269206 15144 269212 15156
rect 107528 15116 269212 15144
rect 107528 15104 107534 15116
rect 269206 15104 269212 15116
rect 269264 15104 269270 15156
rect 103422 15036 103428 15088
rect 103480 15076 103486 15088
rect 267826 15076 267832 15088
rect 103480 15048 267832 15076
rect 103480 15036 103486 15048
rect 267826 15036 267832 15048
rect 267884 15036 267890 15088
rect 99282 14968 99288 15020
rect 99340 15008 99346 15020
rect 266446 15008 266452 15020
rect 99340 14980 266452 15008
rect 99340 14968 99346 14980
rect 266446 14968 266452 14980
rect 266504 14968 266510 15020
rect 96522 14900 96528 14952
rect 96580 14940 96586 14952
rect 265066 14940 265072 14952
rect 96580 14912 265072 14940
rect 96580 14900 96586 14912
rect 265066 14900 265072 14912
rect 265124 14900 265130 14952
rect 92382 14832 92388 14884
rect 92440 14872 92446 14884
rect 263686 14872 263692 14884
rect 92440 14844 263692 14872
rect 92440 14832 92446 14844
rect 263686 14832 263692 14844
rect 263744 14832 263750 14884
rect 89622 14764 89628 14816
rect 89680 14804 89686 14816
rect 262582 14804 262588 14816
rect 89680 14776 262588 14804
rect 89680 14764 89686 14776
rect 262582 14764 262588 14776
rect 262640 14764 262646 14816
rect 85482 14696 85488 14748
rect 85540 14736 85546 14748
rect 261110 14736 261116 14748
rect 85540 14708 261116 14736
rect 85540 14696 85546 14708
rect 261110 14696 261116 14708
rect 261168 14696 261174 14748
rect 82722 14628 82728 14680
rect 82780 14668 82786 14680
rect 259546 14668 259552 14680
rect 82780 14640 259552 14668
rect 82780 14628 82786 14640
rect 259546 14628 259552 14640
rect 259604 14628 259610 14680
rect 78582 14560 78588 14612
rect 78640 14600 78646 14612
rect 258166 14600 258172 14612
rect 78640 14572 258172 14600
rect 78640 14560 78646 14572
rect 258166 14560 258172 14572
rect 258224 14560 258230 14612
rect 74442 14492 74448 14544
rect 74500 14532 74506 14544
rect 256786 14532 256792 14544
rect 74500 14504 256792 14532
rect 74500 14492 74506 14504
rect 256786 14492 256792 14504
rect 256844 14492 256850 14544
rect 31662 14424 31668 14476
rect 31720 14464 31726 14476
rect 241698 14464 241704 14476
rect 31720 14436 241704 14464
rect 31720 14424 31726 14436
rect 241698 14424 241704 14436
rect 241756 14424 241762 14476
rect 110322 14356 110328 14408
rect 110380 14396 110386 14408
rect 270586 14396 270592 14408
rect 110380 14368 270592 14396
rect 110380 14356 110386 14368
rect 270586 14356 270592 14368
rect 270644 14356 270650 14408
rect 114462 14288 114468 14340
rect 114520 14328 114526 14340
rect 271966 14328 271972 14340
rect 114520 14300 271972 14328
rect 114520 14288 114526 14300
rect 271966 14288 271972 14300
rect 272024 14288 272030 14340
rect 117222 14220 117228 14272
rect 117280 14260 117286 14272
rect 273346 14260 273352 14272
rect 117280 14232 273352 14260
rect 117280 14220 117286 14232
rect 273346 14220 273352 14232
rect 273404 14220 273410 14272
rect 121362 14152 121368 14204
rect 121420 14192 121426 14204
rect 274726 14192 274732 14204
rect 121420 14164 274732 14192
rect 121420 14152 121426 14164
rect 274726 14152 274732 14164
rect 274784 14152 274790 14204
rect 125410 14084 125416 14136
rect 125468 14124 125474 14136
rect 276106 14124 276112 14136
rect 125468 14096 276112 14124
rect 125468 14084 125474 14096
rect 276106 14084 276112 14096
rect 276164 14084 276170 14136
rect 197262 14016 197268 14068
rect 197320 14056 197326 14068
rect 303890 14056 303896 14068
rect 197320 14028 303896 14056
rect 197320 14016 197326 14028
rect 303890 14016 303896 14028
rect 303948 14016 303954 14068
rect 190362 13744 190368 13796
rect 190420 13784 190426 13796
rect 301038 13784 301044 13796
rect 190420 13756 301044 13784
rect 190420 13744 190426 13756
rect 301038 13744 301044 13756
rect 301096 13744 301102 13796
rect 186222 13676 186228 13728
rect 186280 13716 186286 13728
rect 299658 13716 299664 13728
rect 186280 13688 299664 13716
rect 186280 13676 186286 13688
rect 299658 13676 299664 13688
rect 299716 13676 299722 13728
rect 183462 13608 183468 13660
rect 183520 13648 183526 13660
rect 298278 13648 298284 13660
rect 183520 13620 298284 13648
rect 183520 13608 183526 13620
rect 298278 13608 298284 13620
rect 298336 13608 298342 13660
rect 179322 13540 179328 13592
rect 179380 13580 179386 13592
rect 296990 13580 296996 13592
rect 179380 13552 296996 13580
rect 179380 13540 179386 13552
rect 296990 13540 296996 13552
rect 297048 13540 297054 13592
rect 176562 13472 176568 13524
rect 176620 13512 176626 13524
rect 295610 13512 295616 13524
rect 176620 13484 295616 13512
rect 176620 13472 176626 13484
rect 295610 13472 295616 13484
rect 295668 13472 295674 13524
rect 172422 13404 172428 13456
rect 172480 13444 172486 13456
rect 294230 13444 294236 13456
rect 172480 13416 294236 13444
rect 172480 13404 172486 13416
rect 294230 13404 294236 13416
rect 294288 13404 294294 13456
rect 160002 13336 160008 13388
rect 160060 13376 160066 13388
rect 288710 13376 288716 13388
rect 160060 13348 288716 13376
rect 160060 13336 160066 13348
rect 288710 13336 288716 13348
rect 288768 13336 288774 13388
rect 155862 13268 155868 13320
rect 155920 13308 155926 13320
rect 287330 13308 287336 13320
rect 155920 13280 287336 13308
rect 155920 13268 155926 13280
rect 287330 13268 287336 13280
rect 287388 13268 287394 13320
rect 135162 13200 135168 13252
rect 135220 13240 135226 13252
rect 280338 13240 280344 13252
rect 135220 13212 280344 13240
rect 135220 13200 135226 13212
rect 280338 13200 280344 13212
rect 280396 13200 280402 13252
rect 71682 13132 71688 13184
rect 71740 13172 71746 13184
rect 255406 13172 255412 13184
rect 71740 13144 255412 13172
rect 71740 13132 71746 13144
rect 255406 13132 255412 13144
rect 255464 13132 255470 13184
rect 23382 13064 23388 13116
rect 23440 13104 23446 13116
rect 237466 13104 237472 13116
rect 23440 13076 237472 13104
rect 23440 13064 23446 13076
rect 237466 13064 237472 13076
rect 237524 13064 237530 13116
rect 194502 12996 194508 13048
rect 194560 13036 194566 13048
rect 302418 13036 302424 13048
rect 194560 13008 302424 13036
rect 194560 12996 194566 13008
rect 302418 12996 302424 13008
rect 302476 12996 302482 13048
rect 211062 12928 211068 12980
rect 211120 12968 211126 12980
rect 308125 12971 308183 12977
rect 308125 12968 308137 12971
rect 211120 12940 308137 12968
rect 211120 12928 211126 12940
rect 308125 12937 308137 12940
rect 308171 12937 308183 12971
rect 308125 12931 308183 12937
rect 213822 12860 213828 12912
rect 213880 12900 213886 12912
rect 309318 12900 309324 12912
rect 213880 12872 309324 12900
rect 213880 12860 213886 12872
rect 309318 12860 309324 12872
rect 309376 12860 309382 12912
rect 217962 12792 217968 12844
rect 218020 12832 218026 12844
rect 310698 12832 310704 12844
rect 218020 12804 310704 12832
rect 218020 12792 218026 12804
rect 310698 12792 310704 12804
rect 310756 12792 310762 12844
rect 220722 12724 220728 12776
rect 220780 12764 220786 12776
rect 312170 12764 312176 12776
rect 220780 12736 312176 12764
rect 220780 12724 220786 12736
rect 312170 12724 312176 12736
rect 312228 12724 312234 12776
rect 224862 12656 224868 12708
rect 224920 12696 224926 12708
rect 313550 12696 313556 12708
rect 224920 12668 313556 12696
rect 224920 12656 224926 12668
rect 313550 12656 313556 12668
rect 313608 12656 313614 12708
rect 229002 12588 229008 12640
rect 229060 12628 229066 12640
rect 314930 12628 314936 12640
rect 229060 12600 314936 12628
rect 229060 12588 229066 12600
rect 314930 12588 314936 12600
rect 314988 12588 314994 12640
rect 231305 12563 231363 12569
rect 231305 12529 231317 12563
rect 231351 12560 231363 12563
rect 316218 12560 316224 12572
rect 231351 12532 316224 12560
rect 231351 12529 231363 12532
rect 231305 12523 231363 12529
rect 316218 12520 316224 12532
rect 316276 12520 316282 12572
rect 234706 12492 234712 12504
rect 234667 12464 234712 12492
rect 234706 12452 234712 12464
rect 234764 12452 234770 12504
rect 290090 12492 290096 12504
rect 290051 12464 290096 12492
rect 290090 12452 290096 12464
rect 290148 12452 290154 12504
rect 325970 12492 325976 12504
rect 325896 12464 325976 12492
rect 325896 12436 325924 12464
rect 325970 12452 325976 12464
rect 326028 12452 326034 12504
rect 173802 12384 173808 12436
rect 173860 12424 173866 12436
rect 294046 12424 294052 12436
rect 173860 12396 294052 12424
rect 173860 12384 173866 12396
rect 294046 12384 294052 12396
rect 294104 12384 294110 12436
rect 325878 12384 325884 12436
rect 325936 12384 325942 12436
rect 169386 12316 169392 12368
rect 169444 12356 169450 12368
rect 292942 12356 292948 12368
rect 169444 12328 292948 12356
rect 169444 12316 169450 12328
rect 292942 12316 292948 12328
rect 293000 12316 293006 12368
rect 328457 12359 328515 12365
rect 328457 12325 328469 12359
rect 328503 12356 328515 12359
rect 328546 12356 328552 12368
rect 328503 12328 328552 12356
rect 328503 12325 328515 12328
rect 328457 12319 328515 12325
rect 328546 12316 328552 12328
rect 328604 12316 328610 12368
rect 165890 12248 165896 12300
rect 165948 12288 165954 12300
rect 291654 12288 291660 12300
rect 165948 12260 291660 12288
rect 165948 12248 165954 12260
rect 291654 12248 291660 12260
rect 291712 12248 291718 12300
rect 162302 12180 162308 12232
rect 162360 12220 162366 12232
rect 290093 12223 290151 12229
rect 290093 12220 290105 12223
rect 162360 12192 290105 12220
rect 162360 12180 162366 12192
rect 290093 12189 290105 12192
rect 290139 12189 290151 12223
rect 290093 12183 290151 12189
rect 151722 12112 151728 12164
rect 151780 12152 151786 12164
rect 285858 12152 285864 12164
rect 151780 12124 285864 12152
rect 151780 12112 151786 12124
rect 285858 12112 285864 12124
rect 285916 12112 285922 12164
rect 148962 12044 148968 12096
rect 149020 12084 149026 12096
rect 285950 12084 285956 12096
rect 149020 12056 285956 12084
rect 149020 12044 149026 12056
rect 285950 12044 285956 12056
rect 286008 12044 286014 12096
rect 144822 11976 144828 12028
rect 144880 12016 144886 12028
rect 284478 12016 284484 12028
rect 144880 11988 284484 12016
rect 144880 11976 144886 11988
rect 284478 11976 284484 11988
rect 284536 11976 284542 12028
rect 140866 11908 140872 11960
rect 140924 11948 140930 11960
rect 283098 11948 283104 11960
rect 140924 11920 283104 11948
rect 140924 11908 140930 11920
rect 283098 11908 283104 11920
rect 283156 11908 283162 11960
rect 128262 11840 128268 11892
rect 128320 11880 128326 11892
rect 277486 11880 277492 11892
rect 128320 11852 277492 11880
rect 128320 11840 128326 11852
rect 277486 11840 277492 11852
rect 277544 11840 277550 11892
rect 126882 11772 126888 11824
rect 126940 11812 126946 11824
rect 277578 11812 277584 11824
rect 126940 11784 277584 11812
rect 126940 11772 126946 11784
rect 277578 11772 277584 11784
rect 277636 11772 277642 11824
rect 18322 11704 18328 11756
rect 18380 11744 18386 11756
rect 236086 11744 236092 11756
rect 18380 11716 236092 11744
rect 18380 11704 18386 11716
rect 236086 11704 236092 11716
rect 236144 11704 236150 11756
rect 176378 11636 176384 11688
rect 176436 11676 176442 11688
rect 295426 11676 295432 11688
rect 176436 11648 295432 11676
rect 176436 11636 176442 11648
rect 295426 11636 295432 11648
rect 295484 11636 295490 11688
rect 180702 11568 180708 11620
rect 180760 11608 180766 11620
rect 296806 11608 296812 11620
rect 180760 11580 296812 11608
rect 180760 11568 180766 11580
rect 296806 11568 296812 11580
rect 296864 11568 296870 11620
rect 184750 11500 184756 11552
rect 184808 11540 184814 11552
rect 298646 11540 298652 11552
rect 184808 11512 298652 11540
rect 184808 11500 184814 11512
rect 298646 11500 298652 11512
rect 298704 11500 298710 11552
rect 187602 11432 187608 11484
rect 187660 11472 187666 11484
rect 299842 11472 299848 11484
rect 187660 11444 299848 11472
rect 187660 11432 187666 11444
rect 299842 11432 299848 11444
rect 299900 11432 299906 11484
rect 191742 11364 191748 11416
rect 191800 11404 191806 11416
rect 300946 11404 300952 11416
rect 191800 11376 300952 11404
rect 191800 11364 191806 11376
rect 300946 11364 300952 11376
rect 301004 11364 301010 11416
rect 194410 11296 194416 11348
rect 194468 11336 194474 11348
rect 302326 11336 302332 11348
rect 194468 11308 302332 11336
rect 194468 11296 194474 11308
rect 302326 11296 302332 11308
rect 302384 11296 302390 11348
rect 198642 11228 198648 11280
rect 198700 11268 198706 11280
rect 303798 11268 303804 11280
rect 198700 11240 303804 11268
rect 198700 11228 198706 11240
rect 303798 11228 303804 11240
rect 303856 11228 303862 11280
rect 234706 11200 234712 11212
rect 234667 11172 234712 11200
rect 234706 11160 234712 11172
rect 234764 11160 234770 11212
rect 108942 10956 108948 11008
rect 109000 10996 109006 11008
rect 270678 10996 270684 11008
rect 109000 10968 270684 10996
rect 109000 10956 109006 10968
rect 270678 10956 270684 10968
rect 270736 10956 270742 11008
rect 106182 10888 106188 10940
rect 106240 10928 106246 10940
rect 269298 10928 269304 10940
rect 106240 10900 269304 10928
rect 106240 10888 106246 10900
rect 269298 10888 269304 10900
rect 269356 10888 269362 10940
rect 102042 10820 102048 10872
rect 102100 10860 102106 10872
rect 267918 10860 267924 10872
rect 102100 10832 267924 10860
rect 102100 10820 102106 10832
rect 267918 10820 267924 10832
rect 267976 10820 267982 10872
rect 99190 10752 99196 10804
rect 99248 10792 99254 10804
rect 266538 10792 266544 10804
rect 99248 10764 266544 10792
rect 99248 10752 99254 10764
rect 266538 10752 266544 10764
rect 266596 10752 266602 10804
rect 95142 10684 95148 10736
rect 95200 10724 95206 10736
rect 265158 10724 265164 10736
rect 95200 10696 265164 10724
rect 95200 10684 95206 10696
rect 265158 10684 265164 10696
rect 265216 10684 265222 10736
rect 91002 10616 91008 10668
rect 91060 10656 91066 10668
rect 263778 10656 263784 10668
rect 91060 10628 263784 10656
rect 91060 10616 91066 10628
rect 263778 10616 263784 10628
rect 263836 10616 263842 10668
rect 63586 10548 63592 10600
rect 63644 10588 63650 10600
rect 252646 10588 252652 10600
rect 63644 10560 252652 10588
rect 63644 10548 63650 10560
rect 252646 10548 252652 10560
rect 252704 10548 252710 10600
rect 59998 10480 60004 10532
rect 60056 10520 60062 10532
rect 251266 10520 251272 10532
rect 60056 10492 251272 10520
rect 60056 10480 60062 10492
rect 251266 10480 251272 10492
rect 251324 10480 251330 10532
rect 56410 10412 56416 10464
rect 56468 10452 56474 10464
rect 249886 10452 249892 10464
rect 56468 10424 249892 10452
rect 56468 10412 56474 10424
rect 249886 10412 249892 10424
rect 249944 10412 249950 10464
rect 52822 10344 52828 10396
rect 52880 10384 52886 10396
rect 248598 10384 248604 10396
rect 52880 10356 248604 10384
rect 52880 10344 52886 10356
rect 248598 10344 248604 10356
rect 248656 10344 248662 10396
rect 49326 10276 49332 10328
rect 49384 10316 49390 10328
rect 248506 10316 248512 10328
rect 49384 10288 248512 10316
rect 49384 10276 49390 10288
rect 248506 10276 248512 10288
rect 248564 10276 248570 10328
rect 113082 10208 113088 10260
rect 113140 10248 113146 10260
rect 272058 10248 272064 10260
rect 113140 10220 272064 10248
rect 113140 10208 113146 10220
rect 272058 10208 272064 10220
rect 272116 10208 272122 10260
rect 117130 10140 117136 10192
rect 117188 10180 117194 10192
rect 273438 10180 273444 10192
rect 117188 10152 273444 10180
rect 117188 10140 117194 10152
rect 273438 10140 273444 10152
rect 273496 10140 273502 10192
rect 119982 10072 119988 10124
rect 120040 10112 120046 10124
rect 274818 10112 274824 10124
rect 120040 10084 274824 10112
rect 120040 10072 120046 10084
rect 274818 10072 274824 10084
rect 274876 10072 274882 10124
rect 124122 10004 124128 10056
rect 124180 10044 124186 10056
rect 276198 10044 276204 10056
rect 124180 10016 276204 10044
rect 124180 10004 124186 10016
rect 276198 10004 276204 10016
rect 276256 10004 276262 10056
rect 154482 9936 154488 9988
rect 154540 9976 154546 9988
rect 287146 9976 287152 9988
rect 154540 9948 287152 9976
rect 154540 9936 154546 9948
rect 287146 9936 287152 9948
rect 287204 9936 287210 9988
rect 158622 9868 158628 9920
rect 158680 9908 158686 9920
rect 288526 9908 288532 9920
rect 158680 9880 288532 9908
rect 158680 9868 158686 9880
rect 288526 9868 288532 9880
rect 288584 9868 288590 9920
rect 161382 9800 161388 9852
rect 161440 9840 161446 9852
rect 289906 9840 289912 9852
rect 161440 9812 289912 9840
rect 161440 9800 161446 9812
rect 289906 9800 289912 9812
rect 289964 9800 289970 9852
rect 231302 9704 231308 9716
rect 231263 9676 231308 9704
rect 231302 9664 231308 9676
rect 231360 9664 231366 9716
rect 252738 9704 252744 9716
rect 252699 9676 252744 9704
rect 252738 9664 252744 9676
rect 252796 9664 252802 9716
rect 254118 9704 254124 9716
rect 254079 9676 254124 9704
rect 254118 9664 254124 9676
rect 254176 9664 254182 9716
rect 327258 9704 327264 9716
rect 327219 9676 327264 9704
rect 327258 9664 327264 9676
rect 327316 9664 327322 9716
rect 342438 9704 342444 9716
rect 342399 9676 342444 9704
rect 342438 9664 342444 9676
rect 342496 9664 342502 9716
rect 345198 9704 345204 9716
rect 345159 9676 345204 9704
rect 345198 9664 345204 9676
rect 345256 9664 345262 9716
rect 363230 9704 363236 9716
rect 363191 9676 363236 9704
rect 363230 9664 363236 9676
rect 363288 9664 363294 9716
rect 203886 9596 203892 9648
rect 203944 9636 203950 9648
rect 306558 9636 306564 9648
rect 203944 9608 306564 9636
rect 203944 9596 203950 9608
rect 306558 9596 306564 9608
rect 306616 9596 306622 9648
rect 405550 9596 405556 9648
rect 405608 9636 405614 9648
rect 463234 9636 463240 9648
rect 405608 9608 463240 9636
rect 405608 9596 405614 9608
rect 463234 9596 463240 9608
rect 463292 9596 463298 9648
rect 200390 9528 200396 9580
rect 200448 9568 200454 9580
rect 305086 9568 305092 9580
rect 200448 9540 305092 9568
rect 200448 9528 200454 9540
rect 305086 9528 305092 9540
rect 305144 9528 305150 9580
rect 406930 9528 406936 9580
rect 406988 9568 406994 9580
rect 466822 9568 466828 9580
rect 406988 9540 466828 9568
rect 406988 9528 406994 9540
rect 466822 9528 466828 9540
rect 466880 9528 466886 9580
rect 150434 9460 150440 9512
rect 150492 9500 150498 9512
rect 285766 9500 285772 9512
rect 150492 9472 285772 9500
rect 150492 9460 150498 9472
rect 285766 9460 285772 9472
rect 285824 9460 285830 9512
rect 408310 9460 408316 9512
rect 408368 9500 408374 9512
rect 470318 9500 470324 9512
rect 408368 9472 470324 9500
rect 408368 9460 408374 9472
rect 470318 9460 470324 9472
rect 470376 9460 470382 9512
rect 146846 9392 146852 9444
rect 146904 9432 146910 9444
rect 284386 9432 284392 9444
rect 146904 9404 284392 9432
rect 146904 9392 146910 9404
rect 284386 9392 284392 9404
rect 284444 9392 284450 9444
rect 439958 9392 439964 9444
rect 440016 9432 440022 9444
rect 555970 9432 555976 9444
rect 440016 9404 555976 9432
rect 440016 9392 440022 9404
rect 555970 9392 555976 9404
rect 556028 9392 556034 9444
rect 143258 9324 143264 9376
rect 143316 9364 143322 9376
rect 283006 9364 283012 9376
rect 143316 9336 283012 9364
rect 143316 9324 143322 9336
rect 283006 9324 283012 9336
rect 283064 9324 283070 9376
rect 441430 9324 441436 9376
rect 441488 9364 441494 9376
rect 559558 9364 559564 9376
rect 441488 9336 559564 9364
rect 441488 9324 441494 9336
rect 559558 9324 559564 9336
rect 559616 9324 559622 9376
rect 139670 9256 139676 9308
rect 139728 9296 139734 9308
rect 281718 9296 281724 9308
rect 139728 9268 281724 9296
rect 139728 9256 139734 9268
rect 281718 9256 281724 9268
rect 281776 9256 281782 9308
rect 442718 9256 442724 9308
rect 442776 9296 442782 9308
rect 563146 9296 563152 9308
rect 442776 9268 563152 9296
rect 442776 9256 442782 9268
rect 563146 9256 563152 9268
rect 563204 9256 563210 9308
rect 136082 9188 136088 9240
rect 136140 9228 136146 9240
rect 280430 9228 280436 9240
rect 136140 9200 280436 9228
rect 136140 9188 136146 9200
rect 280430 9188 280436 9200
rect 280488 9188 280494 9240
rect 444006 9188 444012 9240
rect 444064 9228 444070 9240
rect 566734 9228 566740 9240
rect 444064 9200 566740 9228
rect 444064 9188 444070 9200
rect 566734 9188 566740 9200
rect 566792 9188 566798 9240
rect 44542 9120 44548 9172
rect 44600 9160 44606 9172
rect 245746 9160 245752 9172
rect 44600 9132 245752 9160
rect 44600 9120 44606 9132
rect 245746 9120 245752 9132
rect 245804 9120 245810 9172
rect 250346 9120 250352 9172
rect 250404 9160 250410 9172
rect 323210 9160 323216 9172
rect 250404 9132 323216 9160
rect 250404 9120 250410 9132
rect 323210 9120 323216 9132
rect 323268 9120 323274 9172
rect 445478 9120 445484 9172
rect 445536 9160 445542 9172
rect 570230 9160 570236 9172
rect 445536 9132 570236 9160
rect 445536 9120 445542 9132
rect 570230 9120 570236 9132
rect 570288 9120 570294 9172
rect 40954 9052 40960 9104
rect 41012 9092 41018 9104
rect 244458 9092 244464 9104
rect 41012 9064 244464 9092
rect 41012 9052 41018 9064
rect 244458 9052 244464 9064
rect 244516 9052 244522 9104
rect 246758 9052 246764 9104
rect 246816 9092 246822 9104
rect 323118 9092 323124 9104
rect 246816 9064 323124 9092
rect 246816 9052 246822 9064
rect 323118 9052 323124 9064
rect 323176 9052 323182 9104
rect 446950 9052 446956 9104
rect 447008 9092 447014 9104
rect 573818 9092 573824 9104
rect 447008 9064 573824 9092
rect 447008 9052 447014 9064
rect 573818 9052 573824 9064
rect 573876 9052 573882 9104
rect 27890 8984 27896 9036
rect 27948 9024 27954 9036
rect 233878 9024 233884 9036
rect 27948 8996 233884 9024
rect 27948 8984 27954 8996
rect 233878 8984 233884 8996
rect 233936 8984 233942 9036
rect 239582 8984 239588 9036
rect 239640 9024 239646 9036
rect 320358 9024 320364 9036
rect 239640 8996 320364 9024
rect 239640 8984 239646 8996
rect 320358 8984 320364 8996
rect 320416 8984 320422 9036
rect 448330 8984 448336 9036
rect 448388 9024 448394 9036
rect 577406 9024 577412 9036
rect 448388 8996 577412 9024
rect 448388 8984 448394 8996
rect 577406 8984 577412 8996
rect 577464 8984 577470 9036
rect 13630 8916 13636 8968
rect 13688 8956 13694 8968
rect 234801 8959 234859 8965
rect 234801 8956 234813 8959
rect 13688 8928 234813 8956
rect 13688 8916 13694 8928
rect 234801 8925 234813 8928
rect 234847 8925 234859 8959
rect 234801 8919 234859 8925
rect 235994 8916 236000 8968
rect 236052 8956 236058 8968
rect 318978 8956 318984 8968
rect 236052 8928 318984 8956
rect 236052 8916 236058 8928
rect 318978 8916 318984 8928
rect 319036 8916 319042 8968
rect 400030 8916 400036 8968
rect 400088 8956 400094 8968
rect 448974 8956 448980 8968
rect 400088 8928 448980 8956
rect 400088 8916 400094 8928
rect 448974 8916 448980 8928
rect 449032 8916 449038 8968
rect 449710 8916 449716 8968
rect 449768 8956 449774 8968
rect 580994 8956 581000 8968
rect 449768 8928 581000 8956
rect 449768 8916 449774 8928
rect 580994 8916 581000 8928
rect 581052 8916 581058 8968
rect 207474 8848 207480 8900
rect 207532 8888 207538 8900
rect 307846 8888 307852 8900
rect 207532 8860 307852 8888
rect 207532 8848 207538 8860
rect 307846 8848 307852 8860
rect 307904 8848 307910 8900
rect 404170 8848 404176 8900
rect 404228 8888 404234 8900
rect 459646 8888 459652 8900
rect 404228 8860 459652 8888
rect 404228 8848 404234 8860
rect 459646 8848 459652 8860
rect 459704 8848 459710 8900
rect 210878 8780 210884 8832
rect 210936 8820 210942 8832
rect 309226 8820 309232 8832
rect 210936 8792 309232 8820
rect 210936 8780 210942 8792
rect 309226 8780 309232 8792
rect 309284 8780 309290 8832
rect 402790 8780 402796 8832
rect 402848 8820 402854 8832
rect 456058 8820 456064 8832
rect 402848 8792 456064 8820
rect 402848 8780 402854 8792
rect 456058 8780 456064 8792
rect 456116 8780 456122 8832
rect 214650 8712 214656 8764
rect 214708 8752 214714 8764
rect 310606 8752 310612 8764
rect 214708 8724 310612 8752
rect 214708 8712 214714 8724
rect 310606 8712 310612 8724
rect 310664 8712 310670 8764
rect 401410 8712 401416 8764
rect 401468 8752 401474 8764
rect 452470 8752 452476 8764
rect 401468 8724 452476 8752
rect 401468 8712 401474 8724
rect 452470 8712 452476 8724
rect 452528 8712 452534 8764
rect 218146 8644 218152 8696
rect 218204 8684 218210 8696
rect 311986 8684 311992 8696
rect 218204 8656 311992 8684
rect 218204 8644 218210 8656
rect 311986 8644 311992 8656
rect 312044 8644 312050 8696
rect 221734 8576 221740 8628
rect 221792 8616 221798 8628
rect 313366 8616 313372 8628
rect 221792 8588 313372 8616
rect 221792 8576 221798 8588
rect 313366 8576 313372 8588
rect 313424 8576 313430 8628
rect 225322 8508 225328 8560
rect 225380 8548 225386 8560
rect 314746 8548 314752 8560
rect 225380 8520 314752 8548
rect 225380 8508 225386 8520
rect 314746 8508 314752 8520
rect 314804 8508 314810 8560
rect 228910 8440 228916 8492
rect 228968 8480 228974 8492
rect 316126 8480 316132 8492
rect 228968 8452 316132 8480
rect 228968 8440 228974 8452
rect 316126 8440 316132 8452
rect 316184 8440 316190 8492
rect 232498 8372 232504 8424
rect 232556 8412 232562 8424
rect 317598 8412 317604 8424
rect 232556 8384 317604 8412
rect 232556 8372 232562 8384
rect 317598 8372 317604 8384
rect 317656 8372 317662 8424
rect 229186 8344 229192 8356
rect 229147 8316 229192 8344
rect 229186 8304 229192 8316
rect 229244 8304 229250 8356
rect 234890 8304 234896 8356
rect 234948 8344 234954 8356
rect 235074 8344 235080 8356
rect 234948 8316 235080 8344
rect 234948 8304 234954 8316
rect 235074 8304 235080 8316
rect 235132 8304 235138 8356
rect 238941 8347 238999 8353
rect 238941 8313 238953 8347
rect 238987 8344 238999 8347
rect 239030 8344 239036 8356
rect 238987 8316 239036 8344
rect 238987 8313 238999 8316
rect 238941 8307 238999 8313
rect 239030 8304 239036 8316
rect 239088 8304 239094 8356
rect 240226 8344 240232 8356
rect 240187 8316 240232 8344
rect 240226 8304 240232 8316
rect 240284 8304 240290 8356
rect 241609 8347 241667 8353
rect 241609 8313 241621 8347
rect 241655 8344 241667 8347
rect 241698 8344 241704 8356
rect 241655 8316 241704 8344
rect 241655 8313 241667 8316
rect 241609 8307 241667 8313
rect 241698 8304 241704 8316
rect 241756 8304 241762 8356
rect 243170 8304 243176 8356
rect 243228 8344 243234 8356
rect 321738 8344 321744 8356
rect 243228 8316 321744 8344
rect 243228 8304 243234 8316
rect 321738 8304 321744 8316
rect 321796 8304 321802 8356
rect 128998 8236 129004 8288
rect 129056 8276 129062 8288
rect 251177 8279 251235 8285
rect 251177 8276 251189 8279
rect 129056 8248 251189 8276
rect 129056 8236 129062 8248
rect 251177 8245 251189 8248
rect 251223 8245 251235 8279
rect 251177 8239 251235 8245
rect 254581 8279 254639 8285
rect 254581 8245 254593 8279
rect 254627 8276 254639 8279
rect 277394 8276 277400 8288
rect 254627 8248 277400 8276
rect 254627 8245 254639 8248
rect 254581 8239 254639 8245
rect 277394 8236 277400 8248
rect 277452 8236 277458 8288
rect 420730 8236 420736 8288
rect 420788 8276 420794 8288
rect 504818 8276 504824 8288
rect 420788 8248 504824 8276
rect 420788 8236 420794 8248
rect 504818 8236 504824 8248
rect 504876 8236 504882 8288
rect 87322 8168 87328 8220
rect 87380 8208 87386 8220
rect 262398 8208 262404 8220
rect 87380 8180 262404 8208
rect 87380 8168 87386 8180
rect 262398 8168 262404 8180
rect 262456 8168 262462 8220
rect 266998 8168 267004 8220
rect 267056 8208 267062 8220
rect 329926 8208 329932 8220
rect 267056 8180 329932 8208
rect 267056 8168 267062 8180
rect 329926 8168 329932 8180
rect 329984 8168 329990 8220
rect 391474 8168 391480 8220
rect 391532 8208 391538 8220
rect 391750 8208 391756 8220
rect 391532 8180 391756 8208
rect 391532 8168 391538 8180
rect 391750 8168 391756 8180
rect 391808 8168 391814 8220
rect 422110 8168 422116 8220
rect 422168 8208 422174 8220
rect 508406 8208 508412 8220
rect 422168 8180 508412 8208
rect 422168 8168 422174 8180
rect 508406 8168 508412 8180
rect 508464 8168 508470 8220
rect 83826 8100 83832 8152
rect 83884 8140 83890 8152
rect 261018 8140 261024 8152
rect 83884 8112 261024 8140
rect 83884 8100 83890 8112
rect 261018 8100 261024 8112
rect 261076 8100 261082 8152
rect 263410 8100 263416 8152
rect 263468 8140 263474 8152
rect 328454 8140 328460 8152
rect 263468 8112 328460 8140
rect 263468 8100 263474 8112
rect 328454 8100 328460 8112
rect 328512 8100 328518 8152
rect 427630 8100 427636 8152
rect 427688 8140 427694 8152
rect 523862 8140 523868 8152
rect 427688 8112 523868 8140
rect 427688 8100 427694 8112
rect 523862 8100 523868 8112
rect 523920 8100 523926 8152
rect 80238 8032 80244 8084
rect 80296 8072 80302 8084
rect 259730 8072 259736 8084
rect 80296 8044 259736 8072
rect 80296 8032 80302 8044
rect 259730 8032 259736 8044
rect 259788 8032 259794 8084
rect 259822 8032 259828 8084
rect 259880 8072 259886 8084
rect 327258 8072 327264 8084
rect 259880 8044 327264 8072
rect 259880 8032 259886 8044
rect 327258 8032 327264 8044
rect 327316 8032 327322 8084
rect 429010 8032 429016 8084
rect 429068 8072 429074 8084
rect 527450 8072 527456 8084
rect 429068 8044 527456 8072
rect 429068 8032 429074 8044
rect 527450 8032 527456 8044
rect 527508 8032 527514 8084
rect 37366 7964 37372 8016
rect 37424 8004 37430 8016
rect 243078 8004 243084 8016
rect 37424 7976 243084 8004
rect 37424 7964 37430 7976
rect 243078 7964 243084 7976
rect 243136 7964 243142 8016
rect 251177 8007 251235 8013
rect 251177 7973 251189 8007
rect 251223 8004 251235 8007
rect 254581 8007 254639 8013
rect 254581 8004 254593 8007
rect 251223 7976 254593 8004
rect 251223 7973 251235 7976
rect 251177 7967 251235 7973
rect 254581 7973 254593 7976
rect 254627 7973 254639 8007
rect 254581 7967 254639 7973
rect 256234 7964 256240 8016
rect 256292 8004 256298 8016
rect 325878 8004 325884 8016
rect 256292 7976 325884 8004
rect 256292 7964 256298 7976
rect 325878 7964 325884 7976
rect 325936 7964 325942 8016
rect 430390 7964 430396 8016
rect 430448 8004 430454 8016
rect 531038 8004 531044 8016
rect 430448 7976 531044 8004
rect 430448 7964 430454 7976
rect 531038 7964 531044 7976
rect 531096 7964 531102 8016
rect 33870 7896 33876 7948
rect 33928 7936 33934 7948
rect 241698 7936 241704 7948
rect 33928 7908 241704 7936
rect 33928 7896 33934 7908
rect 241698 7896 241704 7908
rect 241756 7896 241762 7948
rect 252646 7896 252652 7948
rect 252704 7936 252710 7948
rect 324590 7936 324596 7948
rect 252704 7908 324596 7936
rect 252704 7896 252710 7908
rect 324590 7896 324596 7908
rect 324648 7896 324654 7948
rect 431770 7896 431776 7948
rect 431828 7936 431834 7948
rect 534534 7936 534540 7948
rect 431828 7908 534540 7936
rect 431828 7896 431834 7908
rect 534534 7896 534540 7908
rect 534592 7896 534598 7948
rect 30282 7828 30288 7880
rect 30340 7868 30346 7880
rect 240226 7868 240232 7880
rect 30340 7840 240232 7868
rect 30340 7828 30346 7840
rect 240226 7828 240232 7840
rect 240284 7828 240290 7880
rect 249150 7828 249156 7880
rect 249208 7868 249214 7880
rect 323026 7868 323032 7880
rect 249208 7840 323032 7868
rect 249208 7828 249214 7840
rect 323026 7828 323032 7840
rect 323084 7828 323090 7880
rect 433150 7828 433156 7880
rect 433208 7868 433214 7880
rect 538122 7868 538128 7880
rect 433208 7840 538128 7868
rect 433208 7828 433214 7840
rect 538122 7828 538128 7840
rect 538180 7828 538186 7880
rect 26694 7760 26700 7812
rect 26752 7800 26758 7812
rect 239030 7800 239036 7812
rect 26752 7772 239036 7800
rect 26752 7760 26758 7772
rect 239030 7760 239036 7772
rect 239088 7760 239094 7812
rect 245562 7760 245568 7812
rect 245620 7800 245626 7812
rect 321646 7800 321652 7812
rect 245620 7772 321652 7800
rect 245620 7760 245626 7772
rect 321646 7760 321652 7772
rect 321704 7760 321710 7812
rect 434530 7760 434536 7812
rect 434588 7800 434594 7812
rect 541710 7800 541716 7812
rect 434588 7772 541716 7800
rect 434588 7760 434594 7772
rect 541710 7760 541716 7772
rect 541768 7760 541774 7812
rect 21910 7692 21916 7744
rect 21968 7732 21974 7744
rect 237650 7732 237656 7744
rect 21968 7704 237656 7732
rect 21968 7692 21974 7704
rect 237650 7692 237656 7704
rect 237708 7692 237714 7744
rect 241974 7692 241980 7744
rect 242032 7732 242038 7744
rect 320266 7732 320272 7744
rect 242032 7704 320272 7732
rect 242032 7692 242038 7704
rect 320266 7692 320272 7704
rect 320324 7692 320330 7744
rect 435910 7692 435916 7744
rect 435968 7732 435974 7744
rect 545298 7732 545304 7744
rect 435968 7704 545304 7732
rect 435968 7692 435974 7704
rect 545298 7692 545304 7704
rect 545356 7692 545362 7744
rect 17218 7624 17224 7676
rect 17276 7664 17282 7676
rect 236178 7664 236184 7676
rect 17276 7636 236184 7664
rect 17276 7624 17282 7636
rect 236178 7624 236184 7636
rect 236236 7624 236242 7676
rect 238386 7624 238392 7676
rect 238444 7664 238450 7676
rect 319162 7664 319168 7676
rect 238444 7636 319168 7664
rect 238444 7624 238450 7636
rect 319162 7624 319168 7636
rect 319220 7624 319226 7676
rect 437290 7624 437296 7676
rect 437348 7664 437354 7676
rect 548886 7664 548892 7676
rect 437348 7636 548892 7664
rect 437348 7624 437354 7636
rect 548886 7624 548892 7636
rect 548944 7624 548950 7676
rect 8846 7556 8852 7608
rect 8904 7596 8910 7608
rect 227625 7599 227683 7605
rect 227625 7596 227637 7599
rect 8904 7568 227637 7596
rect 8904 7556 8910 7568
rect 227625 7565 227637 7568
rect 227671 7565 227683 7599
rect 227625 7559 227683 7565
rect 227714 7556 227720 7608
rect 227772 7596 227778 7608
rect 229002 7596 229008 7608
rect 227772 7568 229008 7596
rect 227772 7556 227778 7568
rect 229002 7556 229008 7568
rect 229060 7556 229066 7608
rect 234798 7556 234804 7608
rect 234856 7596 234862 7608
rect 317782 7596 317788 7608
rect 234856 7568 317788 7596
rect 234856 7556 234862 7568
rect 317782 7556 317788 7568
rect 317840 7556 317846 7608
rect 438670 7556 438676 7608
rect 438728 7596 438734 7608
rect 552382 7596 552388 7608
rect 438728 7568 552388 7596
rect 438728 7556 438734 7568
rect 552382 7556 552388 7568
rect 552440 7556 552446 7608
rect 138474 7488 138480 7540
rect 138532 7528 138538 7540
rect 281810 7528 281816 7540
rect 138532 7500 281816 7528
rect 138532 7488 138538 7500
rect 281810 7488 281816 7500
rect 281868 7488 281874 7540
rect 419350 7488 419356 7540
rect 419408 7528 419414 7540
rect 501230 7528 501236 7540
rect 419408 7500 501236 7528
rect 419408 7488 419414 7500
rect 501230 7488 501236 7500
rect 501288 7488 501294 7540
rect 142062 7420 142068 7472
rect 142120 7460 142126 7472
rect 283190 7460 283196 7472
rect 142120 7432 283196 7460
rect 142120 7420 142126 7432
rect 283190 7420 283196 7432
rect 283248 7420 283254 7472
rect 417970 7420 417976 7472
rect 418028 7460 418034 7472
rect 497734 7460 497740 7472
rect 418028 7432 497740 7460
rect 418028 7420 418034 7432
rect 497734 7420 497740 7432
rect 497792 7420 497798 7472
rect 145650 7352 145656 7404
rect 145708 7392 145714 7404
rect 284570 7392 284576 7404
rect 145708 7364 284576 7392
rect 145708 7352 145714 7364
rect 284570 7352 284576 7364
rect 284628 7352 284634 7404
rect 416498 7352 416504 7404
rect 416556 7392 416562 7404
rect 494146 7392 494152 7404
rect 416556 7364 494152 7392
rect 416556 7352 416562 7364
rect 494146 7352 494152 7364
rect 494204 7352 494210 7404
rect 149238 7284 149244 7336
rect 149296 7324 149302 7336
rect 286042 7324 286048 7336
rect 149296 7296 286048 7324
rect 149296 7284 149302 7296
rect 286042 7284 286048 7296
rect 286100 7284 286106 7336
rect 415210 7284 415216 7336
rect 415268 7324 415274 7336
rect 490558 7324 490564 7336
rect 415268 7296 490564 7324
rect 415268 7284 415274 7296
rect 490558 7284 490564 7296
rect 490616 7284 490622 7336
rect 152734 7216 152740 7268
rect 152792 7256 152798 7268
rect 287054 7256 287060 7268
rect 152792 7228 287060 7256
rect 152792 7216 152798 7228
rect 287054 7216 287060 7228
rect 287112 7216 287118 7268
rect 413830 7216 413836 7268
rect 413888 7256 413894 7268
rect 486970 7256 486976 7268
rect 413888 7228 486976 7256
rect 413888 7216 413894 7228
rect 486970 7216 486976 7228
rect 487028 7216 487034 7268
rect 156322 7148 156328 7200
rect 156380 7188 156386 7200
rect 288434 7188 288440 7200
rect 156380 7160 288440 7188
rect 156380 7148 156386 7160
rect 288434 7148 288440 7160
rect 288492 7148 288498 7200
rect 412542 7148 412548 7200
rect 412600 7188 412606 7200
rect 483474 7188 483480 7200
rect 412600 7160 483480 7188
rect 412600 7148 412606 7160
rect 483474 7148 483480 7160
rect 483532 7148 483538 7200
rect 158714 7080 158720 7132
rect 158772 7120 158778 7132
rect 160002 7120 160008 7132
rect 158772 7092 160008 7120
rect 158772 7080 158778 7092
rect 160002 7080 160008 7092
rect 160060 7080 160066 7132
rect 289814 7120 289820 7132
rect 160112 7092 289820 7120
rect 159910 7012 159916 7064
rect 159968 7052 159974 7064
rect 160112 7052 160140 7092
rect 289814 7080 289820 7092
rect 289872 7080 289878 7132
rect 398558 7080 398564 7132
rect 398616 7120 398622 7132
rect 445386 7120 445392 7132
rect 398616 7092 445392 7120
rect 398616 7080 398622 7092
rect 445386 7080 445392 7092
rect 445444 7080 445450 7132
rect 159968 7024 160140 7052
rect 159968 7012 159974 7024
rect 164694 7012 164700 7064
rect 164752 7052 164758 7064
rect 291286 7052 291292 7064
rect 164752 7024 291292 7052
rect 164752 7012 164758 7024
rect 291286 7012 291292 7024
rect 291344 7012 291350 7064
rect 168190 6944 168196 6996
rect 168248 6984 168254 6996
rect 292666 6984 292672 6996
rect 168248 6956 292672 6984
rect 168248 6944 168254 6956
rect 292666 6944 292672 6956
rect 292724 6944 292730 6996
rect 175366 6876 175372 6928
rect 175424 6916 175430 6928
rect 176562 6916 176568 6928
rect 175424 6888 176568 6916
rect 175424 6876 175430 6888
rect 176562 6876 176568 6888
rect 176620 6876 176626 6928
rect 193214 6876 193220 6928
rect 193272 6916 193278 6928
rect 194502 6916 194508 6928
rect 193272 6888 194508 6916
rect 193272 6876 193278 6888
rect 194502 6876 194508 6888
rect 194560 6876 194566 6928
rect 209866 6876 209872 6928
rect 209924 6916 209930 6928
rect 211062 6916 211068 6928
rect 209924 6888 211068 6916
rect 209924 6876 209930 6888
rect 211062 6876 211068 6888
rect 211120 6876 211126 6928
rect 227625 6919 227683 6925
rect 227625 6885 227637 6919
rect 227671 6916 227683 6919
rect 232038 6916 232044 6928
rect 227671 6888 232044 6916
rect 227671 6885 227683 6888
rect 227625 6879 227683 6885
rect 232038 6876 232044 6888
rect 232096 6876 232102 6928
rect 348050 6876 348056 6928
rect 348108 6916 348114 6928
rect 348234 6916 348240 6928
rect 348108 6888 348240 6916
rect 348108 6876 348114 6888
rect 348234 6876 348240 6888
rect 348292 6876 348298 6928
rect 174170 6808 174176 6860
rect 174228 6848 174234 6860
rect 295334 6848 295340 6860
rect 174228 6820 295340 6848
rect 174228 6808 174234 6820
rect 295334 6808 295340 6820
rect 295392 6808 295398 6860
rect 413922 6808 413928 6860
rect 413980 6848 413986 6860
rect 484578 6848 484584 6860
rect 413980 6820 484584 6848
rect 413980 6808 413986 6820
rect 484578 6808 484584 6820
rect 484636 6808 484642 6860
rect 170582 6740 170588 6792
rect 170640 6780 170646 6792
rect 293954 6780 293960 6792
rect 170640 6752 293960 6780
rect 170640 6740 170646 6752
rect 293954 6740 293960 6752
rect 294012 6740 294018 6792
rect 415302 6740 415308 6792
rect 415360 6780 415366 6792
rect 488166 6780 488172 6792
rect 415360 6752 488172 6780
rect 415360 6740 415366 6752
rect 488166 6740 488172 6752
rect 488224 6740 488230 6792
rect 167086 6672 167092 6724
rect 167144 6712 167150 6724
rect 292574 6712 292580 6724
rect 167144 6684 292580 6712
rect 167144 6672 167150 6684
rect 292574 6672 292580 6684
rect 292632 6672 292638 6724
rect 416590 6672 416596 6724
rect 416648 6712 416654 6724
rect 491754 6712 491760 6724
rect 416648 6684 491760 6712
rect 416648 6672 416654 6684
rect 491754 6672 491760 6684
rect 491812 6672 491818 6724
rect 163498 6604 163504 6656
rect 163556 6644 163562 6656
rect 291194 6644 291200 6656
rect 163556 6616 291200 6644
rect 163556 6604 163562 6616
rect 291194 6604 291200 6616
rect 291252 6604 291258 6656
rect 416682 6604 416688 6656
rect 416740 6644 416746 6656
rect 495342 6644 495348 6656
rect 416740 6616 495348 6644
rect 416740 6604 416746 6616
rect 495342 6604 495348 6616
rect 495400 6604 495406 6656
rect 131390 6536 131396 6588
rect 131448 6576 131454 6588
rect 279050 6576 279056 6588
rect 131448 6548 279056 6576
rect 131448 6536 131454 6548
rect 279050 6536 279056 6548
rect 279108 6536 279114 6588
rect 418062 6536 418068 6588
rect 418120 6576 418126 6588
rect 498930 6576 498936 6588
rect 418120 6548 498936 6576
rect 418120 6536 418126 6548
rect 498930 6536 498936 6548
rect 498988 6536 498994 6588
rect 76650 6468 76656 6520
rect 76708 6508 76714 6520
rect 258350 6508 258356 6520
rect 76708 6480 258356 6508
rect 76708 6468 76714 6480
rect 258350 6468 258356 6480
rect 258408 6468 258414 6520
rect 419442 6468 419448 6520
rect 419500 6508 419506 6520
rect 502426 6508 502432 6520
rect 419500 6480 502432 6508
rect 419500 6468 419506 6480
rect 502426 6468 502432 6480
rect 502484 6468 502490 6520
rect 73062 6400 73068 6452
rect 73120 6440 73126 6452
rect 256970 6440 256976 6452
rect 73120 6412 256976 6440
rect 73120 6400 73126 6412
rect 256970 6400 256976 6412
rect 257028 6400 257034 6452
rect 304994 6400 305000 6452
rect 305052 6440 305058 6452
rect 343726 6440 343732 6452
rect 305052 6412 343732 6440
rect 305052 6400 305058 6412
rect 343726 6400 343732 6412
rect 343784 6400 343790 6452
rect 420822 6400 420828 6452
rect 420880 6440 420886 6452
rect 506014 6440 506020 6452
rect 420880 6412 506020 6440
rect 420880 6400 420886 6412
rect 506014 6400 506020 6412
rect 506072 6400 506078 6452
rect 69474 6332 69480 6384
rect 69532 6372 69538 6384
rect 255406 6372 255412 6384
rect 69532 6344 255412 6372
rect 69532 6332 69538 6344
rect 255406 6332 255412 6344
rect 255464 6332 255470 6384
rect 284202 6332 284208 6384
rect 284260 6372 284266 6384
rect 334158 6372 334164 6384
rect 284260 6344 334164 6372
rect 284260 6332 284266 6344
rect 334158 6332 334164 6344
rect 334216 6332 334222 6384
rect 422202 6332 422208 6384
rect 422260 6372 422266 6384
rect 509602 6372 509608 6384
rect 422260 6344 509608 6372
rect 422260 6332 422266 6344
rect 509602 6332 509608 6344
rect 509660 6332 509666 6384
rect 65978 6264 65984 6316
rect 66036 6304 66042 6316
rect 254026 6304 254032 6316
rect 66036 6276 254032 6304
rect 66036 6264 66042 6276
rect 254026 6264 254032 6276
rect 254084 6264 254090 6316
rect 261018 6264 261024 6316
rect 261076 6304 261082 6316
rect 327166 6304 327172 6316
rect 261076 6276 327172 6304
rect 261076 6264 261082 6276
rect 327166 6264 327172 6276
rect 327224 6264 327230 6316
rect 423490 6264 423496 6316
rect 423548 6304 423554 6316
rect 513190 6304 513196 6316
rect 423548 6276 513196 6304
rect 423548 6264 423554 6276
rect 513190 6264 513196 6276
rect 513248 6264 513254 6316
rect 62390 6196 62396 6248
rect 62448 6236 62454 6248
rect 252738 6236 252744 6248
rect 62448 6208 252744 6236
rect 62448 6196 62454 6208
rect 252738 6196 252744 6208
rect 252796 6196 252802 6248
rect 257430 6196 257436 6248
rect 257488 6236 257494 6248
rect 325786 6236 325792 6248
rect 257488 6208 325792 6236
rect 257488 6196 257494 6208
rect 325786 6196 325792 6208
rect 325844 6196 325850 6248
rect 424870 6196 424876 6248
rect 424928 6236 424934 6248
rect 516778 6236 516784 6248
rect 424928 6208 516784 6236
rect 424928 6196 424934 6208
rect 516778 6196 516784 6208
rect 516836 6196 516842 6248
rect 58802 6128 58808 6180
rect 58860 6168 58866 6180
rect 251266 6168 251272 6180
rect 58860 6140 251272 6168
rect 58860 6128 58866 6140
rect 251266 6128 251272 6140
rect 251324 6128 251330 6180
rect 253842 6128 253848 6180
rect 253900 6168 253906 6180
rect 324406 6168 324412 6180
rect 253900 6140 324412 6168
rect 253900 6128 253906 6140
rect 324406 6128 324412 6140
rect 324464 6128 324470 6180
rect 426250 6128 426256 6180
rect 426308 6168 426314 6180
rect 520274 6168 520280 6180
rect 426308 6140 520280 6168
rect 426308 6128 426314 6140
rect 520274 6128 520280 6140
rect 520332 6128 520338 6180
rect 177758 6060 177764 6112
rect 177816 6100 177822 6112
rect 296714 6100 296720 6112
rect 177816 6072 296720 6100
rect 177816 6060 177822 6072
rect 296714 6060 296720 6072
rect 296772 6060 296778 6112
rect 411162 6060 411168 6112
rect 411220 6100 411226 6112
rect 479886 6100 479892 6112
rect 411220 6072 479892 6100
rect 411220 6060 411226 6072
rect 479886 6060 479892 6072
rect 479944 6060 479950 6112
rect 181346 5992 181352 6044
rect 181404 6032 181410 6044
rect 298094 6032 298100 6044
rect 181404 6004 298100 6032
rect 181404 5992 181410 6004
rect 298094 5992 298100 6004
rect 298152 5992 298158 6044
rect 409782 5992 409788 6044
rect 409840 6032 409846 6044
rect 476298 6032 476304 6044
rect 409840 6004 476304 6032
rect 409840 5992 409846 6004
rect 476298 5992 476304 6004
rect 476356 5992 476362 6044
rect 184842 5924 184848 5976
rect 184900 5964 184906 5976
rect 299474 5964 299480 5976
rect 184900 5936 299480 5964
rect 184900 5924 184906 5936
rect 299474 5924 299480 5936
rect 299532 5924 299538 5976
rect 408402 5924 408408 5976
rect 408460 5964 408466 5976
rect 472710 5964 472716 5976
rect 408460 5936 472716 5964
rect 408460 5924 408466 5936
rect 472710 5924 472716 5936
rect 472768 5924 472774 5976
rect 188430 5856 188436 5908
rect 188488 5896 188494 5908
rect 300854 5896 300860 5908
rect 188488 5868 300860 5896
rect 188488 5856 188494 5868
rect 300854 5856 300860 5868
rect 300912 5856 300918 5908
rect 407022 5856 407028 5908
rect 407080 5896 407086 5908
rect 469122 5896 469128 5908
rect 407080 5868 469128 5896
rect 407080 5856 407086 5868
rect 469122 5856 469128 5868
rect 469180 5856 469186 5908
rect 192018 5788 192024 5840
rect 192076 5828 192082 5840
rect 302234 5828 302240 5840
rect 192076 5800 302240 5828
rect 192076 5788 192082 5800
rect 302234 5788 302240 5800
rect 302292 5788 302298 5840
rect 405642 5788 405648 5840
rect 405700 5828 405706 5840
rect 465626 5828 465632 5840
rect 405700 5800 465632 5828
rect 405700 5788 405706 5800
rect 465626 5788 465632 5800
rect 465684 5788 465690 5840
rect 195606 5720 195612 5772
rect 195664 5760 195670 5772
rect 303614 5760 303620 5772
rect 195664 5732 303620 5760
rect 195664 5720 195670 5732
rect 303614 5720 303620 5732
rect 303672 5720 303678 5772
rect 404262 5720 404268 5772
rect 404320 5760 404326 5772
rect 462038 5760 462044 5772
rect 404320 5732 462044 5760
rect 404320 5720 404326 5732
rect 462038 5720 462044 5732
rect 462096 5720 462102 5772
rect 199194 5652 199200 5704
rect 199252 5692 199258 5704
rect 303706 5692 303712 5704
rect 199252 5664 303712 5692
rect 199252 5652 199258 5664
rect 303706 5652 303712 5664
rect 303764 5652 303770 5704
rect 402882 5652 402888 5704
rect 402940 5692 402946 5704
rect 458450 5692 458456 5704
rect 402940 5664 458456 5692
rect 402940 5652 402946 5664
rect 458450 5652 458456 5664
rect 458508 5652 458514 5704
rect 202690 5584 202696 5636
rect 202748 5624 202754 5636
rect 305178 5624 305184 5636
rect 202748 5596 305184 5624
rect 202748 5584 202754 5596
rect 305178 5584 305184 5596
rect 305236 5584 305242 5636
rect 401502 5584 401508 5636
rect 401560 5624 401566 5636
rect 454862 5624 454868 5636
rect 401560 5596 454868 5624
rect 401560 5584 401566 5596
rect 454862 5584 454868 5596
rect 454920 5584 454926 5636
rect 206278 5516 206284 5568
rect 206336 5556 206342 5568
rect 306466 5556 306472 5568
rect 206336 5528 306472 5556
rect 206336 5516 206342 5528
rect 306466 5516 306472 5528
rect 306524 5516 306530 5568
rect 137278 5448 137284 5500
rect 137336 5488 137342 5500
rect 281534 5488 281540 5500
rect 137336 5460 281540 5488
rect 137336 5448 137342 5460
rect 281534 5448 281540 5460
rect 281592 5448 281598 5500
rect 290734 5448 290740 5500
rect 290792 5488 290798 5500
rect 339586 5488 339592 5500
rect 290792 5460 339592 5488
rect 290792 5448 290798 5460
rect 339586 5448 339592 5460
rect 339644 5448 339650 5500
rect 390370 5448 390376 5500
rect 390428 5488 390434 5500
rect 423950 5488 423956 5500
rect 390428 5460 423956 5488
rect 390428 5448 390434 5460
rect 423950 5448 423956 5460
rect 424008 5448 424014 5500
rect 434622 5448 434628 5500
rect 434680 5488 434686 5500
rect 540514 5488 540520 5500
rect 434680 5460 540520 5488
rect 434680 5448 434686 5460
rect 540514 5448 540520 5460
rect 540572 5448 540578 5500
rect 133782 5380 133788 5432
rect 133840 5420 133846 5432
rect 280154 5420 280160 5432
rect 133840 5392 280160 5420
rect 133840 5380 133846 5392
rect 280154 5380 280160 5392
rect 280212 5380 280218 5432
rect 287146 5380 287152 5432
rect 287204 5420 287210 5432
rect 338206 5420 338212 5432
rect 287204 5392 338212 5420
rect 287204 5380 287210 5392
rect 338206 5380 338212 5392
rect 338264 5380 338270 5432
rect 391658 5380 391664 5432
rect 391716 5420 391722 5432
rect 426342 5420 426348 5432
rect 391716 5392 426348 5420
rect 391716 5380 391722 5392
rect 426342 5380 426348 5392
rect 426400 5380 426406 5432
rect 436002 5380 436008 5432
rect 436060 5420 436066 5432
rect 544102 5420 544108 5432
rect 436060 5392 544108 5420
rect 436060 5380 436066 5392
rect 544102 5380 544108 5392
rect 544160 5380 544166 5432
rect 130194 5312 130200 5364
rect 130252 5352 130258 5364
rect 278774 5352 278780 5364
rect 130252 5324 278780 5352
rect 130252 5312 130258 5324
rect 278774 5312 278780 5324
rect 278832 5312 278838 5364
rect 283650 5312 283656 5364
rect 283708 5352 283714 5364
rect 336826 5352 336832 5364
rect 283708 5324 336832 5352
rect 283708 5312 283714 5324
rect 336826 5312 336832 5324
rect 336884 5312 336890 5364
rect 393038 5312 393044 5364
rect 393096 5352 393102 5364
rect 429930 5352 429936 5364
rect 393096 5324 429936 5352
rect 393096 5312 393102 5324
rect 429930 5312 429936 5324
rect 429988 5312 429994 5364
rect 437382 5312 437388 5364
rect 437440 5352 437446 5364
rect 547690 5352 547696 5364
rect 437440 5324 547696 5352
rect 437440 5312 437446 5324
rect 547690 5312 547696 5324
rect 547748 5312 547754 5364
rect 67174 5244 67180 5296
rect 67232 5284 67238 5296
rect 254118 5284 254124 5296
rect 67232 5256 254124 5284
rect 67232 5244 67238 5256
rect 254118 5244 254124 5256
rect 254176 5244 254182 5296
rect 280062 5244 280068 5296
rect 280120 5284 280126 5296
rect 335538 5284 335544 5296
rect 280120 5256 335544 5284
rect 280120 5244 280126 5256
rect 335538 5244 335544 5256
rect 335596 5244 335602 5296
rect 394510 5244 394516 5296
rect 394568 5284 394574 5296
rect 433518 5284 433524 5296
rect 394568 5256 433524 5284
rect 394568 5244 394574 5256
rect 433518 5244 433524 5256
rect 433576 5244 433582 5296
rect 438762 5244 438768 5296
rect 438820 5284 438826 5296
rect 551186 5284 551192 5296
rect 438820 5256 551192 5284
rect 438820 5244 438826 5256
rect 551186 5244 551192 5256
rect 551244 5244 551250 5296
rect 51626 5176 51632 5228
rect 51684 5216 51690 5228
rect 248690 5216 248696 5228
rect 51684 5188 248696 5216
rect 51684 5176 51690 5188
rect 248690 5176 248696 5188
rect 248748 5176 248754 5228
rect 251450 5176 251456 5228
rect 251508 5216 251514 5228
rect 324314 5216 324320 5228
rect 251508 5188 324320 5216
rect 251508 5176 251514 5188
rect 324314 5176 324320 5188
rect 324372 5176 324378 5228
rect 394418 5176 394424 5228
rect 394476 5216 394482 5228
rect 434622 5216 434628 5228
rect 394476 5188 434628 5216
rect 394476 5176 394482 5188
rect 434622 5176 434628 5188
rect 434680 5176 434686 5228
rect 440050 5176 440056 5228
rect 440108 5216 440114 5228
rect 554774 5216 554780 5228
rect 440108 5188 554780 5216
rect 440108 5176 440114 5188
rect 554774 5176 554780 5188
rect 554832 5176 554838 5228
rect 48130 5108 48136 5160
rect 48188 5148 48194 5160
rect 247126 5148 247132 5160
rect 48188 5120 247132 5148
rect 48188 5108 48194 5120
rect 247126 5108 247132 5120
rect 247184 5108 247190 5160
rect 247954 5108 247960 5160
rect 248012 5148 248018 5160
rect 323302 5148 323308 5160
rect 248012 5120 323308 5148
rect 248012 5108 248018 5120
rect 323302 5108 323308 5120
rect 323360 5108 323366 5160
rect 395798 5108 395804 5160
rect 395856 5148 395862 5160
rect 437014 5148 437020 5160
rect 395856 5120 437020 5148
rect 395856 5108 395862 5120
rect 437014 5108 437020 5120
rect 437072 5108 437078 5160
rect 441522 5108 441528 5160
rect 441580 5148 441586 5160
rect 558362 5148 558368 5160
rect 441580 5120 558368 5148
rect 441580 5108 441586 5120
rect 558362 5108 558368 5120
rect 558420 5108 558426 5160
rect 12434 5040 12440 5092
rect 12492 5080 12498 5092
rect 233234 5080 233240 5092
rect 12492 5052 233240 5080
rect 12492 5040 12498 5052
rect 233234 5040 233240 5052
rect 233292 5040 233298 5092
rect 244366 5040 244372 5092
rect 244424 5080 244430 5092
rect 321830 5080 321836 5092
rect 244424 5052 321836 5080
rect 244424 5040 244430 5052
rect 321830 5040 321836 5052
rect 321888 5040 321894 5092
rect 395890 5040 395896 5092
rect 395948 5080 395954 5092
rect 438210 5080 438216 5092
rect 395948 5052 438216 5080
rect 395948 5040 395954 5052
rect 438210 5040 438216 5052
rect 438268 5040 438274 5092
rect 442810 5040 442816 5092
rect 442868 5080 442874 5092
rect 561950 5080 561956 5092
rect 442868 5052 561956 5080
rect 442868 5040 442874 5052
rect 561950 5040 561956 5052
rect 562008 5040 562014 5092
rect 7650 4972 7656 5024
rect 7708 5012 7714 5024
rect 231946 5012 231952 5024
rect 7708 4984 231952 5012
rect 7708 4972 7714 4984
rect 231946 4972 231952 4984
rect 232004 4972 232010 5024
rect 240778 4972 240784 5024
rect 240836 5012 240842 5024
rect 320450 5012 320456 5024
rect 240836 4984 320456 5012
rect 240836 4972 240842 4984
rect 320450 4972 320456 4984
rect 320508 4972 320514 5024
rect 397362 4972 397368 5024
rect 397420 5012 397426 5024
rect 440602 5012 440608 5024
rect 397420 4984 440608 5012
rect 397420 4972 397426 4984
rect 440602 4972 440608 4984
rect 440660 4972 440666 5024
rect 444282 4972 444288 5024
rect 444340 5012 444346 5024
rect 565538 5012 565544 5024
rect 444340 4984 565544 5012
rect 444340 4972 444346 4984
rect 565538 4972 565544 4984
rect 565596 4972 565602 5024
rect 2866 4904 2872 4956
rect 2924 4944 2930 4956
rect 224221 4947 224279 4953
rect 224221 4944 224233 4947
rect 2924 4916 224233 4944
rect 2924 4904 2930 4916
rect 224221 4913 224233 4916
rect 224267 4913 224279 4947
rect 224221 4907 224279 4913
rect 237190 4904 237196 4956
rect 237248 4944 237254 4956
rect 318702 4944 318708 4956
rect 237248 4916 318708 4944
rect 237248 4904 237254 4916
rect 318702 4904 318708 4916
rect 318760 4904 318766 4956
rect 318794 4904 318800 4956
rect 318852 4944 318858 4956
rect 346394 4944 346400 4956
rect 318852 4916 346400 4944
rect 318852 4904 318858 4916
rect 346394 4904 346400 4916
rect 346452 4904 346458 4956
rect 398650 4904 398656 4956
rect 398708 4944 398714 4956
rect 444190 4944 444196 4956
rect 398708 4916 444196 4944
rect 398708 4904 398714 4916
rect 444190 4904 444196 4916
rect 444248 4904 444254 4956
rect 445570 4904 445576 4956
rect 445628 4944 445634 4956
rect 569034 4944 569040 4956
rect 445628 4916 569040 4944
rect 445628 4904 445634 4916
rect 569034 4904 569040 4916
rect 569092 4904 569098 4956
rect 2777 4879 2835 4885
rect 2777 4845 2789 4879
rect 2823 4876 2835 4879
rect 12437 4879 12495 4885
rect 12437 4876 12449 4879
rect 2823 4848 12449 4876
rect 2823 4845 2835 4848
rect 2777 4839 2835 4845
rect 12437 4845 12449 4848
rect 12483 4845 12495 4879
rect 12437 4839 12495 4845
rect 19337 4879 19395 4885
rect 19337 4845 19349 4879
rect 19383 4876 19395 4879
rect 31757 4879 31815 4885
rect 31757 4876 31769 4879
rect 19383 4848 31769 4876
rect 19383 4845 19395 4848
rect 19337 4839 19395 4845
rect 31757 4845 31769 4848
rect 31803 4845 31815 4879
rect 31757 4839 31815 4845
rect 41417 4879 41475 4885
rect 41417 4845 41429 4879
rect 41463 4876 41475 4879
rect 51077 4879 51135 4885
rect 51077 4876 51089 4879
rect 41463 4848 51089 4876
rect 41463 4845 41475 4848
rect 41417 4839 41475 4845
rect 51077 4845 51089 4848
rect 51123 4845 51135 4879
rect 51077 4839 51135 4845
rect 60737 4879 60795 4885
rect 60737 4845 60749 4879
rect 60783 4876 60795 4879
rect 128357 4879 128415 4885
rect 128357 4876 128369 4879
rect 60783 4848 128369 4876
rect 60783 4845 60795 4848
rect 60737 4839 60795 4845
rect 128357 4845 128369 4848
rect 128403 4845 128415 4879
rect 128357 4839 128415 4845
rect 138017 4879 138075 4885
rect 138017 4845 138029 4879
rect 138063 4876 138075 4879
rect 147677 4879 147735 4885
rect 147677 4876 147689 4879
rect 138063 4848 147689 4876
rect 138063 4845 138075 4848
rect 138017 4839 138075 4845
rect 147677 4845 147689 4848
rect 147723 4845 147735 4879
rect 147677 4839 147735 4845
rect 157337 4879 157395 4885
rect 157337 4845 157349 4879
rect 157383 4876 157395 4879
rect 166997 4879 167055 4885
rect 166997 4876 167009 4879
rect 157383 4848 167009 4876
rect 157383 4845 157395 4848
rect 157337 4839 157395 4845
rect 166997 4845 167009 4848
rect 167043 4845 167055 4879
rect 166997 4839 167055 4845
rect 173897 4879 173955 4885
rect 173897 4845 173909 4879
rect 173943 4876 173955 4879
rect 186317 4879 186375 4885
rect 186317 4876 186329 4879
rect 173943 4848 186329 4876
rect 173943 4845 173955 4848
rect 173897 4839 173955 4845
rect 186317 4845 186329 4848
rect 186363 4845 186375 4879
rect 186317 4839 186375 4845
rect 195977 4879 196035 4885
rect 195977 4845 195989 4879
rect 196023 4876 196035 4879
rect 205637 4879 205695 4885
rect 205637 4876 205649 4879
rect 196023 4848 205649 4876
rect 196023 4845 196035 4848
rect 195977 4839 196035 4845
rect 205637 4845 205649 4848
rect 205683 4845 205695 4879
rect 205637 4839 205695 4845
rect 215205 4879 215263 4885
rect 215205 4845 215217 4879
rect 215251 4876 215263 4879
rect 229186 4876 229192 4888
rect 215251 4848 229192 4876
rect 215251 4845 215263 4848
rect 215205 4839 215263 4845
rect 229186 4836 229192 4848
rect 229244 4836 229250 4888
rect 230474 4876 230480 4888
rect 229388 4848 230480 4876
rect 566 4768 572 4820
rect 624 4808 630 4820
rect 224129 4811 224187 4817
rect 224129 4808 224141 4811
rect 624 4780 224141 4808
rect 624 4768 630 4780
rect 224129 4777 224141 4780
rect 224175 4777 224187 4811
rect 224129 4771 224187 4777
rect 224221 4811 224279 4817
rect 224221 4777 224233 4811
rect 224267 4808 224279 4811
rect 229388 4808 229416 4848
rect 230474 4836 230480 4848
rect 230532 4836 230538 4888
rect 233694 4836 233700 4888
rect 233752 4876 233758 4888
rect 317414 4876 317420 4888
rect 233752 4848 317420 4876
rect 233752 4836 233758 4848
rect 317414 4836 317420 4848
rect 317472 4836 317478 4888
rect 320174 4836 320180 4888
rect 320232 4876 320238 4888
rect 347866 4876 347872 4888
rect 320232 4848 347872 4876
rect 320232 4836 320238 4848
rect 347866 4836 347872 4848
rect 347924 4836 347930 4888
rect 397270 4836 397276 4888
rect 397328 4876 397334 4888
rect 441798 4876 441804 4888
rect 397328 4848 441804 4876
rect 397328 4836 397334 4848
rect 441798 4836 441804 4848
rect 441856 4836 441862 4888
rect 447042 4836 447048 4888
rect 447100 4876 447106 4888
rect 572622 4876 572628 4888
rect 447100 4848 572628 4876
rect 447100 4836 447106 4848
rect 572622 4836 572628 4848
rect 572680 4836 572686 4888
rect 224267 4780 229416 4808
rect 224267 4777 224279 4780
rect 224221 4771 224279 4777
rect 230106 4768 230112 4820
rect 230164 4808 230170 4820
rect 316034 4808 316040 4820
rect 230164 4780 316040 4808
rect 230164 4768 230170 4780
rect 316034 4768 316040 4780
rect 316092 4768 316098 4820
rect 316678 4768 316684 4820
rect 316736 4808 316742 4820
rect 345106 4808 345112 4820
rect 316736 4780 345112 4808
rect 316736 4768 316742 4780
rect 345106 4768 345112 4780
rect 345164 4768 345170 4820
rect 398742 4768 398748 4820
rect 398800 4808 398806 4820
rect 447778 4808 447784 4820
rect 398800 4780 447784 4808
rect 398800 4768 398806 4780
rect 447778 4768 447784 4780
rect 447836 4768 447842 4820
rect 448422 4768 448428 4820
rect 448480 4808 448486 4820
rect 576210 4808 576216 4820
rect 448480 4780 576216 4808
rect 448480 4768 448486 4780
rect 576210 4768 576216 4780
rect 576268 4768 576274 4820
rect 1670 4700 1676 4752
rect 1728 4740 1734 4752
rect 2777 4743 2835 4749
rect 2777 4740 2789 4743
rect 1728 4712 2789 4740
rect 1728 4700 1734 4712
rect 2777 4709 2789 4712
rect 2823 4709 2835 4743
rect 2777 4703 2835 4709
rect 12437 4743 12495 4749
rect 12437 4709 12449 4743
rect 12483 4740 12495 4743
rect 19337 4743 19395 4749
rect 19337 4740 19349 4743
rect 12483 4712 19349 4740
rect 12483 4709 12495 4712
rect 12437 4703 12495 4709
rect 19337 4709 19349 4712
rect 19383 4709 19395 4743
rect 19337 4703 19395 4709
rect 31757 4743 31815 4749
rect 31757 4709 31769 4743
rect 31803 4740 31815 4743
rect 41417 4743 41475 4749
rect 41417 4740 41429 4743
rect 31803 4712 41429 4740
rect 31803 4709 31815 4712
rect 31757 4703 31815 4709
rect 41417 4709 41429 4712
rect 41463 4709 41475 4743
rect 41417 4703 41475 4709
rect 51077 4743 51135 4749
rect 51077 4709 51089 4743
rect 51123 4740 51135 4743
rect 60737 4743 60795 4749
rect 60737 4740 60749 4743
rect 51123 4712 60749 4740
rect 51123 4709 51135 4712
rect 51077 4703 51135 4709
rect 60737 4709 60749 4712
rect 60783 4709 60795 4743
rect 60737 4703 60795 4709
rect 128357 4743 128415 4749
rect 128357 4709 128369 4743
rect 128403 4740 128415 4743
rect 138017 4743 138075 4749
rect 138017 4740 138029 4743
rect 128403 4712 138029 4740
rect 128403 4709 128415 4712
rect 128357 4703 128415 4709
rect 138017 4709 138029 4712
rect 138063 4709 138075 4743
rect 138017 4703 138075 4709
rect 147677 4743 147735 4749
rect 147677 4709 147689 4743
rect 147723 4740 147735 4743
rect 157337 4743 157395 4749
rect 157337 4740 157349 4743
rect 147723 4712 157349 4740
rect 147723 4709 147735 4712
rect 147677 4703 147735 4709
rect 157337 4709 157349 4712
rect 157383 4709 157395 4743
rect 157337 4703 157395 4709
rect 166997 4743 167055 4749
rect 166997 4709 167009 4743
rect 167043 4740 167055 4743
rect 173897 4743 173955 4749
rect 173897 4740 173909 4743
rect 167043 4712 173909 4740
rect 167043 4709 167055 4712
rect 166997 4703 167055 4709
rect 173897 4709 173909 4712
rect 173943 4709 173955 4743
rect 173897 4703 173955 4709
rect 186317 4743 186375 4749
rect 186317 4709 186329 4743
rect 186363 4740 186375 4743
rect 195977 4743 196035 4749
rect 195977 4740 195989 4743
rect 186363 4712 195989 4740
rect 186363 4709 186375 4712
rect 186317 4703 186375 4709
rect 195977 4709 195989 4712
rect 196023 4709 196035 4743
rect 195977 4703 196035 4709
rect 208670 4700 208676 4752
rect 208728 4740 208734 4752
rect 305089 4743 305147 4749
rect 208728 4712 305040 4740
rect 208728 4700 208734 4712
rect 212258 4632 212264 4684
rect 212316 4672 212322 4684
rect 305012 4672 305040 4712
rect 305089 4709 305101 4743
rect 305135 4740 305147 4743
rect 306837 4743 306895 4749
rect 306837 4740 306849 4743
rect 305135 4712 306849 4740
rect 305135 4709 305147 4712
rect 305089 4703 305147 4709
rect 306837 4709 306849 4712
rect 306883 4709 306895 4743
rect 306837 4703 306895 4709
rect 306929 4743 306987 4749
rect 306929 4709 306941 4743
rect 306975 4740 306987 4743
rect 314654 4740 314660 4752
rect 306975 4712 314660 4740
rect 306975 4709 306987 4712
rect 306929 4703 306987 4709
rect 314654 4700 314660 4712
rect 314712 4700 314718 4752
rect 315942 4700 315948 4752
rect 316000 4740 316006 4752
rect 331398 4740 331404 4752
rect 316000 4712 331404 4740
rect 316000 4700 316006 4712
rect 331398 4700 331404 4712
rect 331456 4700 331462 4752
rect 390462 4700 390468 4752
rect 390520 4740 390526 4752
rect 422754 4740 422760 4752
rect 390520 4712 422760 4740
rect 390520 4700 390526 4712
rect 422754 4700 422760 4712
rect 422812 4700 422818 4752
rect 433242 4700 433248 4752
rect 433300 4740 433306 4752
rect 536926 4740 536932 4752
rect 433300 4712 536932 4740
rect 433300 4700 433306 4712
rect 536926 4700 536932 4712
rect 536984 4700 536990 4752
rect 307754 4672 307760 4684
rect 212316 4644 304948 4672
rect 305012 4644 307760 4672
rect 212316 4632 212322 4644
rect 205637 4607 205695 4613
rect 205637 4573 205649 4607
rect 205683 4604 205695 4607
rect 215205 4607 215263 4613
rect 215205 4604 215217 4607
rect 205683 4576 215217 4604
rect 205683 4573 205695 4576
rect 205637 4567 205695 4573
rect 215205 4573 215217 4576
rect 215251 4573 215263 4607
rect 215205 4567 215263 4573
rect 215846 4564 215852 4616
rect 215904 4604 215910 4616
rect 304813 4607 304871 4613
rect 304813 4604 304825 4607
rect 215904 4576 304825 4604
rect 215904 4564 215910 4576
rect 304813 4573 304825 4576
rect 304859 4573 304871 4607
rect 304920 4604 304948 4644
rect 307754 4632 307760 4644
rect 307812 4632 307818 4684
rect 310514 4632 310520 4684
rect 310572 4672 310578 4684
rect 327074 4672 327080 4684
rect 310572 4644 327080 4672
rect 310572 4632 310578 4644
rect 327074 4632 327080 4644
rect 327132 4632 327138 4684
rect 387518 4632 387524 4684
rect 387576 4672 387582 4684
rect 415670 4672 415676 4684
rect 387576 4644 415676 4672
rect 387576 4632 387582 4644
rect 415670 4632 415676 4644
rect 415728 4632 415734 4684
rect 431862 4632 431868 4684
rect 431920 4672 431926 4684
rect 533430 4672 533436 4684
rect 431920 4644 533436 4672
rect 431920 4632 431926 4644
rect 533430 4632 533436 4644
rect 533488 4632 533494 4684
rect 309042 4604 309048 4616
rect 304920 4576 309048 4604
rect 304813 4567 304871 4573
rect 309042 4564 309048 4576
rect 309100 4564 309106 4616
rect 309134 4564 309140 4616
rect 309192 4604 309198 4616
rect 325694 4604 325700 4616
rect 309192 4576 325700 4604
rect 309192 4564 309198 4576
rect 325694 4564 325700 4576
rect 325752 4564 325758 4616
rect 386230 4564 386236 4616
rect 386288 4604 386294 4616
rect 413278 4604 413284 4616
rect 386288 4576 413284 4604
rect 386288 4564 386294 4576
rect 413278 4564 413284 4576
rect 413336 4564 413342 4616
rect 430482 4564 430488 4616
rect 430540 4604 430546 4616
rect 529842 4604 529848 4616
rect 430540 4576 529848 4604
rect 430540 4564 430546 4576
rect 529842 4564 529848 4576
rect 529900 4564 529906 4616
rect 219342 4496 219348 4548
rect 219400 4536 219406 4548
rect 311802 4536 311808 4548
rect 219400 4508 311808 4536
rect 219400 4496 219406 4508
rect 311802 4496 311808 4508
rect 311860 4496 311866 4548
rect 314562 4496 314568 4548
rect 314620 4536 314626 4548
rect 330018 4536 330024 4548
rect 314620 4508 330024 4536
rect 314620 4496 314626 4508
rect 330018 4496 330024 4508
rect 330076 4496 330082 4548
rect 429102 4496 429108 4548
rect 429160 4536 429166 4548
rect 526254 4536 526260 4548
rect 429160 4508 526260 4536
rect 429160 4496 429166 4508
rect 526254 4496 526260 4508
rect 526312 4496 526318 4548
rect 222930 4428 222936 4480
rect 222988 4468 222994 4480
rect 307113 4471 307171 4477
rect 222988 4440 307064 4468
rect 222988 4428 222994 4440
rect 226518 4360 226524 4412
rect 226576 4400 226582 4412
rect 306929 4403 306987 4409
rect 306929 4400 306941 4403
rect 226576 4372 306941 4400
rect 226576 4360 226582 4372
rect 306929 4369 306941 4372
rect 306975 4369 306987 4403
rect 307036 4400 307064 4440
rect 307113 4437 307125 4471
rect 307159 4468 307171 4471
rect 310606 4468 310612 4480
rect 307159 4440 310612 4468
rect 307159 4437 307171 4440
rect 307113 4431 307171 4437
rect 310606 4428 310612 4440
rect 310664 4428 310670 4480
rect 313182 4428 313188 4480
rect 313240 4468 313246 4480
rect 328638 4468 328644 4480
rect 313240 4440 328644 4468
rect 313240 4428 313246 4440
rect 328638 4428 328644 4440
rect 328696 4428 328702 4480
rect 427722 4428 427728 4480
rect 427780 4468 427786 4480
rect 522666 4468 522672 4480
rect 427780 4440 522672 4468
rect 427780 4428 427786 4440
rect 522666 4428 522672 4440
rect 522724 4428 522730 4480
rect 313274 4400 313280 4412
rect 307036 4372 313280 4400
rect 306929 4363 306987 4369
rect 313274 4360 313280 4372
rect 313332 4360 313338 4412
rect 317414 4360 317420 4412
rect 317472 4400 317478 4412
rect 332778 4400 332784 4412
rect 317472 4372 332784 4400
rect 317472 4360 317478 4372
rect 332778 4360 332784 4372
rect 332836 4360 332842 4412
rect 426250 4360 426256 4412
rect 426308 4400 426314 4412
rect 519078 4400 519084 4412
rect 426308 4372 519084 4400
rect 426308 4360 426314 4372
rect 519078 4360 519084 4372
rect 519136 4360 519142 4412
rect 201494 4292 201500 4344
rect 201552 4332 201558 4344
rect 267274 4332 267280 4344
rect 201552 4304 267280 4332
rect 201552 4292 201558 4304
rect 267274 4292 267280 4304
rect 267332 4292 267338 4344
rect 294322 4292 294328 4344
rect 294380 4332 294386 4344
rect 340966 4332 340972 4344
rect 294380 4304 340972 4332
rect 294380 4292 294386 4304
rect 340966 4292 340972 4304
rect 341024 4292 341030 4344
rect 424962 4292 424968 4344
rect 425020 4332 425026 4344
rect 515582 4332 515588 4344
rect 425020 4304 515588 4332
rect 425020 4292 425026 4304
rect 515582 4292 515588 4304
rect 515640 4292 515646 4344
rect 224129 4267 224187 4273
rect 224129 4233 224141 4267
rect 224175 4264 224187 4267
rect 229094 4264 229100 4276
rect 224175 4236 229100 4264
rect 224175 4233 224187 4236
rect 224129 4227 224187 4233
rect 229094 4224 229100 4236
rect 229152 4224 229158 4276
rect 298002 4224 298008 4276
rect 298060 4264 298066 4276
rect 341058 4264 341064 4276
rect 298060 4236 341064 4264
rect 298060 4224 298066 4236
rect 341058 4224 341064 4236
rect 341116 4224 341122 4276
rect 423582 4224 423588 4276
rect 423640 4264 423646 4276
rect 511994 4264 512000 4276
rect 423640 4236 512000 4264
rect 423640 4224 423646 4236
rect 511994 4224 512000 4236
rect 512052 4224 512058 4276
rect 124214 4156 124220 4208
rect 124272 4196 124278 4208
rect 125410 4196 125416 4208
rect 124272 4168 125416 4196
rect 124272 4156 124278 4168
rect 125410 4156 125416 4168
rect 125468 4156 125474 4208
rect 301406 4156 301412 4208
rect 301464 4196 301470 4208
rect 342438 4196 342444 4208
rect 301464 4168 342444 4196
rect 301464 4156 301470 4168
rect 342438 4156 342444 4168
rect 342496 4156 342502 4208
rect 344204 4168 345060 4196
rect 5258 4088 5264 4140
rect 5316 4128 5322 4140
rect 10318 4128 10324 4140
rect 5316 4100 10324 4128
rect 5316 4088 5322 4100
rect 10318 4088 10324 4100
rect 10376 4088 10382 4140
rect 36170 4088 36176 4140
rect 36228 4128 36234 4140
rect 39298 4128 39304 4140
rect 36228 4100 39304 4128
rect 36228 4088 36234 4100
rect 39298 4088 39304 4100
rect 39356 4088 39362 4140
rect 57606 4088 57612 4140
rect 57664 4128 57670 4140
rect 249058 4128 249064 4140
rect 57664 4100 249064 4128
rect 57664 4088 57670 4100
rect 249058 4088 249064 4100
rect 249116 4088 249122 4140
rect 268102 4088 268108 4140
rect 268160 4128 268166 4140
rect 269022 4128 269028 4140
rect 268160 4100 269028 4128
rect 268160 4088 268166 4100
rect 269022 4088 269028 4100
rect 269080 4088 269086 4140
rect 274082 4088 274088 4140
rect 274140 4128 274146 4140
rect 274542 4128 274548 4140
rect 274140 4100 274548 4128
rect 274140 4088 274146 4100
rect 274542 4088 274548 4100
rect 274600 4088 274606 4140
rect 275278 4088 275284 4140
rect 275336 4128 275342 4140
rect 276658 4128 276664 4140
rect 275336 4100 276664 4128
rect 275336 4088 275342 4100
rect 276658 4088 276664 4100
rect 276716 4088 276722 4140
rect 278866 4088 278872 4140
rect 278924 4128 278930 4140
rect 279970 4128 279976 4140
rect 278924 4100 279976 4128
rect 278924 4088 278930 4100
rect 279970 4088 279976 4100
rect 280028 4088 280034 4140
rect 281258 4088 281264 4140
rect 281316 4128 281322 4140
rect 284665 4131 284723 4137
rect 284665 4128 284677 4131
rect 281316 4100 284677 4128
rect 281316 4088 281322 4100
rect 284665 4097 284677 4100
rect 284711 4097 284723 4131
rect 284665 4091 284723 4097
rect 284754 4088 284760 4140
rect 284812 4128 284818 4140
rect 285582 4128 285588 4140
rect 284812 4100 285588 4128
rect 284812 4088 284818 4100
rect 285582 4088 285588 4100
rect 285640 4088 285646 4140
rect 291930 4088 291936 4140
rect 291988 4128 291994 4140
rect 292482 4128 292488 4140
rect 291988 4100 292488 4128
rect 291988 4088 291994 4100
rect 292482 4088 292488 4100
rect 292540 4088 292546 4140
rect 296714 4088 296720 4140
rect 296772 4128 296778 4140
rect 297910 4128 297916 4140
rect 296772 4100 297916 4128
rect 296772 4088 296778 4100
rect 297910 4088 297916 4100
rect 297968 4088 297974 4140
rect 307386 4088 307392 4140
rect 307444 4128 307450 4140
rect 344204 4128 344232 4168
rect 307444 4100 344232 4128
rect 307444 4088 307450 4100
rect 344278 4088 344284 4140
rect 344336 4128 344342 4140
rect 344922 4128 344928 4140
rect 344336 4100 344928 4128
rect 344336 4088 344342 4100
rect 344922 4088 344928 4100
rect 344980 4088 344986 4140
rect 345032 4128 345060 4168
rect 400122 4156 400128 4208
rect 400180 4196 400186 4208
rect 451274 4196 451280 4208
rect 400180 4168 451280 4196
rect 400180 4156 400186 4168
rect 451274 4156 451280 4168
rect 451332 4156 451338 4208
rect 477494 4156 477500 4208
rect 477552 4196 477558 4208
rect 478690 4196 478696 4208
rect 477552 4168 478696 4196
rect 477552 4156 477558 4168
rect 478690 4156 478696 4168
rect 478748 4156 478754 4208
rect 345198 4128 345204 4140
rect 345032 4100 345204 4128
rect 345198 4088 345204 4100
rect 345256 4088 345262 4140
rect 345474 4088 345480 4140
rect 345532 4128 345538 4140
rect 349798 4128 349804 4140
rect 345532 4100 349804 4128
rect 345532 4088 345538 4100
rect 349798 4088 349804 4100
rect 349856 4088 349862 4140
rect 349893 4131 349951 4137
rect 349893 4097 349905 4131
rect 349939 4128 349951 4131
rect 355318 4128 355324 4140
rect 349939 4100 355324 4128
rect 349939 4097 349951 4100
rect 349893 4091 349951 4097
rect 355318 4088 355324 4100
rect 355376 4088 355382 4140
rect 362126 4088 362132 4140
rect 362184 4128 362190 4140
rect 362862 4128 362868 4140
rect 362184 4100 362868 4128
rect 362184 4088 362190 4100
rect 362862 4088 362868 4100
rect 362920 4088 362926 4140
rect 364518 4088 364524 4140
rect 364576 4128 364582 4140
rect 366358 4128 366364 4140
rect 364576 4100 366364 4128
rect 364576 4088 364582 4100
rect 366358 4088 366364 4100
rect 366416 4088 366422 4140
rect 368014 4088 368020 4140
rect 368072 4128 368078 4140
rect 368474 4128 368480 4140
rect 368072 4100 368480 4128
rect 368072 4088 368078 4100
rect 368474 4088 368480 4100
rect 368532 4088 368538 4140
rect 368566 4088 368572 4140
rect 368624 4128 368630 4140
rect 369210 4128 369216 4140
rect 368624 4100 369216 4128
rect 368624 4088 368630 4100
rect 369210 4088 369216 4100
rect 369268 4088 369274 4140
rect 371142 4088 371148 4140
rect 371200 4128 371206 4140
rect 373994 4128 374000 4140
rect 371200 4100 374000 4128
rect 371200 4088 371206 4100
rect 373994 4088 374000 4100
rect 374052 4088 374058 4140
rect 381538 4088 381544 4140
rect 381596 4128 381602 4140
rect 384666 4128 384672 4140
rect 381596 4100 384672 4128
rect 381596 4088 381602 4100
rect 384666 4088 384672 4100
rect 384724 4088 384730 4140
rect 387702 4088 387708 4140
rect 387760 4128 387766 4140
rect 417970 4128 417976 4140
rect 387760 4100 417976 4128
rect 387760 4088 387766 4100
rect 417970 4088 417976 4100
rect 418028 4088 418034 4140
rect 421558 4088 421564 4140
rect 421616 4128 421622 4140
rect 503622 4128 503628 4140
rect 421616 4100 503628 4128
rect 421616 4088 421622 4100
rect 503622 4088 503628 4100
rect 503680 4088 503686 4140
rect 507118 4088 507124 4140
rect 507176 4128 507182 4140
rect 521470 4128 521476 4140
rect 507176 4100 521476 4128
rect 507176 4088 507182 4100
rect 521470 4088 521476 4100
rect 521528 4088 521534 4140
rect 525058 4088 525064 4140
rect 525116 4128 525122 4140
rect 560754 4128 560760 4140
rect 525116 4100 560760 4128
rect 525116 4088 525122 4100
rect 560754 4088 560760 4100
rect 560812 4088 560818 4140
rect 50522 4020 50528 4072
rect 50580 4060 50586 4072
rect 247678 4060 247684 4072
rect 50580 4032 247684 4060
rect 50580 4020 50586 4032
rect 247678 4020 247684 4032
rect 247736 4020 247742 4072
rect 269298 4020 269304 4072
rect 269356 4060 269362 4072
rect 315942 4060 315948 4072
rect 269356 4032 315948 4060
rect 269356 4020 269362 4032
rect 315942 4020 315948 4032
rect 316000 4020 316006 4072
rect 319254 4020 319260 4072
rect 319312 4060 319318 4072
rect 344370 4060 344376 4072
rect 319312 4032 344376 4060
rect 319312 4020 319318 4032
rect 344370 4020 344376 4032
rect 344428 4020 344434 4072
rect 346670 4020 346676 4072
rect 346728 4060 346734 4072
rect 356698 4060 356704 4072
rect 346728 4032 356704 4060
rect 346728 4020 346734 4032
rect 356698 4020 356704 4032
rect 356756 4020 356762 4072
rect 387610 4020 387616 4072
rect 387668 4060 387674 4072
rect 394053 4063 394111 4069
rect 387668 4032 394004 4060
rect 387668 4020 387674 4032
rect 46934 3952 46940 4004
rect 46992 3992 46998 4004
rect 247218 3992 247224 4004
rect 46992 3964 247224 3992
rect 46992 3952 46998 3964
rect 247218 3952 247224 3964
rect 247276 3952 247282 4004
rect 265802 3952 265808 4004
rect 265860 3992 265866 4004
rect 265860 3964 271920 3992
rect 265860 3952 265866 3964
rect 20714 3884 20720 3936
rect 20772 3924 20778 3936
rect 42058 3924 42064 3936
rect 20772 3896 42064 3924
rect 20772 3884 20778 3896
rect 42058 3884 42064 3896
rect 42116 3884 42122 3936
rect 45738 3884 45744 3936
rect 45796 3924 45802 3936
rect 246298 3924 246304 3936
rect 45796 3896 246304 3924
rect 45796 3884 45802 3896
rect 246298 3884 246304 3896
rect 246356 3884 246362 3936
rect 39758 3816 39764 3868
rect 39816 3856 39822 3868
rect 244274 3856 244280 3868
rect 39816 3828 244280 3856
rect 39816 3816 39822 3828
rect 244274 3816 244280 3828
rect 244332 3816 244338 3868
rect 270494 3816 270500 3868
rect 270552 3856 270558 3868
rect 271782 3856 271788 3868
rect 270552 3828 271788 3856
rect 270552 3816 270558 3828
rect 271782 3816 271788 3828
rect 271840 3816 271846 3868
rect 271892 3856 271920 3964
rect 272886 3952 272892 4004
rect 272944 3992 272950 4004
rect 317414 3992 317420 4004
rect 272944 3964 317420 3992
rect 272944 3952 272950 3964
rect 317414 3952 317420 3964
rect 317472 3952 317478 4004
rect 320450 3952 320456 4004
rect 320508 3992 320514 4004
rect 321462 3992 321468 4004
rect 320508 3964 321468 3992
rect 320508 3952 320514 3964
rect 321462 3952 321468 3964
rect 321520 3952 321526 4004
rect 321557 3995 321615 4001
rect 321557 3961 321569 3995
rect 321603 3992 321615 3995
rect 327810 3992 327816 4004
rect 321603 3964 327816 3992
rect 321603 3961 321615 3964
rect 321557 3955 321615 3961
rect 327810 3952 327816 3964
rect 327868 3952 327874 4004
rect 330018 3952 330024 4004
rect 330076 3992 330082 4004
rect 331122 3992 331128 4004
rect 330076 3964 331128 3992
rect 330076 3952 330082 3964
rect 331122 3952 331128 3964
rect 331180 3952 331186 4004
rect 335265 3995 335323 4001
rect 335265 3961 335277 3995
rect 335311 3992 335323 3995
rect 352006 3992 352012 4004
rect 335311 3964 352012 3992
rect 335311 3961 335323 3964
rect 335265 3955 335323 3961
rect 352006 3952 352012 3964
rect 352064 3952 352070 4004
rect 360930 3952 360936 4004
rect 360988 3992 360994 4004
rect 362218 3992 362224 4004
rect 360988 3964 362224 3992
rect 360988 3952 360994 3964
rect 362218 3952 362224 3964
rect 362276 3952 362282 4004
rect 389082 3952 389088 4004
rect 389140 3992 389146 4004
rect 393976 3992 394004 4032
rect 394053 4029 394065 4063
rect 394099 4060 394111 4063
rect 414474 4060 414480 4072
rect 394099 4032 414480 4060
rect 394099 4029 394111 4032
rect 394053 4023 394111 4029
rect 414474 4020 414480 4032
rect 414532 4020 414538 4072
rect 428458 4020 428464 4072
rect 428516 4060 428522 4072
rect 510798 4060 510804 4072
rect 428516 4032 510804 4060
rect 428516 4020 428522 4032
rect 510798 4020 510804 4032
rect 510856 4020 510862 4072
rect 527818 4020 527824 4072
rect 527876 4060 527882 4072
rect 567838 4060 567844 4072
rect 527876 4032 567844 4060
rect 527876 4020 527882 4032
rect 567838 4020 567844 4032
rect 567896 4020 567902 4072
rect 416866 3992 416872 4004
rect 389140 3964 393912 3992
rect 393976 3964 416872 3992
rect 389140 3952 389146 3964
rect 284665 3927 284723 3933
rect 284665 3893 284677 3927
rect 284711 3924 284723 3927
rect 290458 3924 290464 3936
rect 284711 3896 290464 3924
rect 284711 3893 284723 3896
rect 284665 3887 284723 3893
rect 290458 3884 290464 3896
rect 290516 3884 290522 3936
rect 293126 3884 293132 3936
rect 293184 3924 293190 3936
rect 339678 3924 339684 3936
rect 293184 3896 339684 3924
rect 293184 3884 293190 3896
rect 339678 3884 339684 3896
rect 339736 3884 339742 3936
rect 343082 3884 343088 3936
rect 343140 3924 343146 3936
rect 344557 3927 344615 3933
rect 343140 3896 344324 3924
rect 343140 3884 343146 3896
rect 314562 3856 314568 3868
rect 271892 3828 314568 3856
rect 314562 3816 314568 3828
rect 314620 3816 314626 3868
rect 316954 3816 316960 3868
rect 317012 3856 317018 3868
rect 344186 3856 344192 3868
rect 317012 3828 344192 3856
rect 317012 3816 317018 3828
rect 344186 3816 344192 3828
rect 344244 3816 344250 3868
rect 344296 3856 344324 3896
rect 344557 3893 344569 3927
rect 344603 3924 344615 3927
rect 352098 3924 352104 3936
rect 344603 3896 352104 3924
rect 344603 3893 344615 3896
rect 344557 3887 344615 3893
rect 352098 3884 352104 3896
rect 352156 3884 352162 3936
rect 384942 3884 384948 3936
rect 385000 3924 385006 3936
rect 388349 3927 388407 3933
rect 388349 3924 388361 3927
rect 385000 3896 388361 3924
rect 385000 3884 385006 3896
rect 388349 3893 388361 3896
rect 388395 3893 388407 3927
rect 388349 3887 388407 3893
rect 388990 3884 388996 3936
rect 389048 3924 389054 3936
rect 393685 3927 393743 3933
rect 393685 3924 393697 3927
rect 389048 3896 393697 3924
rect 389048 3884 389054 3896
rect 393685 3893 393697 3896
rect 393731 3893 393743 3927
rect 393685 3887 393743 3893
rect 349893 3859 349951 3865
rect 349893 3856 349905 3859
rect 344296 3828 349905 3856
rect 349893 3825 349905 3828
rect 349939 3825 349951 3859
rect 349893 3819 349951 3825
rect 376018 3816 376024 3868
rect 376076 3856 376082 3868
rect 383470 3856 383476 3868
rect 376076 3828 383476 3856
rect 376076 3816 376082 3828
rect 383470 3816 383476 3828
rect 383528 3816 383534 3868
rect 387058 3816 387064 3868
rect 387116 3856 387122 3868
rect 393038 3856 393044 3868
rect 387116 3828 393044 3856
rect 387116 3816 387122 3828
rect 393038 3816 393044 3828
rect 393096 3816 393102 3868
rect 393884 3856 393912 3964
rect 416866 3952 416872 3964
rect 416924 3952 416930 4004
rect 429838 3952 429844 4004
rect 429896 3992 429902 4004
rect 517882 3992 517888 4004
rect 429896 3964 517888 3992
rect 429896 3952 429902 3964
rect 517882 3952 517888 3964
rect 517940 3952 517946 4004
rect 529198 3952 529204 4004
rect 529256 3992 529262 4004
rect 575014 3992 575020 4004
rect 529256 3964 575020 3992
rect 529256 3952 529262 3964
rect 575014 3952 575020 3964
rect 575072 3952 575078 4004
rect 393961 3927 394019 3933
rect 393961 3893 393973 3927
rect 394007 3924 394019 3927
rect 420362 3924 420368 3936
rect 394007 3896 420368 3924
rect 394007 3893 394019 3896
rect 393961 3887 394019 3893
rect 420362 3884 420368 3896
rect 420420 3884 420426 3936
rect 434070 3884 434076 3936
rect 434128 3924 434134 3936
rect 525058 3924 525064 3936
rect 434128 3896 525064 3924
rect 434128 3884 434134 3896
rect 525058 3884 525064 3896
rect 525116 3884 525122 3936
rect 530578 3884 530584 3936
rect 530636 3924 530642 3936
rect 582190 3924 582196 3936
rect 530636 3896 582196 3924
rect 530636 3884 530642 3896
rect 582190 3884 582196 3896
rect 582248 3884 582254 3936
rect 421558 3856 421564 3868
rect 393884 3828 421564 3856
rect 421558 3816 421564 3828
rect 421616 3816 421622 3868
rect 436738 3816 436744 3868
rect 436796 3856 436802 3868
rect 532234 3856 532240 3868
rect 436796 3828 532240 3856
rect 436796 3816 436802 3828
rect 532234 3816 532240 3828
rect 532292 3816 532298 3868
rect 38562 3748 38568 3800
rect 38620 3788 38626 3800
rect 244458 3788 244464 3800
rect 38620 3760 244464 3788
rect 38620 3748 38626 3760
rect 244458 3748 244464 3760
rect 244516 3748 244522 3800
rect 262214 3748 262220 3800
rect 262272 3788 262278 3800
rect 313182 3788 313188 3800
rect 262272 3760 313188 3788
rect 262272 3748 262278 3760
rect 313182 3748 313188 3760
rect 313240 3748 313246 3800
rect 315758 3748 315764 3800
rect 315816 3788 315822 3800
rect 320174 3788 320180 3800
rect 315816 3760 320180 3788
rect 315816 3748 315822 3760
rect 320174 3748 320180 3760
rect 320232 3748 320238 3800
rect 325234 3748 325240 3800
rect 325292 3788 325298 3800
rect 330478 3788 330484 3800
rect 325292 3760 330484 3788
rect 325292 3748 325298 3760
rect 330478 3748 330484 3760
rect 330536 3748 330542 3800
rect 330573 3791 330631 3797
rect 330573 3757 330585 3791
rect 330619 3788 330631 3791
rect 350810 3788 350816 3800
rect 330619 3760 350816 3788
rect 330619 3757 330631 3760
rect 330573 3751 330631 3757
rect 350810 3748 350816 3760
rect 350868 3748 350874 3800
rect 374638 3748 374644 3800
rect 374696 3788 374702 3800
rect 381170 3788 381176 3800
rect 374696 3760 381176 3788
rect 374696 3748 374702 3760
rect 381170 3748 381176 3760
rect 381228 3748 381234 3800
rect 384850 3748 384856 3800
rect 384908 3788 384914 3800
rect 394329 3791 394387 3797
rect 394329 3788 394341 3791
rect 384908 3760 394341 3788
rect 384908 3748 384914 3760
rect 394329 3757 394341 3760
rect 394375 3757 394387 3791
rect 394329 3751 394387 3757
rect 394513 3791 394571 3797
rect 394513 3757 394525 3791
rect 394559 3788 394571 3791
rect 427538 3788 427544 3800
rect 394559 3760 427544 3788
rect 394559 3757 394571 3760
rect 394513 3751 394571 3757
rect 427538 3748 427544 3760
rect 427596 3748 427602 3800
rect 435174 3748 435180 3800
rect 435232 3788 435238 3800
rect 539318 3788 539324 3800
rect 435232 3760 539324 3788
rect 435232 3748 435238 3760
rect 539318 3748 539324 3760
rect 539376 3748 539382 3800
rect 32674 3680 32680 3732
rect 32732 3720 32738 3732
rect 241514 3720 241520 3732
rect 32732 3692 241520 3720
rect 32732 3680 32738 3692
rect 241514 3680 241520 3692
rect 241572 3680 241578 3732
rect 264606 3680 264612 3732
rect 264664 3720 264670 3732
rect 276382 3720 276388 3732
rect 264664 3692 276388 3720
rect 264664 3680 264670 3692
rect 276382 3680 276388 3692
rect 276440 3680 276446 3732
rect 276474 3680 276480 3732
rect 276532 3720 276538 3732
rect 284202 3720 284208 3732
rect 276532 3692 284208 3720
rect 276532 3680 276538 3692
rect 284202 3680 284208 3692
rect 284260 3680 284266 3732
rect 285950 3680 285956 3732
rect 286008 3720 286014 3732
rect 326433 3723 326491 3729
rect 326433 3720 326445 3723
rect 286008 3692 326445 3720
rect 286008 3680 286014 3692
rect 326433 3689 326445 3692
rect 326479 3689 326491 3723
rect 326433 3683 326491 3689
rect 328822 3680 328828 3732
rect 328880 3720 328886 3732
rect 334618 3720 334624 3732
rect 328880 3692 334624 3720
rect 328880 3680 328886 3692
rect 334618 3680 334624 3692
rect 334676 3680 334682 3732
rect 337102 3680 337108 3732
rect 337160 3720 337166 3732
rect 338022 3720 338028 3732
rect 337160 3692 338028 3720
rect 337160 3680 337166 3692
rect 338022 3680 338028 3692
rect 338080 3680 338086 3732
rect 339494 3680 339500 3732
rect 339552 3720 339558 3732
rect 357618 3720 357624 3732
rect 339552 3692 357624 3720
rect 339552 3680 339558 3692
rect 357618 3680 357624 3692
rect 357676 3680 357682 3732
rect 376662 3680 376668 3732
rect 376720 3720 376726 3732
rect 385862 3720 385868 3732
rect 376720 3692 385868 3720
rect 376720 3680 376726 3692
rect 385862 3680 385868 3692
rect 385920 3680 385926 3732
rect 386322 3680 386328 3732
rect 386380 3720 386386 3732
rect 386380 3692 387196 3720
rect 386380 3680 386386 3692
rect 25498 3612 25504 3664
rect 25556 3652 25562 3664
rect 238754 3652 238760 3664
rect 25556 3624 238760 3652
rect 25556 3612 25562 3624
rect 238754 3612 238760 3624
rect 238812 3612 238818 3664
rect 277670 3612 277676 3664
rect 277728 3652 277734 3664
rect 287698 3652 287704 3664
rect 277728 3624 287704 3652
rect 277728 3612 277734 3624
rect 287698 3612 287704 3624
rect 287756 3612 287762 3664
rect 288342 3612 288348 3664
rect 288400 3652 288406 3664
rect 338298 3652 338304 3664
rect 288400 3624 338304 3652
rect 288400 3612 288406 3624
rect 338298 3612 338304 3624
rect 338356 3612 338362 3664
rect 341886 3612 341892 3664
rect 341944 3652 341950 3664
rect 358814 3652 358820 3664
rect 341944 3624 358820 3652
rect 341944 3612 341950 3624
rect 358814 3612 358820 3624
rect 358872 3612 358878 3664
rect 377398 3612 377404 3664
rect 377456 3652 377462 3664
rect 387058 3652 387064 3664
rect 377456 3624 387064 3652
rect 377456 3612 377462 3624
rect 387058 3612 387064 3624
rect 387116 3612 387122 3664
rect 387168 3652 387196 3692
rect 393130 3680 393136 3732
rect 393188 3720 393194 3732
rect 394421 3723 394479 3729
rect 393188 3692 394188 3720
rect 393188 3680 393194 3692
rect 394053 3655 394111 3661
rect 394053 3652 394065 3655
rect 387168 3624 394065 3652
rect 394053 3621 394065 3624
rect 394099 3621 394111 3655
rect 394160 3652 394188 3692
rect 394421 3689 394433 3723
rect 394467 3720 394479 3723
rect 428734 3720 428740 3732
rect 394467 3692 428740 3720
rect 394467 3689 394479 3692
rect 394421 3683 394479 3689
rect 428734 3680 428740 3692
rect 428792 3680 428798 3732
rect 436830 3680 436836 3732
rect 436888 3720 436894 3732
rect 546494 3720 546500 3732
rect 436888 3692 546500 3720
rect 436888 3680 436894 3692
rect 546494 3680 546500 3692
rect 546552 3680 546558 3732
rect 431126 3652 431132 3664
rect 394160 3624 431132 3652
rect 394053 3615 394111 3621
rect 431126 3612 431132 3624
rect 431184 3612 431190 3664
rect 440142 3612 440148 3664
rect 440200 3652 440206 3664
rect 557166 3652 557172 3664
rect 440200 3624 557172 3652
rect 440200 3612 440206 3624
rect 557166 3612 557172 3624
rect 557224 3612 557230 3664
rect 11238 3544 11244 3596
rect 11296 3584 11302 3596
rect 19978 3584 19984 3596
rect 11296 3556 19984 3584
rect 11296 3544 11302 3556
rect 19978 3544 19984 3556
rect 20036 3544 20042 3596
rect 24302 3544 24308 3596
rect 24360 3584 24366 3596
rect 238846 3584 238852 3596
rect 24360 3556 238852 3584
rect 24360 3544 24366 3556
rect 238846 3544 238852 3556
rect 238904 3544 238910 3596
rect 258626 3544 258632 3596
rect 258684 3584 258690 3596
rect 310514 3584 310520 3596
rect 258684 3556 310520 3584
rect 258684 3544 258690 3556
rect 310514 3544 310520 3556
rect 310572 3544 310578 3596
rect 312170 3544 312176 3596
rect 312228 3584 312234 3596
rect 318794 3584 318800 3596
rect 312228 3556 318800 3584
rect 312228 3544 312234 3556
rect 318794 3544 318800 3556
rect 318852 3544 318858 3596
rect 324038 3544 324044 3596
rect 324096 3584 324102 3596
rect 344557 3587 344615 3593
rect 344557 3584 344569 3587
rect 324096 3556 344569 3584
rect 324096 3544 324102 3556
rect 344557 3553 344569 3556
rect 344603 3553 344615 3587
rect 344557 3547 344615 3553
rect 347866 3544 347872 3596
rect 347924 3584 347930 3596
rect 349062 3584 349068 3596
rect 347924 3556 349068 3584
rect 347924 3544 347930 3556
rect 349062 3544 349068 3556
rect 349120 3544 349126 3596
rect 353754 3544 353760 3596
rect 353812 3584 353818 3596
rect 358078 3584 358084 3596
rect 353812 3556 358084 3584
rect 353812 3544 353818 3556
rect 358078 3544 358084 3556
rect 358136 3544 358142 3596
rect 378042 3544 378048 3596
rect 378100 3584 378106 3596
rect 389450 3584 389456 3596
rect 378100 3556 389456 3584
rect 378100 3544 378106 3556
rect 389450 3544 389456 3556
rect 389508 3544 389514 3596
rect 391750 3544 391756 3596
rect 391808 3584 391814 3596
rect 391808 3556 391980 3584
rect 391808 3544 391814 3556
rect 16022 3476 16028 3528
rect 16080 3516 16086 3528
rect 235074 3516 235080 3528
rect 16080 3488 235080 3516
rect 16080 3476 16086 3488
rect 235074 3476 235080 3488
rect 235132 3476 235138 3528
rect 263597 3519 263655 3525
rect 263597 3485 263609 3519
rect 263643 3516 263655 3519
rect 290921 3519 290979 3525
rect 263643 3488 270540 3516
rect 263643 3485 263655 3488
rect 263597 3479 263655 3485
rect 14826 3408 14832 3460
rect 14884 3448 14890 3460
rect 234706 3448 234712 3460
rect 14884 3420 234712 3448
rect 14884 3408 14890 3420
rect 234706 3408 234712 3420
rect 234764 3408 234770 3460
rect 255038 3408 255044 3460
rect 255096 3448 255102 3460
rect 270512 3457 270540 3488
rect 290921 3485 290933 3519
rect 290967 3516 290979 3519
rect 326341 3519 326399 3525
rect 326341 3516 326353 3519
rect 290967 3488 326353 3516
rect 290967 3485 290979 3488
rect 290921 3479 290979 3485
rect 326341 3485 326353 3488
rect 326387 3485 326399 3519
rect 326341 3479 326399 3485
rect 326430 3476 326436 3528
rect 326488 3516 326494 3528
rect 330573 3519 330631 3525
rect 330573 3516 330585 3519
rect 326488 3488 330585 3516
rect 326488 3476 326494 3488
rect 330573 3485 330585 3488
rect 330619 3485 330631 3519
rect 334802 3516 334808 3528
rect 330573 3479 330631 3485
rect 331324 3488 334808 3516
rect 263505 3451 263563 3457
rect 263505 3448 263517 3451
rect 255096 3420 263517 3448
rect 255096 3408 255102 3420
rect 263505 3417 263517 3420
rect 263551 3417 263563 3451
rect 263505 3411 263563 3417
rect 270497 3451 270555 3457
rect 270497 3417 270509 3451
rect 270543 3417 270555 3451
rect 270497 3411 270555 3417
rect 270589 3451 270647 3457
rect 270589 3417 270601 3451
rect 270635 3448 270647 3451
rect 280065 3451 280123 3457
rect 280065 3448 280077 3451
rect 270635 3420 280077 3448
rect 270635 3417 270647 3420
rect 270589 3411 270647 3417
rect 280065 3417 280077 3420
rect 280111 3417 280123 3451
rect 280065 3411 280123 3417
rect 289725 3451 289783 3457
rect 289725 3417 289737 3451
rect 289771 3448 289783 3451
rect 292393 3451 292451 3457
rect 292393 3448 292405 3451
rect 289771 3420 292405 3448
rect 289771 3417 289783 3420
rect 289725 3411 289783 3417
rect 292393 3417 292405 3420
rect 292439 3417 292451 3451
rect 292393 3411 292451 3417
rect 292577 3451 292635 3457
rect 292577 3417 292589 3451
rect 292623 3448 292635 3451
rect 302237 3451 302295 3457
rect 302237 3448 302249 3451
rect 292623 3420 302249 3448
rect 292623 3417 292635 3420
rect 292577 3411 292635 3417
rect 302237 3417 302249 3420
rect 302283 3417 302295 3451
rect 302237 3411 302295 3417
rect 309244 3420 311940 3448
rect 19518 3340 19524 3392
rect 19576 3380 19582 3392
rect 28258 3380 28264 3392
rect 19576 3352 28264 3380
rect 19576 3340 19582 3352
rect 28258 3340 28264 3352
rect 28316 3340 28322 3392
rect 34974 3340 34980 3392
rect 35032 3380 35038 3392
rect 57238 3380 57244 3392
rect 35032 3352 57244 3380
rect 35032 3340 35038 3352
rect 57238 3340 57244 3352
rect 57296 3340 57302 3392
rect 64690 3340 64696 3392
rect 64748 3380 64754 3392
rect 250438 3380 250444 3392
rect 64748 3352 250444 3380
rect 64748 3340 64754 3352
rect 250438 3340 250444 3352
rect 250496 3340 250502 3392
rect 290921 3383 290979 3389
rect 290921 3380 290933 3383
rect 287808 3352 290933 3380
rect 10042 3272 10048 3324
rect 10100 3312 10106 3324
rect 13078 3312 13084 3324
rect 10100 3284 13084 3312
rect 10100 3272 10106 3284
rect 13078 3272 13084 3284
rect 13136 3272 13142 3324
rect 29086 3272 29092 3324
rect 29144 3312 29150 3324
rect 35158 3312 35164 3324
rect 29144 3284 35164 3312
rect 29144 3272 29150 3284
rect 35158 3272 35164 3284
rect 35216 3272 35222 3324
rect 42150 3272 42156 3324
rect 42208 3312 42214 3324
rect 66898 3312 66904 3324
rect 42208 3284 66904 3312
rect 42208 3272 42214 3284
rect 66898 3272 66904 3284
rect 66956 3272 66962 3324
rect 70670 3272 70676 3324
rect 70728 3312 70734 3324
rect 71682 3312 71688 3324
rect 70728 3284 71688 3312
rect 70728 3272 70734 3284
rect 71682 3272 71688 3284
rect 71740 3272 71746 3324
rect 71866 3272 71872 3324
rect 71924 3312 71930 3324
rect 251818 3312 251824 3324
rect 71924 3284 251824 3312
rect 71924 3272 71930 3284
rect 251818 3272 251824 3284
rect 251876 3272 251882 3324
rect 280157 3315 280215 3321
rect 280157 3312 280169 3315
rect 280080 3284 280169 3312
rect 43346 3204 43352 3256
rect 43404 3244 43410 3256
rect 61378 3244 61384 3256
rect 43404 3216 61384 3244
rect 43404 3204 43410 3216
rect 61378 3204 61384 3216
rect 61436 3204 61442 3256
rect 77846 3204 77852 3256
rect 77904 3244 77910 3256
rect 78582 3244 78588 3256
rect 77904 3216 78588 3244
rect 77904 3204 77910 3216
rect 78582 3204 78588 3216
rect 78640 3204 78646 3256
rect 81434 3204 81440 3256
rect 81492 3244 81498 3256
rect 82722 3244 82728 3256
rect 81492 3216 82728 3244
rect 81492 3204 81498 3216
rect 82722 3204 82728 3216
rect 82780 3204 82786 3256
rect 84838 3244 84844 3256
rect 82832 3216 84844 3244
rect 54018 3136 54024 3188
rect 54076 3176 54082 3188
rect 71038 3176 71044 3188
rect 54076 3148 71044 3176
rect 54076 3136 54082 3148
rect 71038 3136 71044 3148
rect 71096 3136 71102 3188
rect 75454 3136 75460 3188
rect 75512 3176 75518 3188
rect 79318 3176 79324 3188
rect 75512 3148 79324 3176
rect 75512 3136 75518 3148
rect 79318 3136 79324 3148
rect 79376 3136 79382 3188
rect 82630 3136 82636 3188
rect 82688 3176 82694 3188
rect 82832 3176 82860 3216
rect 84838 3204 84844 3216
rect 84896 3204 84902 3256
rect 84930 3204 84936 3256
rect 84988 3244 84994 3256
rect 85482 3244 85488 3256
rect 84988 3216 85488 3244
rect 84988 3204 84994 3216
rect 85482 3204 85488 3216
rect 85540 3204 85546 3256
rect 88518 3204 88524 3256
rect 88576 3244 88582 3256
rect 89622 3244 89628 3256
rect 88576 3216 89628 3244
rect 88576 3204 88582 3216
rect 89622 3204 89628 3216
rect 89680 3204 89686 3256
rect 253198 3244 253204 3256
rect 89732 3216 253204 3244
rect 82688 3148 82860 3176
rect 82909 3179 82967 3185
rect 82688 3136 82694 3148
rect 82909 3145 82921 3179
rect 82955 3176 82967 3179
rect 89732 3176 89760 3216
rect 253198 3204 253204 3216
rect 253256 3204 253262 3256
rect 280080 3253 280108 3284
rect 280157 3281 280169 3284
rect 280203 3281 280215 3315
rect 280157 3275 280215 3281
rect 280065 3247 280123 3253
rect 280065 3213 280077 3247
rect 280111 3213 280123 3247
rect 280065 3207 280123 3213
rect 254578 3176 254584 3188
rect 82955 3148 89760 3176
rect 93872 3148 254584 3176
rect 82955 3145 82967 3148
rect 82909 3139 82967 3145
rect 61194 3068 61200 3120
rect 61252 3108 61258 3120
rect 77938 3108 77944 3120
rect 61252 3080 77944 3108
rect 61252 3068 61258 3080
rect 77938 3068 77944 3080
rect 77996 3068 78002 3120
rect 89714 3068 89720 3120
rect 89772 3108 89778 3120
rect 93872 3108 93900 3148
rect 254578 3136 254584 3148
rect 254636 3136 254642 3188
rect 282454 3136 282460 3188
rect 282512 3176 282518 3188
rect 287808 3176 287836 3352
rect 290921 3349 290933 3352
rect 290967 3349 290979 3383
rect 290921 3343 290979 3349
rect 299106 3272 299112 3324
rect 299164 3312 299170 3324
rect 309244 3312 309272 3420
rect 311912 3380 311940 3420
rect 314562 3408 314568 3460
rect 314620 3448 314626 3460
rect 331217 3451 331275 3457
rect 331217 3448 331229 3451
rect 314620 3420 331229 3448
rect 314620 3408 314626 3420
rect 331217 3417 331229 3420
rect 331263 3417 331275 3451
rect 331217 3411 331275 3417
rect 321557 3383 321615 3389
rect 321557 3380 321569 3383
rect 311912 3352 321569 3380
rect 321557 3349 321569 3352
rect 321603 3349 321615 3383
rect 321557 3343 321615 3349
rect 321646 3340 321652 3392
rect 321704 3380 321710 3392
rect 326246 3380 326252 3392
rect 321704 3352 326252 3380
rect 321704 3340 321710 3352
rect 326246 3340 326252 3352
rect 326304 3340 326310 3392
rect 326341 3383 326399 3389
rect 326341 3349 326353 3383
rect 326387 3380 326399 3383
rect 331324 3380 331352 3488
rect 334802 3476 334808 3488
rect 334860 3476 334866 3528
rect 351362 3476 351368 3528
rect 351420 3516 351426 3528
rect 351822 3516 351828 3528
rect 351420 3488 351828 3516
rect 351420 3476 351426 3488
rect 351822 3476 351828 3488
rect 351880 3476 351886 3528
rect 352558 3476 352564 3528
rect 352616 3516 352622 3528
rect 353202 3516 353208 3528
rect 352616 3488 353208 3516
rect 352616 3476 352622 3488
rect 353202 3476 353208 3488
rect 353260 3476 353266 3528
rect 354950 3476 354956 3528
rect 355008 3516 355014 3528
rect 355962 3516 355968 3528
rect 355008 3488 355968 3516
rect 355008 3476 355014 3488
rect 355962 3476 355968 3488
rect 356020 3476 356026 3528
rect 361758 3516 361764 3528
rect 358188 3488 361764 3516
rect 331401 3451 331459 3457
rect 331401 3417 331413 3451
rect 331447 3448 331459 3451
rect 348050 3448 348056 3460
rect 331447 3420 348056 3448
rect 331447 3417 331459 3420
rect 331401 3411 331459 3417
rect 348050 3408 348056 3420
rect 348108 3408 348114 3460
rect 350258 3408 350264 3460
rect 350316 3448 350322 3460
rect 358188 3448 358216 3488
rect 361758 3476 361764 3488
rect 361816 3476 361822 3528
rect 363322 3476 363328 3528
rect 363380 3516 363386 3528
rect 364242 3516 364248 3528
rect 363380 3488 364248 3516
rect 363380 3476 363386 3488
rect 364242 3476 364248 3488
rect 364300 3476 364306 3528
rect 371050 3476 371056 3528
rect 371108 3516 371114 3528
rect 371602 3516 371608 3528
rect 371108 3488 371608 3516
rect 371108 3476 371114 3488
rect 371602 3476 371608 3488
rect 371660 3476 371666 3528
rect 373258 3476 373264 3528
rect 373316 3516 373322 3528
rect 377582 3516 377588 3528
rect 373316 3488 377588 3516
rect 373316 3476 373322 3488
rect 377582 3476 377588 3488
rect 377640 3476 377646 3528
rect 377950 3476 377956 3528
rect 378008 3516 378014 3528
rect 387153 3519 387211 3525
rect 387153 3516 387165 3519
rect 378008 3488 387165 3516
rect 378008 3476 378014 3488
rect 387153 3485 387165 3488
rect 387199 3485 387211 3519
rect 387153 3479 387211 3485
rect 388438 3476 388444 3528
rect 388496 3516 388502 3528
rect 391842 3516 391848 3528
rect 388496 3488 391848 3516
rect 388496 3476 388502 3488
rect 391842 3476 391848 3488
rect 391900 3476 391906 3528
rect 391952 3516 391980 3556
rect 393222 3544 393228 3596
rect 393280 3584 393286 3596
rect 432322 3584 432328 3596
rect 393280 3556 432328 3584
rect 393280 3544 393286 3556
rect 432322 3544 432328 3556
rect 432380 3544 432386 3596
rect 435450 3544 435456 3596
rect 435508 3584 435514 3596
rect 442261 3587 442319 3593
rect 442261 3584 442273 3587
rect 435508 3556 442273 3584
rect 435508 3544 435514 3556
rect 442261 3553 442273 3556
rect 442307 3553 442319 3587
rect 442261 3547 442319 3553
rect 442902 3544 442908 3596
rect 442960 3584 442966 3596
rect 564342 3584 564348 3596
rect 442960 3556 564348 3584
rect 442960 3544 442966 3556
rect 564342 3544 564348 3556
rect 564400 3544 564406 3596
rect 394421 3519 394479 3525
rect 394421 3516 394433 3519
rect 391952 3488 394433 3516
rect 394421 3485 394433 3488
rect 394467 3485 394479 3519
rect 394421 3479 394479 3485
rect 394602 3476 394608 3528
rect 394660 3516 394666 3528
rect 435818 3516 435824 3528
rect 394660 3488 435824 3516
rect 394660 3476 394666 3488
rect 435818 3476 435824 3488
rect 435876 3476 435882 3528
rect 438118 3476 438124 3528
rect 438176 3516 438182 3528
rect 446677 3519 446735 3525
rect 446677 3516 446689 3519
rect 438176 3488 446689 3516
rect 438176 3476 438182 3488
rect 446677 3485 446689 3488
rect 446723 3485 446735 3519
rect 446677 3479 446735 3485
rect 449158 3476 449164 3528
rect 449216 3516 449222 3528
rect 456153 3519 456211 3525
rect 449216 3488 456104 3516
rect 449216 3476 449222 3488
rect 350316 3420 358216 3448
rect 350316 3408 350322 3420
rect 373902 3408 373908 3460
rect 373960 3448 373966 3460
rect 378778 3448 378784 3460
rect 373960 3420 378784 3448
rect 373960 3408 373966 3420
rect 378778 3408 378784 3420
rect 378836 3408 378842 3460
rect 380158 3408 380164 3460
rect 380216 3448 380222 3460
rect 394234 3448 394240 3460
rect 380216 3420 394240 3448
rect 380216 3408 380222 3420
rect 394234 3408 394240 3420
rect 394292 3408 394298 3460
rect 394513 3451 394571 3457
rect 394513 3448 394525 3451
rect 394344 3420 394525 3448
rect 326387 3352 331352 3380
rect 326387 3349 326399 3352
rect 326341 3343 326399 3349
rect 332410 3340 332416 3392
rect 332468 3380 332474 3392
rect 354858 3380 354864 3392
rect 332468 3352 354864 3380
rect 332468 3340 332474 3352
rect 354858 3340 354864 3352
rect 354916 3340 354922 3392
rect 387153 3383 387211 3389
rect 387153 3349 387165 3383
rect 387199 3380 387211 3383
rect 390646 3380 390652 3392
rect 387199 3352 390652 3380
rect 387199 3349 387211 3352
rect 387153 3343 387211 3349
rect 390646 3340 390652 3352
rect 390704 3340 390710 3392
rect 391474 3340 391480 3392
rect 391532 3380 391538 3392
rect 394344 3380 394372 3420
rect 394513 3417 394525 3420
rect 394559 3417 394571 3451
rect 394513 3411 394571 3417
rect 395338 3408 395344 3460
rect 395396 3448 395402 3460
rect 400214 3448 400220 3460
rect 395396 3420 400220 3448
rect 395396 3408 395402 3420
rect 400214 3408 400220 3420
rect 400272 3408 400278 3460
rect 400309 3451 400367 3457
rect 400309 3417 400321 3451
rect 400355 3448 400367 3451
rect 439406 3448 439412 3460
rect 400355 3420 439412 3448
rect 400355 3417 400367 3420
rect 400309 3411 400367 3417
rect 439406 3408 439412 3420
rect 439464 3408 439470 3460
rect 442169 3451 442227 3457
rect 442169 3417 442181 3451
rect 442215 3448 442227 3451
rect 453666 3448 453672 3460
rect 442215 3420 453672 3448
rect 442215 3417 442227 3420
rect 442169 3411 442227 3417
rect 453666 3408 453672 3420
rect 453724 3408 453730 3460
rect 456076 3448 456104 3488
rect 456153 3485 456165 3519
rect 456199 3516 456211 3519
rect 571426 3516 571432 3528
rect 456199 3488 571432 3516
rect 456199 3485 456211 3488
rect 456153 3479 456211 3485
rect 571426 3476 571432 3488
rect 571484 3476 571490 3528
rect 578602 3448 578608 3460
rect 456076 3420 578608 3448
rect 578602 3408 578608 3420
rect 578660 3408 578666 3460
rect 391532 3352 394372 3380
rect 394421 3383 394479 3389
rect 391532 3340 391538 3352
rect 394421 3349 394433 3383
rect 394467 3380 394479 3383
rect 404909 3383 404967 3389
rect 404909 3380 404921 3383
rect 394467 3352 404921 3380
rect 394467 3349 394479 3352
rect 394421 3343 394479 3349
rect 404909 3349 404921 3352
rect 404955 3349 404967 3383
rect 404909 3343 404967 3349
rect 404998 3340 405004 3392
rect 405056 3380 405062 3392
rect 406102 3380 406108 3392
rect 405056 3352 406108 3380
rect 405056 3340 405062 3352
rect 406102 3340 406108 3352
rect 406160 3340 406166 3392
rect 422389 3383 422447 3389
rect 422389 3349 422401 3383
rect 422435 3380 422447 3383
rect 427173 3383 427231 3389
rect 427173 3380 427185 3383
rect 422435 3352 427185 3380
rect 422435 3349 422447 3352
rect 422389 3343 422447 3349
rect 427173 3349 427185 3352
rect 427219 3349 427231 3383
rect 427173 3343 427231 3349
rect 431218 3340 431224 3392
rect 431276 3380 431282 3392
rect 496538 3380 496544 3392
rect 431276 3352 496544 3380
rect 431276 3340 431282 3352
rect 496538 3340 496544 3352
rect 496596 3340 496602 3392
rect 500218 3340 500224 3392
rect 500276 3380 500282 3392
rect 507210 3380 507216 3392
rect 500276 3352 507216 3380
rect 500276 3340 500282 3352
rect 507210 3340 507216 3352
rect 507268 3340 507274 3392
rect 514386 3380 514392 3392
rect 507320 3352 514392 3380
rect 299164 3284 309272 3312
rect 299164 3272 299170 3284
rect 309778 3272 309784 3324
rect 309836 3312 309842 3324
rect 338758 3312 338764 3324
rect 309836 3284 338764 3312
rect 309836 3272 309842 3284
rect 338758 3272 338764 3284
rect 338816 3272 338822 3324
rect 349062 3272 349068 3324
rect 349120 3312 349126 3324
rect 351178 3312 351184 3324
rect 349120 3284 351184 3312
rect 349120 3272 349126 3284
rect 351178 3272 351184 3284
rect 351236 3272 351242 3324
rect 356146 3272 356152 3324
rect 356204 3312 356210 3324
rect 363230 3312 363236 3324
rect 356204 3284 363236 3312
rect 356204 3272 356210 3284
rect 363230 3272 363236 3284
rect 363288 3272 363294 3324
rect 365714 3272 365720 3324
rect 365772 3312 365778 3324
rect 366910 3312 366916 3324
rect 365772 3284 366916 3312
rect 365772 3272 365778 3284
rect 366910 3272 366916 3284
rect 366968 3272 366974 3324
rect 375282 3272 375288 3324
rect 375340 3312 375346 3324
rect 382366 3312 382372 3324
rect 375340 3284 382372 3312
rect 375340 3272 375346 3284
rect 382366 3272 382372 3284
rect 382424 3272 382430 3324
rect 383562 3272 383568 3324
rect 383620 3312 383626 3324
rect 407298 3312 407304 3324
rect 383620 3284 407304 3312
rect 383620 3272 383626 3284
rect 407298 3272 407304 3284
rect 407356 3272 407362 3324
rect 407758 3272 407764 3324
rect 407816 3312 407822 3324
rect 419166 3312 419172 3324
rect 407816 3284 419172 3312
rect 407816 3272 407822 3284
rect 419166 3272 419172 3284
rect 419224 3272 419230 3324
rect 420178 3272 420184 3324
rect 420236 3312 420242 3324
rect 475102 3312 475108 3324
rect 420236 3284 475108 3312
rect 420236 3272 420242 3284
rect 475102 3272 475108 3284
rect 475160 3272 475166 3324
rect 306190 3204 306196 3256
rect 306248 3244 306254 3256
rect 326341 3247 326399 3253
rect 326341 3244 326353 3247
rect 306248 3216 326353 3244
rect 306248 3204 306254 3216
rect 326341 3213 326353 3216
rect 326387 3213 326399 3247
rect 326341 3207 326399 3213
rect 326433 3247 326491 3253
rect 326433 3213 326445 3247
rect 326479 3244 326491 3247
rect 336918 3244 336924 3256
rect 326479 3216 336924 3244
rect 326479 3213 326491 3216
rect 326433 3207 326491 3213
rect 336918 3204 336924 3216
rect 336976 3204 336982 3256
rect 338298 3204 338304 3256
rect 338356 3244 338362 3256
rect 348418 3244 348424 3256
rect 338356 3216 348424 3244
rect 338356 3204 338362 3216
rect 348418 3204 348424 3216
rect 348476 3204 348482 3256
rect 384298 3204 384304 3256
rect 384356 3244 384362 3256
rect 388254 3244 388260 3256
rect 384356 3216 388260 3244
rect 384356 3204 384362 3216
rect 388254 3204 388260 3216
rect 388312 3204 388318 3256
rect 388349 3247 388407 3253
rect 388349 3213 388361 3247
rect 388395 3244 388407 3247
rect 408494 3244 408500 3256
rect 388395 3216 408500 3244
rect 388395 3213 388407 3216
rect 388349 3207 388407 3213
rect 408494 3204 408500 3216
rect 408552 3204 408558 3256
rect 409138 3204 409144 3256
rect 409196 3244 409202 3256
rect 412542 3244 412548 3256
rect 409196 3216 412548 3244
rect 409196 3204 409202 3216
rect 412542 3204 412548 3216
rect 412600 3204 412606 3256
rect 422297 3247 422355 3253
rect 422297 3213 422309 3247
rect 422343 3244 422355 3247
rect 427081 3247 427139 3253
rect 427081 3244 427093 3247
rect 422343 3216 427093 3244
rect 422343 3213 422355 3216
rect 422297 3207 422355 3213
rect 427081 3213 427093 3216
rect 427127 3213 427139 3247
rect 427081 3207 427139 3213
rect 427173 3247 427231 3253
rect 427173 3213 427185 3247
rect 427219 3244 427231 3247
rect 432509 3247 432567 3253
rect 432509 3244 432521 3247
rect 427219 3216 432521 3244
rect 427219 3213 427231 3216
rect 427173 3207 427231 3213
rect 432509 3213 432521 3216
rect 432555 3213 432567 3247
rect 432509 3207 432567 3213
rect 432601 3247 432659 3253
rect 432601 3213 432613 3247
rect 432647 3244 432659 3247
rect 441985 3247 442043 3253
rect 441985 3244 441997 3247
rect 432647 3216 441997 3244
rect 432647 3213 432659 3216
rect 432601 3207 432659 3213
rect 441985 3213 441997 3216
rect 442031 3213 442043 3247
rect 441985 3207 442043 3213
rect 442261 3247 442319 3253
rect 442261 3213 442273 3247
rect 442307 3244 442319 3247
rect 489362 3244 489368 3256
rect 442307 3216 489368 3244
rect 442307 3213 442319 3216
rect 442261 3207 442319 3213
rect 489362 3204 489368 3216
rect 489420 3204 489426 3256
rect 502978 3204 502984 3256
rect 503036 3244 503042 3256
rect 507320 3244 507348 3352
rect 514386 3340 514392 3352
rect 514444 3340 514450 3392
rect 523678 3340 523684 3392
rect 523736 3380 523742 3392
rect 553578 3380 553584 3392
rect 523736 3352 553584 3380
rect 523736 3340 523742 3352
rect 553578 3340 553584 3352
rect 553636 3340 553642 3392
rect 520918 3272 520924 3324
rect 520976 3312 520982 3324
rect 550082 3312 550088 3324
rect 520976 3284 550088 3312
rect 520976 3272 520982 3284
rect 550082 3272 550088 3284
rect 550140 3272 550146 3324
rect 503036 3216 507348 3244
rect 503036 3204 503042 3216
rect 518158 3204 518164 3256
rect 518216 3244 518222 3256
rect 542906 3244 542912 3256
rect 518216 3216 542912 3244
rect 518216 3204 518222 3216
rect 542906 3204 542912 3216
rect 542964 3204 542970 3256
rect 282512 3148 287836 3176
rect 282512 3136 282518 3148
rect 289538 3136 289544 3188
rect 289596 3176 289602 3188
rect 316586 3176 316592 3188
rect 289596 3148 316592 3176
rect 289596 3136 289602 3148
rect 316586 3136 316592 3148
rect 316644 3136 316650 3188
rect 327626 3136 327632 3188
rect 327684 3176 327690 3188
rect 352466 3176 352472 3188
rect 327684 3148 352472 3176
rect 327684 3136 327690 3148
rect 352466 3136 352472 3148
rect 352524 3136 352530 3188
rect 382090 3136 382096 3188
rect 382148 3176 382154 3188
rect 403710 3176 403716 3188
rect 382148 3148 403716 3176
rect 382148 3136 382154 3148
rect 403710 3136 403716 3148
rect 403768 3136 403774 3188
rect 404909 3179 404967 3185
rect 404909 3145 404921 3179
rect 404955 3176 404967 3179
rect 409690 3176 409696 3188
rect 404955 3148 409696 3176
rect 404955 3145 404967 3148
rect 404909 3139 404967 3145
rect 409690 3136 409696 3148
rect 409748 3136 409754 3188
rect 411898 3136 411904 3188
rect 411956 3176 411962 3188
rect 411956 3148 412220 3176
rect 411956 3136 411962 3148
rect 89772 3080 93900 3108
rect 89772 3068 89778 3080
rect 94498 3068 94504 3120
rect 94556 3108 94562 3120
rect 95142 3108 95148 3120
rect 94556 3080 95148 3108
rect 94556 3068 94562 3080
rect 95142 3068 95148 3080
rect 95200 3068 95206 3120
rect 95694 3068 95700 3120
rect 95752 3108 95758 3120
rect 96522 3108 96528 3120
rect 95752 3080 96528 3108
rect 95752 3068 95758 3080
rect 96522 3068 96528 3080
rect 96580 3068 96586 3120
rect 98086 3068 98092 3120
rect 98144 3108 98150 3120
rect 99190 3108 99196 3120
rect 98144 3080 99196 3108
rect 98144 3068 98150 3080
rect 99190 3068 99196 3080
rect 99248 3068 99254 3120
rect 101582 3068 101588 3120
rect 101640 3108 101646 3120
rect 102042 3108 102048 3120
rect 101640 3080 102048 3108
rect 101640 3068 101646 3080
rect 102042 3068 102048 3080
rect 102100 3068 102106 3120
rect 102778 3068 102784 3120
rect 102836 3108 102842 3120
rect 103422 3108 103428 3120
rect 102836 3080 103428 3108
rect 102836 3068 102842 3080
rect 103422 3068 103428 3080
rect 103480 3068 103486 3120
rect 105170 3068 105176 3120
rect 105228 3108 105234 3120
rect 106182 3108 106188 3120
rect 105228 3080 106188 3108
rect 105228 3068 105234 3080
rect 106182 3068 106188 3080
rect 106240 3068 106246 3120
rect 106366 3068 106372 3120
rect 106424 3108 106430 3120
rect 107470 3108 107476 3120
rect 106424 3080 107476 3108
rect 106424 3068 106430 3080
rect 107470 3068 107476 3080
rect 107528 3068 107534 3120
rect 254670 3108 254676 3120
rect 108316 3080 254676 3108
rect 68278 3000 68284 3052
rect 68336 3040 68342 3052
rect 102594 3040 102600 3052
rect 68336 3012 102600 3040
rect 68336 3000 68342 3012
rect 102594 3000 102600 3012
rect 102652 3000 102658 3052
rect 79042 2932 79048 2984
rect 79100 2972 79106 2984
rect 82909 2975 82967 2981
rect 82909 2972 82921 2975
rect 79100 2944 82921 2972
rect 79100 2932 79106 2944
rect 82909 2941 82921 2944
rect 82955 2941 82967 2975
rect 82909 2935 82967 2941
rect 86126 2932 86132 2984
rect 86184 2972 86190 2984
rect 102781 2975 102839 2981
rect 86184 2944 97488 2972
rect 86184 2932 86190 2944
rect 93302 2864 93308 2916
rect 93360 2904 93366 2916
rect 97258 2904 97264 2916
rect 93360 2876 97264 2904
rect 93360 2864 93366 2876
rect 97258 2864 97264 2876
rect 97316 2864 97322 2916
rect 96890 2796 96896 2848
rect 96948 2836 96954 2848
rect 97460 2836 97488 2944
rect 102781 2941 102793 2975
rect 102827 2972 102839 2975
rect 108316 2972 108344 3080
rect 254670 3068 254676 3080
rect 254728 3068 254734 3120
rect 280157 3111 280215 3117
rect 280157 3077 280169 3111
rect 280203 3108 280215 3111
rect 289725 3111 289783 3117
rect 289725 3108 289737 3111
rect 280203 3080 289737 3108
rect 280203 3077 280215 3080
rect 280157 3071 280215 3077
rect 289725 3077 289737 3080
rect 289771 3077 289783 3111
rect 289725 3071 289783 3077
rect 295518 3068 295524 3120
rect 295576 3108 295582 3120
rect 312538 3108 312544 3120
rect 295576 3080 312544 3108
rect 295576 3068 295582 3080
rect 312538 3068 312544 3080
rect 312596 3068 312602 3120
rect 319438 3108 319444 3120
rect 313292 3080 319444 3108
rect 255958 3040 255964 3052
rect 102827 2944 108344 2972
rect 108408 3012 255964 3040
rect 102827 2941 102839 2944
rect 102781 2935 102839 2941
rect 103974 2864 103980 2916
rect 104032 2904 104038 2916
rect 108408 2904 108436 3012
rect 255958 3000 255964 3012
rect 256016 3000 256022 3052
rect 300302 3000 300308 3052
rect 300360 3040 300366 3052
rect 313292 3040 313320 3080
rect 319438 3068 319444 3080
rect 319496 3068 319502 3120
rect 341518 3108 341524 3120
rect 326448 3080 341524 3108
rect 300360 3012 313320 3040
rect 300360 3000 300366 3012
rect 313366 3000 313372 3052
rect 313424 3040 313430 3052
rect 326448 3040 326476 3080
rect 341518 3068 341524 3080
rect 341576 3068 341582 3120
rect 357342 3068 357348 3120
rect 357400 3108 357406 3120
rect 359458 3108 359464 3120
rect 357400 3080 359464 3108
rect 357400 3068 357406 3080
rect 359458 3068 359464 3080
rect 359516 3068 359522 3120
rect 382182 3068 382188 3120
rect 382240 3108 382246 3120
rect 401318 3108 401324 3120
rect 382240 3080 401324 3108
rect 382240 3068 382246 3080
rect 401318 3068 401324 3080
rect 401376 3068 401382 3120
rect 405090 3068 405096 3120
rect 405148 3108 405154 3120
rect 412082 3108 412088 3120
rect 405148 3080 412088 3108
rect 405148 3068 405154 3080
rect 412082 3068 412088 3080
rect 412140 3068 412146 3120
rect 412192 3108 412220 3148
rect 417418 3136 417424 3188
rect 417476 3176 417482 3188
rect 467926 3176 467932 3188
rect 417476 3148 467932 3176
rect 417476 3136 417482 3148
rect 467926 3136 467932 3148
rect 467984 3136 467990 3188
rect 496078 3136 496084 3188
rect 496136 3176 496142 3188
rect 500126 3176 500132 3188
rect 496136 3148 500132 3176
rect 496136 3136 496142 3148
rect 500126 3136 500132 3148
rect 500184 3136 500190 3188
rect 514018 3136 514024 3188
rect 514076 3176 514082 3188
rect 535730 3176 535736 3188
rect 514076 3148 535736 3176
rect 514076 3136 514082 3148
rect 535730 3136 535736 3148
rect 535788 3136 535794 3188
rect 460842 3108 460848 3120
rect 412192 3080 460848 3108
rect 460842 3068 460848 3080
rect 460900 3068 460906 3120
rect 511258 3068 511264 3120
rect 511316 3108 511322 3120
rect 528646 3108 528652 3120
rect 511316 3080 528652 3108
rect 511316 3068 511322 3080
rect 528646 3068 528652 3080
rect 528704 3068 528710 3120
rect 313424 3012 326476 3040
rect 326525 3043 326583 3049
rect 313424 3000 313430 3012
rect 326525 3009 326537 3043
rect 326571 3040 326583 3043
rect 345750 3040 345756 3052
rect 326571 3012 345756 3040
rect 326571 3009 326583 3012
rect 326525 3003 326583 3009
rect 345750 3000 345756 3012
rect 345808 3000 345814 3052
rect 380802 3000 380808 3052
rect 380860 3040 380866 3052
rect 397822 3040 397828 3052
rect 380860 3012 397828 3040
rect 380860 3000 380866 3012
rect 397822 3000 397828 3012
rect 397880 3000 397886 3052
rect 402606 3000 402612 3052
rect 402664 3040 402670 3052
rect 425146 3040 425152 3052
rect 402664 3012 425152 3040
rect 402664 3000 402670 3012
rect 425146 3000 425152 3012
rect 425204 3000 425210 3052
rect 427081 3043 427139 3049
rect 427081 3009 427093 3043
rect 427127 3040 427139 3043
rect 432601 3043 432659 3049
rect 432601 3040 432613 3043
rect 427127 3012 432613 3040
rect 427127 3009 427139 3012
rect 427081 3003 427139 3009
rect 432601 3009 432613 3012
rect 432647 3009 432659 3043
rect 432601 3003 432659 3009
rect 433978 3000 433984 3052
rect 434036 3040 434042 3052
rect 481082 3040 481088 3052
rect 434036 3012 481088 3040
rect 434036 3000 434042 3012
rect 481082 3000 481088 3012
rect 481140 3000 481146 3052
rect 112346 2932 112352 2984
rect 112404 2972 112410 2984
rect 113082 2972 113088 2984
rect 112404 2944 113088 2972
rect 112404 2932 112410 2944
rect 113082 2932 113088 2944
rect 113140 2932 113146 2984
rect 113542 2932 113548 2984
rect 113600 2972 113606 2984
rect 114462 2972 114468 2984
rect 113600 2944 114468 2972
rect 113600 2932 113606 2944
rect 114462 2932 114468 2944
rect 114520 2932 114526 2984
rect 115934 2932 115940 2984
rect 115992 2972 115998 2984
rect 116946 2972 116952 2984
rect 115992 2944 116952 2972
rect 115992 2932 115998 2944
rect 116946 2932 116952 2944
rect 117004 2932 117010 2984
rect 119430 2932 119436 2984
rect 119488 2972 119494 2984
rect 119982 2972 119988 2984
rect 119488 2944 119988 2972
rect 119488 2932 119494 2944
rect 119982 2932 119988 2944
rect 120040 2932 120046 2984
rect 120626 2932 120632 2984
rect 120684 2972 120690 2984
rect 121362 2972 121368 2984
rect 120684 2944 121368 2972
rect 120684 2932 120690 2944
rect 121362 2932 121368 2944
rect 121420 2932 121426 2984
rect 257338 2972 257344 2984
rect 121472 2944 257344 2972
rect 104032 2876 108436 2904
rect 104032 2864 104038 2876
rect 111150 2864 111156 2916
rect 111208 2904 111214 2916
rect 121472 2904 121500 2944
rect 257338 2932 257344 2944
rect 257396 2932 257402 2984
rect 271690 2932 271696 2984
rect 271748 2972 271754 2984
rect 273898 2972 273904 2984
rect 271748 2944 273904 2972
rect 271748 2932 271754 2944
rect 273898 2932 273904 2944
rect 273956 2932 273962 2984
rect 302237 2975 302295 2981
rect 302237 2941 302249 2975
rect 302283 2972 302295 2975
rect 302283 2944 303660 2972
rect 302283 2941 302295 2944
rect 302237 2935 302295 2941
rect 258718 2904 258724 2916
rect 111208 2876 121500 2904
rect 121564 2876 258724 2904
rect 111208 2864 111214 2876
rect 105538 2836 105544 2848
rect 96948 2808 97396 2836
rect 97460 2808 105544 2836
rect 96948 2796 96954 2808
rect 97368 2768 97396 2808
rect 105538 2796 105544 2808
rect 105596 2796 105602 2848
rect 114738 2796 114744 2848
rect 114796 2836 114802 2848
rect 121564 2836 121592 2876
rect 258718 2864 258724 2876
rect 258776 2864 258782 2916
rect 302602 2864 302608 2916
rect 302660 2904 302666 2916
rect 303522 2904 303528 2916
rect 302660 2876 303528 2904
rect 302660 2864 302666 2876
rect 303522 2864 303528 2876
rect 303580 2864 303586 2916
rect 303632 2904 303660 2944
rect 303798 2932 303804 2984
rect 303856 2972 303862 2984
rect 322198 2972 322204 2984
rect 303856 2944 322204 2972
rect 303856 2932 303862 2944
rect 322198 2932 322204 2944
rect 322256 2932 322262 2984
rect 326154 2972 326160 2984
rect 322768 2944 326160 2972
rect 309134 2904 309140 2916
rect 303632 2876 309140 2904
rect 309134 2864 309140 2876
rect 309192 2864 309198 2916
rect 310974 2864 310980 2916
rect 311032 2904 311038 2916
rect 322768 2904 322796 2944
rect 326154 2932 326160 2944
rect 326212 2932 326218 2984
rect 326341 2975 326399 2981
rect 326341 2941 326353 2975
rect 326387 2972 326399 2975
rect 334618 2972 334624 2984
rect 326387 2944 334624 2972
rect 326387 2941 326399 2944
rect 326341 2935 326399 2941
rect 334618 2932 334624 2944
rect 334676 2932 334682 2984
rect 334710 2932 334716 2984
rect 334768 2972 334774 2984
rect 356422 2972 356428 2984
rect 334768 2944 356428 2972
rect 334768 2932 334774 2944
rect 356422 2932 356428 2944
rect 356480 2932 356486 2984
rect 381630 2932 381636 2984
rect 381688 2972 381694 2984
rect 395430 2972 395436 2984
rect 381688 2944 395436 2972
rect 381688 2932 381694 2944
rect 395430 2932 395436 2944
rect 395488 2932 395494 2984
rect 395982 2932 395988 2984
rect 396040 2972 396046 2984
rect 400309 2975 400367 2981
rect 400309 2972 400321 2975
rect 396040 2944 400321 2972
rect 396040 2932 396046 2944
rect 400309 2941 400321 2944
rect 400355 2941 400367 2975
rect 400309 2935 400367 2941
rect 410518 2932 410524 2984
rect 410576 2972 410582 2984
rect 410576 2944 412496 2972
rect 410576 2932 410582 2944
rect 311032 2876 322796 2904
rect 311032 2864 311038 2876
rect 322842 2864 322848 2916
rect 322900 2904 322906 2916
rect 326525 2907 326583 2913
rect 326525 2904 326537 2907
rect 322900 2876 326537 2904
rect 322900 2864 322906 2876
rect 326525 2873 326537 2876
rect 326571 2873 326583 2907
rect 326525 2867 326583 2873
rect 326617 2907 326675 2913
rect 326617 2873 326629 2907
rect 326663 2904 326675 2907
rect 327718 2904 327724 2916
rect 326663 2876 327724 2904
rect 326663 2873 326675 2876
rect 326617 2867 326675 2873
rect 327718 2864 327724 2876
rect 327776 2864 327782 2916
rect 331214 2864 331220 2916
rect 331272 2904 331278 2916
rect 345658 2904 345664 2916
rect 331272 2876 345664 2904
rect 331272 2864 331278 2876
rect 345658 2864 345664 2876
rect 345716 2864 345722 2916
rect 392578 2864 392584 2916
rect 392636 2904 392642 2916
rect 396626 2904 396632 2916
rect 392636 2876 396632 2904
rect 392636 2864 392642 2876
rect 396626 2864 396632 2876
rect 396684 2864 396690 2916
rect 399478 2864 399484 2916
rect 399536 2904 399542 2916
rect 410886 2904 410892 2916
rect 399536 2876 410892 2904
rect 399536 2864 399542 2876
rect 410886 2864 410892 2876
rect 410944 2864 410950 2916
rect 412468 2904 412496 2944
rect 412542 2932 412548 2984
rect 412600 2972 412606 2984
rect 422297 2975 422355 2981
rect 422297 2972 422309 2975
rect 412600 2944 422309 2972
rect 412600 2932 412606 2944
rect 422297 2941 422309 2944
rect 422343 2941 422355 2975
rect 422297 2935 422355 2941
rect 441985 2975 442043 2981
rect 441985 2941 441997 2975
rect 442031 2972 442043 2975
rect 446582 2972 446588 2984
rect 442031 2944 446588 2972
rect 442031 2941 442043 2944
rect 441985 2935 442043 2941
rect 446582 2932 446588 2944
rect 446640 2932 446646 2984
rect 446677 2975 446735 2981
rect 446677 2941 446689 2975
rect 446723 2972 446735 2975
rect 482278 2972 482284 2984
rect 446723 2944 482284 2972
rect 446723 2941 446735 2944
rect 446677 2935 446735 2941
rect 482278 2932 482284 2944
rect 482336 2932 482342 2984
rect 422389 2907 422447 2913
rect 422389 2904 422401 2907
rect 412468 2876 422401 2904
rect 422389 2873 422401 2876
rect 422435 2873 422447 2907
rect 422389 2867 422447 2873
rect 432509 2907 432567 2913
rect 432509 2873 432521 2907
rect 432555 2904 432567 2907
rect 442169 2907 442227 2913
rect 442169 2904 442181 2907
rect 432555 2876 442181 2904
rect 432555 2873 432567 2876
rect 432509 2867 432567 2873
rect 442169 2873 442181 2876
rect 442215 2873 442227 2907
rect 442169 2867 442227 2873
rect 442258 2864 442264 2916
rect 442316 2904 442322 2916
rect 446309 2907 446367 2913
rect 446309 2904 446321 2907
rect 442316 2876 446321 2904
rect 442316 2864 442322 2876
rect 446309 2873 446321 2876
rect 446355 2873 446367 2907
rect 456153 2907 456211 2913
rect 456153 2904 456165 2907
rect 446309 2867 446367 2873
rect 447980 2876 456165 2904
rect 114796 2808 121592 2836
rect 114796 2796 114802 2808
rect 121822 2796 121828 2848
rect 121880 2836 121886 2848
rect 258810 2836 258816 2848
rect 121880 2808 258816 2836
rect 121880 2796 121886 2808
rect 258810 2796 258816 2808
rect 258868 2796 258874 2848
rect 308582 2796 308588 2848
rect 308640 2836 308646 2848
rect 316678 2836 316684 2848
rect 308640 2808 316684 2836
rect 308640 2796 308646 2808
rect 316678 2796 316684 2808
rect 316736 2796 316742 2848
rect 318058 2796 318064 2848
rect 318116 2836 318122 2848
rect 326341 2839 326399 2845
rect 326341 2836 326353 2839
rect 318116 2808 326353 2836
rect 318116 2796 318122 2808
rect 326341 2805 326353 2808
rect 326387 2805 326399 2839
rect 326341 2799 326399 2805
rect 326430 2796 326436 2848
rect 326488 2836 326494 2848
rect 335265 2839 335323 2845
rect 335265 2836 335277 2839
rect 326488 2808 335277 2836
rect 326488 2796 326494 2808
rect 335265 2805 335277 2808
rect 335311 2805 335323 2839
rect 335265 2799 335323 2805
rect 335906 2796 335912 2848
rect 335964 2836 335970 2848
rect 356514 2836 356520 2848
rect 335964 2808 356520 2836
rect 335964 2796 335970 2808
rect 356514 2796 356520 2808
rect 356572 2796 356578 2848
rect 393958 2796 393964 2848
rect 394016 2836 394022 2848
rect 404906 2836 404912 2848
rect 394016 2808 404912 2836
rect 394016 2796 394022 2808
rect 404906 2796 404912 2808
rect 404964 2796 404970 2848
rect 406378 2796 406384 2848
rect 406436 2836 406442 2848
rect 442994 2836 443000 2848
rect 406436 2808 443000 2836
rect 406436 2796 406442 2808
rect 442994 2796 443000 2808
rect 443052 2796 443058 2848
rect 445662 2796 445668 2848
rect 445720 2836 445726 2848
rect 447980 2836 448008 2876
rect 456153 2873 456165 2876
rect 456199 2873 456211 2907
rect 456153 2867 456211 2873
rect 473906 2836 473912 2848
rect 445720 2808 448008 2836
rect 448072 2808 473912 2836
rect 445720 2796 445726 2808
rect 102781 2771 102839 2777
rect 102781 2768 102793 2771
rect 97368 2740 102793 2768
rect 102781 2737 102793 2740
rect 102827 2737 102839 2771
rect 102781 2731 102839 2737
rect 446309 2771 446367 2777
rect 446309 2737 446321 2771
rect 446355 2768 446367 2771
rect 448072 2768 448100 2808
rect 473906 2796 473912 2808
rect 473964 2796 473970 2848
rect 446355 2740 448100 2768
rect 446355 2737 446367 2740
rect 446309 2731 446367 2737
rect 23106 552 23112 604
rect 23164 592 23170 604
rect 23382 592 23388 604
rect 23164 564 23388 592
rect 23164 552 23170 564
rect 23382 552 23388 564
rect 23440 552 23446 604
rect 148042 552 148048 604
rect 148100 592 148106 604
rect 148962 592 148968 604
rect 148100 564 148968 592
rect 148100 552 148106 564
rect 148962 552 148968 564
rect 149020 552 149026 604
rect 151538 552 151544 604
rect 151596 592 151602 604
rect 151722 592 151728 604
rect 151596 564 151728 592
rect 151596 552 151602 564
rect 151722 552 151728 564
rect 151780 552 151786 604
rect 153930 552 153936 604
rect 153988 592 153994 604
rect 154482 592 154488 604
rect 153988 564 154488 592
rect 153988 552 153994 564
rect 154482 552 154488 564
rect 154540 552 154546 604
rect 155126 552 155132 604
rect 155184 592 155190 604
rect 155862 592 155868 604
rect 155184 564 155868 592
rect 155184 552 155190 564
rect 155862 552 155868 564
rect 155920 552 155926 604
rect 157518 552 157524 604
rect 157576 592 157582 604
rect 158622 592 158628 604
rect 157576 564 158628 592
rect 157576 552 157582 564
rect 158622 552 158628 564
rect 158680 552 158686 604
rect 161106 552 161112 604
rect 161164 592 161170 604
rect 161382 592 161388 604
rect 161164 564 161388 592
rect 161164 552 161170 564
rect 161382 552 161388 564
rect 161440 552 161446 604
rect 171778 552 171784 604
rect 171836 592 171842 604
rect 172422 592 172428 604
rect 171836 564 172428 592
rect 171836 552 171842 564
rect 172422 552 172428 564
rect 172480 552 172486 604
rect 172974 552 172980 604
rect 173032 592 173038 604
rect 173802 592 173808 604
rect 173032 564 173808 592
rect 173032 552 173038 564
rect 173802 552 173808 564
rect 173860 552 173866 604
rect 178954 552 178960 604
rect 179012 592 179018 604
rect 179322 592 179328 604
rect 179012 564 179328 592
rect 179012 552 179018 564
rect 179322 552 179328 564
rect 179380 552 179386 604
rect 180150 552 180156 604
rect 180208 592 180214 604
rect 180702 592 180708 604
rect 180208 564 180708 592
rect 180208 552 180214 564
rect 180702 552 180708 564
rect 180760 552 180766 604
rect 182542 552 182548 604
rect 182600 592 182606 604
rect 183462 592 183468 604
rect 182600 564 183468 592
rect 182600 552 182606 564
rect 183462 552 183468 564
rect 183520 552 183526 604
rect 183738 552 183744 604
rect 183796 592 183802 604
rect 184750 592 184756 604
rect 183796 564 184756 592
rect 183796 552 183802 564
rect 184750 552 184756 564
rect 184808 552 184814 604
rect 189626 552 189632 604
rect 189684 592 189690 604
rect 190362 592 190368 604
rect 189684 564 190368 592
rect 189684 552 189690 564
rect 190362 552 190368 564
rect 190420 552 190426 604
rect 190822 552 190828 604
rect 190880 592 190886 604
rect 191742 592 191748 604
rect 190880 564 191748 592
rect 190880 552 190886 564
rect 191742 552 191748 564
rect 191800 552 191806 604
rect 196802 552 196808 604
rect 196860 592 196866 604
rect 197262 592 197268 604
rect 196860 564 197268 592
rect 196860 552 196866 564
rect 197262 552 197268 564
rect 197320 552 197326 604
rect 197998 552 198004 604
rect 198056 592 198062 604
rect 198642 592 198648 604
rect 198056 564 198648 592
rect 198056 552 198062 564
rect 198642 552 198648 564
rect 198700 552 198706 604
rect 217042 552 217048 604
rect 217100 592 217106 604
rect 217962 592 217968 604
rect 217100 564 217968 592
rect 217100 552 217106 564
rect 217962 552 217968 564
rect 218020 552 218026 604
rect 220538 552 220544 604
rect 220596 592 220602 604
rect 220722 592 220728 604
rect 220596 564 220728 592
rect 220596 552 220602 564
rect 220722 552 220728 564
rect 220780 552 220786 604
rect 224126 552 224132 604
rect 224184 592 224190 604
rect 224862 592 224868 604
rect 224184 564 224868 592
rect 224184 552 224190 564
rect 224862 552 224868 564
rect 224920 552 224926 604
rect 358538 552 358544 604
rect 358596 592 358602 604
rect 358722 592 358728 604
rect 358596 564 358728 592
rect 358596 552 358602 564
rect 358722 552 358728 564
rect 358780 552 358786 604
rect 379606 552 379612 604
rect 379664 592 379670 604
rect 379974 592 379980 604
rect 379664 564 379980 592
rect 379664 552 379670 564
rect 379974 552 379980 564
rect 380032 552 380038 604
rect 492674 552 492680 604
rect 492732 592 492738 604
rect 492950 592 492956 604
rect 492732 564 492956 592
rect 492732 552 492738 564
rect 492950 552 492956 564
rect 493008 552 493014 604
<< via1 >>
rect 328368 700952 328420 701004
rect 478512 700952 478564 701004
rect 170312 700884 170364 700936
rect 351920 700884 351972 700936
rect 154120 700816 154172 700868
rect 356060 700816 356112 700868
rect 320088 700748 320140 700800
rect 527180 700748 527232 700800
rect 137836 700680 137888 700732
rect 353300 700680 353352 700732
rect 321468 700612 321520 700664
rect 543464 700612 543516 700664
rect 105452 700544 105504 700596
rect 357440 700544 357492 700596
rect 89168 700476 89220 700528
rect 361580 700476 361632 700528
rect 72976 700408 73028 700460
rect 358820 700408 358872 700460
rect 40500 700340 40552 700392
rect 362960 700340 363012 700392
rect 24308 700272 24360 700324
rect 367100 700272 367152 700324
rect 202788 700204 202840 700256
rect 347872 700204 347924 700256
rect 348424 700204 348476 700256
rect 364984 700204 365036 700256
rect 325608 700136 325660 700188
rect 462320 700136 462372 700188
rect 218980 700068 219032 700120
rect 349160 700068 349212 700120
rect 235172 700000 235224 700052
rect 346400 700000 346452 700052
rect 333888 699932 333940 699984
rect 413652 699932 413704 699984
rect 267648 699864 267700 699916
rect 342260 699864 342312 699916
rect 331128 699796 331180 699848
rect 397460 699796 397512 699848
rect 283840 699728 283892 699780
rect 343640 699728 343692 699780
rect 300124 699660 300176 699712
rect 300768 699660 300820 699712
rect 332508 699660 332560 699712
rect 336740 699660 336792 699712
rect 339408 699660 339460 699712
rect 348792 699660 348844 699712
rect 314568 696940 314620 696992
rect 580172 696940 580224 696992
rect 429384 688576 429436 688628
rect 429844 688576 429896 688628
rect 559104 688576 559156 688628
rect 559656 688576 559708 688628
rect 315948 685856 316000 685908
rect 580172 685856 580224 685908
rect 429292 684428 429344 684480
rect 559012 684428 559064 684480
rect 3516 681708 3568 681760
rect 368480 681708 368532 681760
rect 494060 676175 494112 676184
rect 494060 676141 494069 676175
rect 494069 676141 494103 676175
rect 494103 676141 494112 676175
rect 494060 676132 494112 676141
rect 311808 673480 311860 673532
rect 580172 673480 580224 673532
rect 3424 667904 3476 667956
rect 372620 667904 372672 667956
rect 429660 666544 429712 666596
rect 494152 666544 494204 666596
rect 559380 666544 559432 666596
rect 494060 654100 494112 654152
rect 494244 654100 494296 654152
rect 3056 652740 3108 652792
rect 371240 652740 371292 652792
rect 309048 650020 309100 650072
rect 580172 650020 580224 650072
rect 429384 647232 429436 647284
rect 429476 647232 429528 647284
rect 559104 647232 559156 647284
rect 559196 647232 559248 647284
rect 429384 640364 429436 640416
rect 429476 640364 429528 640416
rect 559104 640364 559156 640416
rect 559196 640364 559248 640416
rect 310428 638936 310480 638988
rect 580172 638936 580224 638988
rect 494060 634788 494112 634840
rect 494244 634788 494296 634840
rect 429292 630640 429344 630692
rect 429476 630640 429528 630692
rect 559012 630640 559064 630692
rect 559196 630640 559248 630692
rect 306288 626560 306340 626612
rect 580172 626560 580224 626612
rect 3424 623772 3476 623824
rect 375380 623772 375432 623824
rect 494060 615476 494112 615528
rect 494244 615476 494296 615528
rect 429292 611328 429344 611380
rect 429476 611328 429528 611380
rect 559012 611328 559064 611380
rect 559196 611328 559248 611380
rect 3424 609968 3476 610020
rect 378140 609968 378192 610020
rect 429384 608583 429436 608592
rect 429384 608549 429393 608583
rect 429393 608549 429427 608583
rect 429427 608549 429436 608583
rect 429384 608540 429436 608549
rect 559104 608583 559156 608592
rect 559104 608549 559113 608583
rect 559113 608549 559147 608583
rect 559147 608549 559156 608583
rect 559104 608540 559156 608549
rect 302148 603100 302200 603152
rect 580172 603100 580224 603152
rect 429568 601672 429620 601724
rect 559288 601672 559340 601724
rect 429568 598927 429620 598936
rect 429568 598893 429577 598927
rect 429577 598893 429611 598927
rect 429611 598893 429620 598927
rect 429568 598884 429620 598893
rect 559288 598927 559340 598936
rect 559288 598893 559297 598927
rect 559297 598893 559331 598927
rect 559331 598893 559340 598927
rect 559288 598884 559340 598893
rect 494060 596164 494112 596216
rect 494244 596164 494296 596216
rect 3240 594804 3292 594856
rect 376760 594804 376812 594856
rect 304908 592016 304960 592068
rect 580172 592016 580224 592068
rect 429660 589296 429712 589348
rect 559380 589296 559432 589348
rect 300676 579640 300728 579692
rect 580172 579640 580224 579692
rect 429568 579572 429620 579624
rect 494060 579615 494112 579624
rect 494060 579581 494069 579615
rect 494069 579581 494103 579615
rect 494103 579581 494112 579615
rect 494060 579572 494112 579581
rect 559288 579615 559340 579624
rect 559288 579581 559297 579615
rect 559297 579581 559331 579615
rect 559331 579581 559340 579615
rect 559288 579572 559340 579581
rect 429476 569959 429528 569968
rect 429476 569925 429485 569959
rect 429485 569925 429519 569959
rect 429519 569925 429528 569959
rect 429476 569916 429528 569925
rect 494244 569916 494296 569968
rect 559380 569916 559432 569968
rect 3424 567196 3476 567248
rect 380900 567196 380952 567248
rect 307760 565088 307812 565140
rect 309048 565088 309100 565140
rect 309140 565088 309192 565140
rect 310428 565088 310480 565140
rect 310520 565088 310572 565140
rect 311808 565088 311860 565140
rect 313280 565088 313332 565140
rect 314568 565088 314620 565140
rect 314660 565088 314712 565140
rect 315948 565088 316000 565140
rect 327080 565088 327132 565140
rect 328368 565088 328420 565140
rect 329840 565088 329892 565140
rect 331128 565088 331180 565140
rect 332600 565088 332652 565140
rect 333888 565088 333940 565140
rect 333980 563932 334032 563984
rect 348424 563932 348476 563984
rect 300768 563864 300820 563916
rect 340696 563864 340748 563916
rect 328460 563796 328512 563848
rect 429476 563796 429528 563848
rect 323308 563728 323360 563780
rect 494244 563728 494296 563780
rect 317512 563660 317564 563712
rect 559380 563660 559432 563712
rect 289820 562980 289872 563032
rect 298284 562912 298336 562964
rect 412088 562980 412140 563032
rect 310520 562912 310572 562964
rect 311716 562912 311768 562964
rect 450452 562912 450504 562964
rect 255780 562844 255832 562896
rect 286968 562844 287020 562896
rect 292488 562844 292540 562896
rect 450360 562844 450412 562896
rect 284760 562776 284812 562828
rect 451096 562776 451148 562828
rect 280896 562708 280948 562760
rect 450728 562708 450780 562760
rect 278964 562640 279016 562692
rect 451004 562640 451056 562692
rect 261576 562572 261628 562624
rect 278780 562572 278832 562624
rect 286692 562572 286744 562624
rect 462964 562572 463016 562624
rect 273168 562504 273220 562556
rect 450636 562504 450688 562556
rect 259644 562436 259696 562488
rect 580908 562436 580960 562488
rect 6552 562368 6604 562420
rect 388904 562368 388956 562420
rect 3056 562300 3108 562352
rect 386972 562300 387024 562352
rect 6644 562232 6696 562284
rect 390836 562232 390888 562284
rect 3148 562164 3200 562216
rect 392768 562164 392820 562216
rect 5448 562096 5500 562148
rect 394700 562096 394752 562148
rect 417884 562096 417936 562148
rect 6460 562028 6512 562080
rect 396632 562028 396684 562080
rect 3240 561960 3292 562012
rect 398564 561960 398616 562012
rect 5356 561892 5408 561944
rect 400496 561892 400548 561944
rect 6368 561824 6420 561876
rect 402428 561824 402480 561876
rect 3332 561756 3384 561808
rect 408224 561756 408276 561808
rect 6276 561688 6328 561740
rect 414020 561688 414072 561740
rect 390652 561008 390704 561060
rect 4068 560940 4120 560992
rect 289820 560940 289872 560992
rect 296352 560940 296404 560992
rect 450820 560940 450872 560992
rect 290556 560872 290608 560924
rect 451188 560872 451240 560924
rect 282828 560804 282880 560856
rect 450268 560804 450320 560856
rect 277032 560736 277084 560788
rect 400220 560736 400272 560788
rect 400588 560736 400640 560788
rect 449624 560736 449676 560788
rect 271236 560668 271288 560720
rect 450544 560668 450596 560720
rect 286968 560600 287020 560652
rect 294420 560600 294472 560652
rect 548524 560600 548576 560652
rect 5264 560532 5316 560584
rect 410156 560532 410208 560584
rect 411352 560532 411404 560584
rect 424324 560532 424376 560584
rect 5172 560464 5224 560516
rect 421748 560464 421800 560516
rect 4988 560396 5040 560448
rect 427544 560396 427596 560448
rect 4804 560328 4856 560380
rect 400220 560328 400272 560380
rect 400588 560328 400640 560380
rect 433340 560328 433392 560380
rect 6184 560260 6236 560312
rect 439136 560260 439188 560312
rect 400220 560192 400272 560244
rect 400588 560192 400640 560244
rect 579804 560192 579856 560244
rect 278780 560124 278832 560176
rect 580080 560124 580132 560176
rect 275100 560056 275152 560108
rect 400220 560056 400272 560108
rect 400588 560056 400640 560108
rect 579896 560056 579948 560108
rect 269672 559988 269724 560040
rect 579988 559988 580040 560040
rect 267648 559920 267700 559972
rect 400220 559920 400272 559972
rect 400588 559920 400640 559972
rect 577596 559920 577648 559972
rect 265808 559852 265860 559904
rect 372252 559852 372304 559904
rect 389088 559852 389140 559904
rect 400312 559852 400364 559904
rect 400680 559852 400732 559904
rect 409880 559852 409932 559904
rect 419356 559852 419408 559904
rect 577504 559852 577556 559904
rect 263600 559784 263652 559836
rect 580172 559784 580224 559836
rect 3884 559716 3936 559768
rect 390560 559716 390612 559768
rect 258080 559648 258132 559700
rect 580724 559648 580776 559700
rect 5540 559376 5592 559428
rect 248788 559580 248840 559632
rect 252192 559580 252244 559632
rect 580632 559580 580684 559632
rect 246488 559512 246540 559564
rect 580448 559512 580500 559564
rect 240140 559444 240192 559496
rect 240600 559444 240652 559496
rect 580264 559444 580316 559496
rect 3700 559308 3752 559360
rect 384856 559376 384908 559428
rect 369860 559308 369912 559360
rect 396356 559376 396408 559428
rect 385132 559308 385184 559360
rect 396080 559308 396132 559360
rect 434996 559376 435048 559428
rect 431132 559308 431184 559360
rect 3516 559104 3568 559156
rect 450820 557472 450872 557524
rect 579712 557472 579764 557524
rect 450268 557268 450320 557320
rect 450912 557268 450964 557320
rect 450360 557132 450412 557184
rect 451096 557132 451148 557184
rect 2780 553052 2832 553104
rect 5540 553052 5592 553104
rect 579804 552644 579856 552696
rect 580816 552644 580868 552696
rect 450452 546388 450504 546440
rect 579804 546388 579856 546440
rect 548524 534012 548576 534064
rect 579804 534012 579856 534064
rect 451188 510552 451240 510604
rect 579804 510552 579856 510604
rect 451096 499468 451148 499520
rect 579804 499468 579856 499520
rect 3056 495524 3108 495576
rect 6644 495524 6696 495576
rect 3056 481108 3108 481160
rect 6552 481108 6604 481160
rect 451004 463632 451056 463684
rect 579804 463632 579856 463684
rect 462964 452548 463016 452600
rect 579804 452548 579856 452600
rect 450912 440172 450964 440224
rect 579804 440172 579856 440224
rect 3148 438676 3200 438728
rect 6460 438676 6512 438728
rect 2780 424668 2832 424720
rect 5448 424668 5500 424720
rect 450820 416712 450872 416764
rect 579804 416712 579856 416764
rect 450728 405628 450780 405680
rect 579804 405628 579856 405680
rect 449716 393252 449768 393304
rect 579804 393252 579856 393304
rect 3148 380604 3200 380656
rect 6368 380604 6420 380656
rect 450636 369792 450688 369844
rect 579804 369792 579856 369844
rect 2780 366936 2832 366988
rect 5356 366936 5408 366988
rect 450544 346332 450596 346384
rect 579896 346332 579948 346384
rect 363052 340076 363104 340128
rect 363880 340076 363932 340128
rect 345204 339056 345256 339108
rect 345756 339056 345808 339108
rect 270592 338376 270644 338428
rect 271236 338376 271288 338428
rect 239128 338104 239180 338156
rect 239864 338104 239916 338156
rect 79324 338036 79376 338088
rect 258264 338036 258316 338088
rect 292488 338036 292540 338088
rect 341800 338036 341852 338088
rect 348240 338036 348292 338088
rect 349804 338036 349856 338088
rect 71044 337968 71096 338020
rect 250168 337968 250220 338020
rect 263600 337968 263652 338020
rect 335912 337968 335964 338020
rect 344468 337968 344520 338020
rect 349068 337968 349120 338020
rect 357440 338036 357492 338088
rect 363052 338036 363104 338088
rect 363144 338036 363196 338088
rect 377680 338036 377732 338088
rect 360200 337968 360252 338020
rect 376300 337968 376352 338020
rect 66904 337900 66956 337952
rect 245660 337900 245712 337952
rect 251824 337900 251876 337952
rect 256884 337900 256936 337952
rect 259552 337900 259604 337952
rect 266360 337900 266412 337952
rect 334532 337900 334584 337952
rect 334716 337900 334768 337952
rect 345388 337900 345440 337952
rect 345756 337900 345808 337952
rect 351644 337900 351696 337952
rect 351828 337900 351880 337952
rect 61384 337832 61436 337884
rect 246120 337832 246172 337884
rect 250444 337832 250496 337884
rect 254216 337832 254268 337884
rect 57244 337764 57296 337816
rect 242992 337764 243044 337816
rect 339960 337832 340012 337884
rect 349436 337832 349488 337884
rect 352012 337832 352064 337884
rect 352748 337832 352800 337884
rect 361028 337900 361080 337952
rect 379428 337900 379480 337952
rect 384856 338036 384908 338088
rect 418528 338036 418580 338088
rect 431040 338104 431092 338156
rect 431224 338036 431276 338088
rect 434076 338104 434128 338156
rect 502984 338036 503036 338088
rect 390284 337968 390336 338020
rect 397000 337968 397052 338020
rect 406384 337968 406436 338020
rect 421196 337968 421248 338020
rect 500224 337968 500276 338020
rect 355324 337832 355376 337884
rect 359280 337832 359332 337884
rect 370044 337832 370096 337884
rect 371056 337832 371108 337884
rect 380808 337832 380860 337884
rect 393964 337900 394016 337952
rect 388444 337832 388496 337884
rect 395344 337832 395396 337884
rect 254584 337764 254636 337816
rect 42064 337696 42116 337748
rect 233976 337696 234028 337748
rect 260932 337764 260984 337816
rect 285588 337764 285640 337816
rect 337292 337764 337344 337816
rect 344008 337764 344060 337816
rect 344928 337764 344980 337816
rect 359740 337764 359792 337816
rect 374552 337764 374604 337816
rect 376024 337764 376076 337816
rect 276756 337696 276808 337748
rect 329656 337696 329708 337748
rect 331128 337696 331180 337748
rect 39304 337628 39356 337680
rect 243452 337628 243504 337680
rect 254860 337628 254912 337680
rect 259460 337628 259512 337680
rect 35164 337560 35216 337612
rect 240784 337560 240836 337612
rect 258816 337560 258868 337612
rect 275744 337560 275796 337612
rect 276664 337560 276716 337612
rect 333704 337628 333756 337680
rect 330392 337560 330444 337612
rect 330484 337560 330536 337612
rect 352564 337696 352616 337748
rect 353392 337696 353444 337748
rect 356704 337696 356756 337748
rect 360568 337696 360620 337748
rect 372252 337696 372304 337748
rect 373264 337696 373316 337748
rect 374092 337696 374144 337748
rect 375288 337696 375340 337748
rect 377220 337696 377272 337748
rect 377956 337696 378008 337748
rect 379888 337696 379940 337748
rect 380808 337696 380860 337748
rect 381268 337696 381320 337748
rect 382188 337696 382240 337748
rect 382648 337764 382700 337816
rect 393872 337764 393924 337816
rect 394424 337764 394476 337816
rect 383936 337696 383988 337748
rect 384948 337696 385000 337748
rect 389364 337696 389416 337748
rect 390468 337696 390520 337748
rect 399484 337900 399536 337952
rect 406752 337900 406804 337952
rect 398288 337832 398340 337884
rect 409144 337832 409196 337884
rect 415860 337900 415912 337952
rect 427176 337900 427228 337952
rect 428464 337900 428516 337952
rect 429108 337900 429160 337952
rect 417424 337832 417476 337884
rect 423864 337832 423916 337884
rect 340788 337628 340840 337680
rect 358360 337628 358412 337680
rect 372712 337628 372764 337680
rect 373908 337628 373960 337680
rect 375840 337628 375892 337680
rect 377404 337628 377456 337680
rect 378600 337628 378652 337680
rect 380164 337628 380216 337680
rect 380348 337628 380400 337680
rect 399116 337764 399168 337816
rect 403716 337764 403768 337816
rect 411904 337764 411956 337816
rect 396540 337696 396592 337748
rect 397276 337696 397328 337748
rect 397828 337696 397880 337748
rect 398564 337696 398616 337748
rect 399208 337696 399260 337748
rect 400036 337696 400088 337748
rect 400588 337696 400640 337748
rect 401416 337696 401468 337748
rect 401876 337696 401928 337748
rect 402796 337696 402848 337748
rect 403256 337696 403308 337748
rect 404176 337696 404228 337748
rect 404636 337696 404688 337748
rect 405556 337696 405608 337748
rect 405924 337696 405976 337748
rect 406936 337696 406988 337748
rect 407304 337696 407356 337748
rect 408316 337696 408368 337748
rect 409052 337696 409104 337748
rect 420184 337764 420236 337816
rect 422576 337764 422628 337816
rect 414020 337696 414072 337748
rect 415308 337696 415360 337748
rect 423036 337696 423088 337748
rect 423588 337696 423640 337748
rect 424324 337696 424376 337748
rect 424968 337696 425020 337748
rect 396080 337628 396132 337680
rect 397368 337628 397420 337680
rect 397460 337628 397512 337680
rect 398656 337628 398708 337680
rect 401048 337628 401100 337680
rect 410524 337628 410576 337680
rect 412640 337628 412692 337680
rect 413928 337628 413980 337680
rect 414480 337628 414532 337680
rect 417148 337628 417200 337680
rect 425704 337696 425756 337748
rect 426348 337696 426400 337748
rect 426624 337764 426676 337816
rect 507124 337900 507176 337952
rect 437388 337832 437440 337884
rect 514024 337832 514076 337884
rect 511264 337764 511316 337816
rect 426992 337696 427044 337748
rect 427084 337696 427136 337748
rect 427728 337696 427780 337748
rect 427912 337696 427964 337748
rect 429108 337696 429160 337748
rect 429292 337696 429344 337748
rect 425244 337628 425296 337680
rect 429844 337628 429896 337680
rect 431960 337696 432012 337748
rect 438768 337696 438820 337748
rect 444104 337696 444156 337748
rect 436376 337628 436428 337680
rect 436468 337628 436520 337680
rect 437388 337628 437440 337680
rect 441436 337628 441488 337680
rect 444840 337628 444892 337680
rect 445944 337628 445996 337680
rect 447048 337628 447100 337680
rect 356980 337560 357032 337612
rect 358084 337560 358136 337612
rect 363328 337560 363380 337612
rect 375380 337560 375432 337612
rect 376668 337560 376720 337612
rect 379060 337560 379112 337612
rect 381636 337560 381688 337612
rect 28264 337492 28316 337544
rect 19984 337424 20036 337476
rect 237564 337492 237616 337544
rect 258724 337492 258776 337544
rect 273076 337492 273128 337544
rect 274548 337492 274600 337544
rect 333244 337492 333296 337544
rect 334624 337492 334676 337544
rect 348424 337492 348476 337544
rect 353208 337492 353260 337544
rect 362408 337492 362460 337544
rect 371424 337492 371476 337544
rect 374092 337492 374144 337544
rect 378140 337492 378192 337544
rect 384304 337492 384356 337544
rect 386604 337560 386656 337612
rect 387524 337560 387576 337612
rect 390652 337560 390704 337612
rect 391664 337560 391716 337612
rect 392032 337560 392084 337612
rect 393044 337560 393096 337612
rect 387064 337492 387116 337544
rect 387984 337492 388036 337544
rect 407764 337560 407816 337612
rect 408684 337560 408736 337612
rect 438216 337560 438268 337612
rect 518164 337696 518216 337748
rect 447232 337628 447284 337680
rect 448428 337628 448480 337680
rect 448612 337628 448664 337680
rect 449808 337628 449860 337680
rect 447324 337560 447376 337612
rect 529204 337628 529256 337680
rect 527824 337560 527876 337612
rect 405096 337492 405148 337544
rect 411812 337492 411864 337544
rect 237196 337424 237248 337476
rect 13084 337356 13136 337408
rect 233608 337356 233660 337408
rect 234160 337356 234212 337408
rect 240324 337356 240376 337408
rect 138020 337288 138072 337340
rect 147588 337288 147640 337340
rect 157340 337288 157392 337340
rect 166908 337288 166960 337340
rect 176660 337288 176712 337340
rect 186228 337288 186280 337340
rect 195980 337288 196032 337340
rect 205548 337288 205600 337340
rect 215300 337288 215352 337340
rect 224868 337288 224920 337340
rect 257344 337424 257396 337476
rect 271696 337424 271748 337476
rect 271788 337424 271840 337476
rect 331864 337424 331916 337476
rect 333888 337424 333940 337476
rect 355692 337424 355744 337476
rect 362868 337424 362920 337476
rect 373172 337424 373224 337476
rect 77944 337220 77996 337272
rect 252836 337356 252888 337408
rect 255964 337288 256016 337340
rect 268660 337356 268712 337408
rect 269028 337356 269080 337408
rect 334532 337356 334584 337408
rect 334808 337356 334860 337408
rect 336372 337356 336424 337408
rect 352196 337356 352248 337408
rect 355968 337356 356020 337408
rect 363788 337356 363840 337408
rect 376760 337424 376812 337476
rect 378048 337424 378100 337476
rect 381728 337424 381780 337476
rect 379612 337356 379664 337408
rect 383016 337356 383068 337408
rect 279976 337288 280028 337340
rect 288072 337288 288124 337340
rect 303528 337288 303580 337340
rect 338028 337288 338080 337340
rect 347136 337288 347188 337340
rect 351184 337288 351236 337340
rect 361488 337288 361540 337340
rect 375012 337288 375064 337340
rect 381544 337288 381596 337340
rect 385316 337288 385368 337340
rect 394700 337424 394752 337476
rect 395804 337424 395856 337476
rect 402244 337424 402296 337476
rect 415400 337424 415452 337476
rect 416596 337424 416648 337476
rect 433984 337492 434036 337544
rect 433340 337424 433392 337476
rect 435088 337424 435140 337476
rect 444840 337492 444892 337544
rect 525064 337492 525116 337544
rect 520924 337424 520976 337476
rect 405004 337356 405056 337408
rect 411352 337356 411404 337408
rect 428372 337356 428424 337408
rect 429108 337356 429160 337408
rect 429752 337356 429804 337408
rect 430488 337356 430540 337408
rect 431132 337356 431184 337408
rect 431868 337356 431920 337408
rect 432420 337356 432472 337408
rect 433248 337356 433300 337408
rect 433800 337356 433852 337408
rect 434628 337356 434680 337408
rect 436008 337356 436060 337408
rect 436836 337356 436888 337408
rect 437848 337356 437900 337408
rect 438768 337356 438820 337408
rect 439136 337356 439188 337408
rect 440056 337356 440108 337408
rect 440516 337356 440568 337408
rect 441528 337356 441580 337408
rect 441896 337356 441948 337408
rect 442816 337356 442868 337408
rect 443184 337356 443236 337408
rect 444288 337356 444340 337408
rect 444564 337356 444616 337408
rect 445576 337356 445628 337408
rect 523684 337356 523736 337408
rect 401876 337288 401928 337340
rect 496084 337288 496136 337340
rect 246304 337220 246356 337272
rect 247040 337220 247092 337272
rect 247776 337220 247828 337272
rect 248788 337220 248840 337272
rect 249064 337220 249116 337272
rect 251548 337220 251600 337272
rect 253204 337220 253256 337272
rect 259644 337220 259696 337272
rect 305828 337220 305880 337272
rect 97264 337152 97316 337204
rect 264980 337152 265032 337204
rect 297916 337152 297968 337204
rect 312728 337152 312780 337204
rect 84844 337084 84896 337136
rect 100668 337084 100720 337136
rect 267648 337084 267700 337136
rect 321468 337084 321520 337136
rect 350724 337220 350776 337272
rect 392584 337220 392636 337272
rect 408040 337220 408092 337272
rect 419908 337220 419960 337272
rect 421564 337220 421616 337272
rect 492680 337220 492732 337272
rect 341340 337152 341392 337204
rect 345664 337152 345716 337204
rect 354772 337152 354824 337204
rect 365536 337152 365588 337204
rect 370504 337152 370556 337204
rect 372712 337152 372764 337204
rect 413100 337152 413152 337204
rect 485780 337152 485832 337204
rect 107568 337016 107620 337068
rect 270408 337016 270460 337068
rect 105544 336948 105596 337000
rect 262312 336948 262364 337000
rect 319536 336948 319588 337000
rect 343088 337084 343140 337136
rect 339040 337016 339092 337068
rect 346676 337084 346728 337136
rect 358728 337084 358780 337136
rect 365076 337084 365128 337136
rect 393412 337084 393464 337136
rect 394516 337084 394568 337136
rect 399668 337084 399720 337136
rect 410432 337084 410484 337136
rect 477500 337084 477552 337136
rect 327724 336948 327776 337000
rect 118608 336880 118660 336932
rect 274456 336880 274508 336932
rect 316776 336880 316828 336932
rect 102784 336812 102836 336864
rect 255596 336812 255648 336864
rect 326344 336812 326396 336864
rect 338764 336812 338816 336864
rect 353852 337016 353904 337068
rect 359464 337016 359516 337068
rect 364616 337016 364668 337068
rect 371792 337016 371844 337068
rect 375656 337016 375708 337068
rect 389824 337016 389876 337068
rect 390376 337016 390428 337068
rect 409972 337016 410024 337068
rect 477592 337016 477644 337068
rect 341984 336948 342036 337000
rect 348056 336948 348108 337000
rect 360108 336948 360160 337000
rect 364248 336948 364300 337000
rect 366916 336948 366968 337000
rect 470600 336948 470652 337000
rect 344744 336880 344796 336932
rect 350264 336880 350316 336932
rect 366364 336880 366416 336932
rect 367376 336880 367428 336932
rect 373632 336880 373684 336932
rect 374644 336880 374696 336932
rect 402336 336880 402388 336932
rect 344652 336812 344704 336864
rect 349344 336812 349396 336864
rect 362224 336812 362276 336864
rect 365996 336812 366048 336864
rect 366916 336812 366968 336864
rect 367836 336812 367888 336864
rect 405372 336880 405424 336932
rect 463700 336880 463752 336932
rect 456800 336812 456852 336864
rect 125508 336744 125560 336796
rect 277124 336744 277176 336796
rect 322296 336744 322348 336796
rect 327816 336744 327868 336796
rect 342628 336744 342680 336796
rect 354312 336744 354364 336796
rect 362868 336744 362920 336796
rect 366456 336744 366508 336796
rect 367008 336744 367060 336796
rect 368204 336744 368256 336796
rect 239128 336719 239180 336728
rect 239128 336685 239137 336719
rect 239137 336685 239171 336719
rect 239171 336685 239180 336719
rect 239128 336676 239180 336685
rect 324688 336719 324740 336728
rect 324688 336685 324697 336719
rect 324697 336685 324731 336719
rect 324731 336685 324740 336719
rect 324688 336676 324740 336685
rect 435364 336676 435416 336728
rect 449900 336676 449952 336728
rect 438124 336608 438176 336660
rect 442264 336472 442316 336524
rect 311900 335724 311952 335776
rect 312268 335724 312320 335776
rect 232044 335656 232096 335708
rect 232780 335656 232832 335708
rect 277400 335656 277452 335708
rect 278136 335656 278188 335708
rect 285864 335656 285916 335708
rect 286692 335656 286744 335708
rect 303712 335656 303764 335708
rect 304632 335656 304684 335708
rect 306472 335656 306524 335708
rect 307300 335656 307352 335708
rect 317420 335656 317472 335708
rect 317604 335656 317656 335708
rect 323032 335656 323084 335708
rect 323492 335656 323544 335708
rect 231952 335588 232004 335640
rect 232412 335588 232464 335640
rect 234712 335588 234764 335640
rect 234988 335588 235040 335640
rect 236092 335588 236144 335640
rect 236460 335588 236512 335640
rect 237472 335588 237524 335640
rect 238116 335588 238168 335640
rect 241520 335588 241572 335640
rect 241796 335588 241848 335640
rect 247132 335588 247184 335640
rect 247684 335588 247736 335640
rect 249892 335588 249944 335640
rect 250812 335588 250864 335640
rect 251272 335588 251324 335640
rect 252100 335588 252152 335640
rect 252652 335588 252704 335640
rect 253388 335588 253440 335640
rect 255412 335588 255464 335640
rect 256148 335588 256200 335640
rect 258172 335588 258224 335640
rect 258908 335588 258960 335640
rect 259552 335588 259604 335640
rect 260196 335588 260248 335640
rect 263692 335588 263744 335640
rect 264244 335588 264296 335640
rect 266452 335588 266504 335640
rect 267004 335588 267056 335640
rect 267832 335588 267884 335640
rect 268292 335588 268344 335640
rect 269212 335588 269264 335640
rect 269580 335588 269632 335640
rect 271972 335588 272024 335640
rect 272340 335588 272392 335640
rect 274732 335588 274784 335640
rect 274916 335588 274968 335640
rect 277492 335588 277544 335640
rect 277676 335588 277728 335640
rect 278964 335588 279016 335640
rect 279516 335588 279568 335640
rect 281724 335588 281776 335640
rect 282184 335588 282236 335640
rect 283012 335588 283064 335640
rect 283564 335588 283616 335640
rect 285772 335588 285824 335640
rect 286140 335588 286192 335640
rect 294052 335588 294104 335640
rect 294788 335588 294840 335640
rect 296812 335588 296864 335640
rect 297364 335588 297416 335640
rect 302332 335588 302384 335640
rect 302884 335588 302936 335640
rect 303804 335588 303856 335640
rect 304172 335588 304224 335640
rect 306380 335588 306432 335640
rect 306932 335588 306984 335640
rect 307760 335588 307812 335640
rect 308220 335588 308272 335640
rect 309140 335588 309192 335640
rect 309508 335588 309560 335640
rect 310520 335588 310572 335640
rect 310980 335588 311032 335640
rect 313280 335588 313332 335640
rect 313556 335588 313608 335640
rect 320272 335588 320324 335640
rect 320732 335588 320784 335640
rect 321652 335588 321704 335640
rect 322204 335588 322256 335640
rect 323216 335588 323268 335640
rect 323860 335588 323912 335640
rect 325792 335588 325844 335640
rect 326620 335588 326672 335640
rect 327172 335588 327224 335640
rect 327908 335588 327960 335640
rect 329932 335588 329984 335640
rect 330300 335588 330352 335640
rect 345112 335588 345164 335640
rect 345940 335588 345992 335640
rect 435456 335588 435508 335640
rect 436008 335588 436060 335640
rect 344560 335520 344612 335572
rect 273536 335384 273588 335436
rect 314660 335248 314712 335300
rect 315028 335248 315080 335300
rect 273444 335180 273496 335232
rect 324412 334976 324464 335028
rect 325332 334976 325384 335028
rect 234068 334432 234120 334484
rect 265072 334296 265124 334348
rect 265532 334296 265584 334348
rect 287980 334296 288032 334348
rect 312176 334296 312228 334348
rect 312636 334296 312688 334348
rect 319444 334160 319496 334212
rect 256792 334024 256844 334076
rect 257436 334024 257488 334076
rect 238668 333276 238720 333328
rect 239036 333276 239088 333328
rect 273352 333276 273404 333328
rect 273628 333276 273680 333328
rect 347872 333276 347924 333328
rect 348700 333276 348752 333328
rect 284392 333140 284444 333192
rect 284852 333140 284904 333192
rect 318800 333140 318852 333192
rect 319076 333140 319128 333192
rect 300952 332800 301004 332852
rect 301412 332800 301464 332852
rect 248604 332392 248656 332444
rect 249340 332392 249392 332444
rect 235448 331916 235500 331968
rect 295432 331576 295484 331628
rect 296076 331576 296128 331628
rect 298468 331440 298520 331492
rect 298928 331440 298980 331492
rect 244464 331304 244516 331356
rect 244372 331236 244424 331288
rect 244280 331168 244332 331220
rect 327448 331211 327500 331220
rect 327448 331177 327457 331211
rect 327457 331177 327491 331211
rect 327491 331177 327500 331211
rect 327448 331168 327500 331177
rect 244372 331100 244424 331152
rect 316040 330964 316092 331016
rect 316316 330964 316368 331016
rect 314936 330216 314988 330268
rect 315396 330216 315448 330268
rect 290464 329400 290516 329452
rect 233516 328491 233568 328500
rect 233516 328457 233525 328491
rect 233525 328457 233559 328491
rect 233559 328457 233568 328491
rect 233516 328448 233568 328457
rect 262680 328448 262732 328500
rect 263048 328448 263100 328500
rect 267004 328491 267056 328500
rect 267004 328457 267013 328491
rect 267013 328457 267047 328491
rect 267047 328457 267056 328491
rect 267004 328448 267056 328457
rect 288808 328448 288860 328500
rect 289544 328448 289596 328500
rect 290004 328448 290056 328500
rect 290648 328448 290700 328500
rect 291568 328448 291620 328500
rect 292120 328448 292172 328500
rect 292764 328448 292816 328500
rect 293592 328448 293644 328500
rect 305368 328448 305420 328500
rect 306104 328448 306156 328500
rect 308128 328448 308180 328500
rect 308680 328448 308732 328500
rect 310888 328448 310940 328500
rect 311440 328448 311492 328500
rect 316408 328448 316460 328500
rect 316592 328448 316644 328500
rect 319168 328491 319220 328500
rect 319168 328457 319177 328491
rect 319177 328457 319211 328491
rect 319211 328457 319220 328491
rect 319168 328448 319220 328457
rect 327448 328491 327500 328500
rect 327448 328457 327457 328491
rect 327457 328457 327491 328491
rect 327491 328457 327500 328491
rect 327448 328448 327500 328457
rect 328552 328448 328604 328500
rect 328828 328448 328880 328500
rect 343824 328491 343876 328500
rect 343824 328457 343833 328491
rect 343833 328457 343867 328491
rect 343867 328457 343876 328491
rect 343824 328448 343876 328457
rect 346584 328448 346636 328500
rect 347320 328448 347372 328500
rect 347964 328491 348016 328500
rect 347964 328457 347973 328491
rect 347973 328457 348007 328491
rect 348007 328457 348016 328491
rect 347964 328448 348016 328457
rect 251456 328380 251508 328432
rect 251640 328380 251692 328432
rect 254216 328380 254268 328432
rect 254308 328380 254360 328432
rect 363236 328423 363288 328432
rect 363236 328389 363245 328423
rect 363245 328389 363279 328423
rect 363279 328389 363288 328423
rect 363236 328380 363288 328389
rect 324780 328312 324832 328364
rect 347964 328355 348016 328364
rect 347964 328321 347973 328355
rect 347973 328321 348007 328355
rect 348007 328321 348016 328355
rect 347964 328312 348016 328321
rect 235080 327131 235132 327140
rect 235080 327097 235089 327131
rect 235089 327097 235123 327131
rect 235123 327097 235132 327131
rect 235080 327088 235132 327097
rect 240416 327088 240468 327140
rect 240876 327088 240928 327140
rect 241888 327088 241940 327140
rect 242164 327088 242216 327140
rect 245936 327088 245988 327140
rect 246212 327088 246264 327140
rect 287428 327131 287480 327140
rect 287428 327097 287437 327131
rect 287437 327097 287471 327131
rect 287471 327097 287480 327131
rect 287428 327088 287480 327097
rect 234804 327063 234856 327072
rect 234804 327029 234813 327063
rect 234813 327029 234847 327063
rect 234847 327029 234856 327063
rect 234804 327020 234856 327029
rect 248880 325660 248932 325712
rect 249248 325660 249300 325712
rect 577596 322872 577648 322924
rect 579896 322872 579948 322924
rect 248788 322192 248840 322244
rect 249248 322192 249300 322244
rect 255688 321580 255740 321632
rect 261208 321580 261260 321632
rect 229284 321512 229336 321564
rect 229468 321512 229520 321564
rect 238760 321512 238812 321564
rect 238944 321512 238996 321564
rect 255688 321376 255740 321428
rect 267096 321580 267148 321632
rect 290004 321580 290056 321632
rect 292764 321580 292816 321632
rect 325976 321580 326028 321632
rect 290096 321444 290148 321496
rect 292856 321444 292908 321496
rect 261300 321376 261352 321428
rect 267004 321376 267056 321428
rect 326068 321376 326120 321428
rect 239128 318835 239180 318844
rect 239128 318801 239137 318835
rect 239137 318801 239171 318835
rect 239171 318801 239180 318835
rect 239128 318792 239180 318801
rect 251640 318860 251692 318912
rect 280528 318792 280580 318844
rect 280620 318792 280672 318844
rect 316408 318860 316460 318912
rect 317880 318860 317932 318912
rect 317788 318792 317840 318844
rect 347964 318835 348016 318844
rect 347964 318801 347973 318835
rect 347973 318801 348007 318835
rect 348007 318801 348016 318835
rect 347964 318792 348016 318801
rect 363328 318792 363380 318844
rect 434352 318792 434404 318844
rect 434444 318792 434496 318844
rect 444104 318792 444156 318844
rect 444196 318792 444248 318844
rect 251456 318724 251508 318776
rect 262680 318767 262732 318776
rect 262680 318733 262689 318767
rect 262689 318733 262723 318767
rect 262723 318733 262732 318767
rect 262680 318724 262732 318733
rect 292856 318767 292908 318776
rect 292856 318733 292865 318767
rect 292865 318733 292899 318767
rect 292899 318733 292908 318767
rect 292856 318724 292908 318733
rect 298468 318724 298520 318776
rect 298560 318724 298612 318776
rect 316316 318724 316368 318776
rect 327448 318767 327500 318776
rect 327448 318733 327457 318767
rect 327457 318733 327491 318767
rect 327491 318733 327500 318767
rect 327448 318724 327500 318733
rect 328552 318724 328604 318776
rect 328736 318724 328788 318776
rect 342536 318767 342588 318776
rect 342536 318733 342545 318767
rect 342545 318733 342579 318767
rect 342579 318733 342588 318767
rect 342536 318724 342588 318733
rect 345204 318767 345256 318776
rect 345204 318733 345213 318767
rect 345213 318733 345247 318767
rect 345247 318733 345256 318767
rect 345204 318724 345256 318733
rect 324596 318656 324648 318708
rect 324780 318656 324832 318708
rect 234896 317432 234948 317484
rect 287336 317407 287388 317416
rect 287336 317373 287345 317407
rect 287345 317373 287379 317407
rect 287379 317373 287388 317407
rect 287336 317364 287388 317373
rect 298468 317407 298520 317416
rect 298468 317373 298477 317407
rect 298477 317373 298511 317407
rect 298511 317373 298520 317407
rect 298468 317364 298520 317373
rect 435364 316684 435416 316736
rect 435548 316684 435600 316736
rect 249984 316072 250036 316124
rect 250168 316072 250220 316124
rect 250168 315936 250220 315988
rect 290096 315911 290148 315920
rect 290096 315877 290105 315911
rect 290105 315877 290139 315911
rect 290139 315877 290148 315911
rect 290096 315868 290148 315877
rect 229468 313896 229520 313948
rect 229652 313896 229704 313948
rect 305368 312740 305420 312792
rect 305644 312740 305696 312792
rect 262680 312171 262732 312180
rect 262680 312137 262689 312171
rect 262689 312137 262723 312171
rect 262723 312137 262732 312171
rect 262680 312128 262732 312137
rect 248880 311924 248932 311976
rect 444104 311924 444156 311976
rect 444196 311924 444248 311976
rect 328644 311856 328696 311908
rect 287336 311831 287388 311840
rect 287336 311797 287345 311831
rect 287345 311797 287379 311831
rect 287379 311797 287388 311831
rect 287336 311788 287388 311797
rect 328644 311652 328696 311704
rect 238852 309748 238904 309800
rect 238852 309612 238904 309664
rect 347964 309272 348016 309324
rect 266912 309136 266964 309188
rect 267004 309136 267056 309188
rect 291476 309136 291528 309188
rect 291568 309136 291620 309188
rect 292856 309179 292908 309188
rect 292856 309145 292865 309179
rect 292865 309145 292899 309179
rect 292899 309145 292908 309179
rect 292856 309136 292908 309145
rect 327448 309179 327500 309188
rect 327448 309145 327457 309179
rect 327457 309145 327491 309179
rect 327491 309145 327500 309179
rect 327448 309136 327500 309145
rect 342536 309179 342588 309188
rect 342536 309145 342545 309179
rect 342545 309145 342579 309179
rect 342579 309145 342588 309179
rect 342536 309136 342588 309145
rect 345296 309136 345348 309188
rect 347964 309136 348016 309188
rect 362960 309136 363012 309188
rect 363328 309136 363380 309188
rect 229468 309068 229520 309120
rect 229652 309068 229704 309120
rect 235080 309111 235132 309120
rect 235080 309077 235089 309111
rect 235089 309077 235123 309111
rect 235123 309077 235132 309111
rect 235080 309068 235132 309077
rect 308036 309068 308088 309120
rect 308220 309068 308272 309120
rect 434536 309068 434588 309120
rect 267004 309043 267056 309052
rect 267004 309009 267013 309043
rect 267013 309009 267047 309043
rect 267047 309009 267056 309043
rect 267004 309000 267056 309009
rect 347964 309043 348016 309052
rect 347964 309009 347973 309043
rect 347973 309009 348007 309043
rect 348007 309009 348016 309043
rect 347964 309000 348016 309009
rect 290280 307776 290332 307828
rect 298468 307819 298520 307828
rect 298468 307785 298477 307819
rect 298477 307785 298511 307819
rect 298511 307785 298520 307819
rect 298468 307776 298520 307785
rect 234896 307751 234948 307760
rect 234896 307717 234905 307751
rect 234905 307717 234939 307751
rect 234939 307717 234948 307751
rect 234896 307708 234948 307717
rect 305552 307708 305604 307760
rect 316316 307751 316368 307760
rect 316316 307717 316325 307751
rect 316325 307717 316359 307751
rect 316359 307717 316368 307751
rect 316316 307708 316368 307717
rect 342444 307751 342496 307760
rect 342444 307717 342453 307751
rect 342453 307717 342487 307751
rect 342487 307717 342496 307751
rect 342444 307708 342496 307717
rect 254124 306416 254176 306468
rect 254308 306416 254360 306468
rect 313464 306348 313516 306400
rect 313556 306348 313608 306400
rect 288716 302268 288768 302320
rect 233332 302200 233384 302252
rect 233516 302200 233568 302252
rect 280436 302200 280488 302252
rect 280620 302200 280672 302252
rect 435364 302200 435416 302252
rect 435548 302200 435600 302252
rect 444012 302200 444064 302252
rect 444196 302200 444248 302252
rect 288716 302132 288768 302184
rect 362960 302064 363012 302116
rect 363236 302064 363288 302116
rect 229468 299548 229520 299600
rect 244188 299548 244240 299600
rect 347964 299591 348016 299600
rect 347964 299557 347973 299591
rect 347973 299557 348007 299591
rect 348007 299557 348016 299591
rect 347964 299548 348016 299557
rect 235080 299523 235132 299532
rect 235080 299489 235089 299523
rect 235089 299489 235123 299523
rect 235123 299489 235132 299523
rect 235080 299480 235132 299489
rect 244280 299480 244332 299532
rect 248788 299523 248840 299532
rect 248788 299489 248797 299523
rect 248797 299489 248831 299523
rect 248831 299489 248840 299523
rect 248788 299480 248840 299489
rect 250076 299523 250128 299532
rect 250076 299489 250085 299523
rect 250085 299489 250119 299523
rect 250119 299489 250128 299523
rect 250076 299480 250128 299489
rect 267280 299480 267332 299532
rect 290096 299480 290148 299532
rect 290280 299480 290332 299532
rect 434260 299523 434312 299532
rect 434260 299489 434269 299523
rect 434269 299489 434303 299523
rect 434303 299489 434312 299523
rect 434260 299480 434312 299489
rect 262680 299412 262732 299464
rect 287336 299455 287388 299464
rect 287336 299421 287345 299455
rect 287345 299421 287379 299455
rect 287379 299421 287388 299455
rect 287336 299412 287388 299421
rect 291476 299412 291528 299464
rect 291568 299412 291620 299464
rect 298560 299412 298612 299464
rect 324688 299412 324740 299464
rect 327264 299412 327316 299464
rect 327448 299412 327500 299464
rect 347964 299412 348016 299464
rect 348056 299412 348108 299464
rect 577504 299412 577556 299464
rect 579896 299412 579948 299464
rect 229284 298163 229336 298172
rect 229284 298129 229293 298163
rect 229293 298129 229327 298163
rect 229327 298129 229336 298163
rect 229284 298120 229336 298129
rect 234896 298163 234948 298172
rect 234896 298129 234905 298163
rect 234905 298129 234939 298163
rect 234939 298129 234948 298163
rect 234896 298120 234948 298129
rect 305460 298163 305512 298172
rect 305460 298129 305469 298163
rect 305469 298129 305503 298163
rect 305503 298129 305512 298163
rect 305460 298120 305512 298129
rect 310888 298120 310940 298172
rect 316316 298163 316368 298172
rect 316316 298129 316325 298163
rect 316325 298129 316359 298163
rect 316359 298129 316368 298163
rect 316316 298120 316368 298129
rect 342536 298120 342588 298172
rect 235080 298095 235132 298104
rect 235080 298061 235089 298095
rect 235089 298061 235123 298095
rect 235123 298061 235132 298095
rect 235080 298052 235132 298061
rect 239036 298052 239088 298104
rect 239128 298052 239180 298104
rect 240416 298095 240468 298104
rect 240416 298061 240425 298095
rect 240425 298061 240459 298095
rect 240459 298061 240468 298095
rect 240416 298052 240468 298061
rect 241888 298095 241940 298104
rect 241888 298061 241897 298095
rect 241897 298061 241931 298095
rect 241931 298061 241940 298095
rect 241888 298052 241940 298061
rect 291476 298095 291528 298104
rect 291476 298061 291485 298095
rect 291485 298061 291519 298095
rect 291519 298061 291528 298095
rect 291476 298052 291528 298061
rect 308128 298052 308180 298104
rect 308220 298052 308272 298104
rect 327264 298095 327316 298104
rect 327264 298061 327273 298095
rect 327273 298061 327307 298095
rect 327307 298061 327316 298095
rect 327264 298052 327316 298061
rect 435364 297372 435416 297424
rect 435548 297372 435600 297424
rect 253940 296692 253992 296744
rect 254216 296692 254268 296744
rect 310796 296735 310848 296744
rect 310796 296701 310805 296735
rect 310805 296701 310839 296735
rect 310839 296701 310848 296735
rect 310796 296692 310848 296701
rect 310796 295740 310848 295792
rect 310980 295740 311032 295792
rect 2780 295196 2832 295248
rect 5264 295196 5316 295248
rect 326068 294652 326120 294704
rect 254216 292612 254268 292664
rect 342536 292612 342588 292664
rect 267004 292544 267056 292596
rect 267280 292544 267332 292596
rect 328552 292544 328604 292596
rect 328736 292544 328788 292596
rect 254216 292476 254268 292528
rect 342536 292476 342588 292528
rect 229376 292408 229428 292460
rect 229560 292408 229612 292460
rect 262588 289935 262640 289944
rect 262588 289901 262597 289935
rect 262597 289901 262631 289935
rect 262631 289901 262640 289935
rect 262588 289892 262640 289901
rect 324596 289935 324648 289944
rect 324596 289901 324605 289935
rect 324605 289901 324639 289935
rect 324639 289901 324648 289935
rect 324596 289892 324648 289901
rect 261208 289824 261260 289876
rect 261300 289824 261352 289876
rect 287336 289867 287388 289876
rect 287336 289833 287345 289867
rect 287345 289833 287379 289867
rect 287379 289833 287388 289867
rect 287336 289824 287388 289833
rect 288716 289824 288768 289876
rect 288992 289824 289044 289876
rect 298468 289867 298520 289876
rect 298468 289833 298477 289867
rect 298477 289833 298511 289867
rect 298511 289833 298520 289867
rect 298468 289824 298520 289833
rect 305460 289824 305512 289876
rect 325976 289867 326028 289876
rect 325976 289833 325985 289867
rect 325985 289833 326019 289867
rect 326019 289833 326028 289867
rect 325976 289824 326028 289833
rect 267004 289756 267056 289808
rect 267280 289756 267332 289808
rect 324596 289756 324648 289808
rect 345204 289799 345256 289808
rect 345204 289765 345213 289799
rect 345213 289765 345247 289799
rect 345247 289765 345256 289799
rect 345204 289756 345256 289765
rect 347780 289756 347832 289808
rect 347964 289756 348016 289808
rect 434352 289756 434404 289808
rect 288716 289731 288768 289740
rect 288716 289697 288725 289731
rect 288725 289697 288759 289731
rect 288759 289697 288768 289731
rect 288716 289688 288768 289697
rect 305460 289688 305512 289740
rect 324780 289688 324832 289740
rect 316316 288464 316368 288516
rect 240416 288439 240468 288448
rect 240416 288405 240425 288439
rect 240425 288405 240459 288439
rect 240459 288405 240468 288439
rect 240416 288396 240468 288405
rect 241888 288439 241940 288448
rect 241888 288405 241897 288439
rect 241897 288405 241931 288439
rect 241931 288405 241940 288439
rect 241888 288396 241940 288405
rect 291476 288439 291528 288448
rect 291476 288405 291485 288439
rect 291485 288405 291519 288439
rect 291519 288405 291528 288439
rect 291476 288396 291528 288405
rect 327540 288396 327592 288448
rect 262588 288328 262640 288380
rect 316224 287079 316276 287088
rect 316224 287045 316233 287079
rect 316233 287045 316267 287079
rect 316267 287045 316276 287079
rect 316224 287036 316276 287045
rect 229376 282956 229428 283008
rect 233332 282888 233384 282940
rect 233516 282888 233568 282940
rect 280436 282888 280488 282940
rect 280620 282888 280672 282940
rect 298468 282888 298520 282940
rect 435364 282888 435416 282940
rect 435548 282888 435600 282940
rect 444012 282888 444064 282940
rect 444196 282888 444248 282940
rect 288716 282863 288768 282872
rect 288716 282829 288725 282863
rect 288725 282829 288759 282863
rect 288759 282829 288768 282863
rect 288716 282820 288768 282829
rect 229376 282752 229428 282804
rect 298560 282752 298612 282804
rect 345204 280279 345256 280288
rect 345204 280245 345213 280279
rect 345213 280245 345247 280279
rect 345247 280245 345256 280279
rect 345204 280236 345256 280245
rect 235080 280211 235132 280220
rect 235080 280177 235089 280211
rect 235089 280177 235123 280211
rect 235123 280177 235132 280211
rect 235080 280168 235132 280177
rect 434260 280211 434312 280220
rect 434260 280177 434269 280211
rect 434269 280177 434303 280211
rect 434303 280177 434312 280211
rect 434260 280168 434312 280177
rect 3148 280100 3200 280152
rect 6276 280100 6328 280152
rect 229376 280143 229428 280152
rect 229376 280109 229385 280143
rect 229385 280109 229419 280143
rect 229419 280109 229428 280143
rect 229376 280100 229428 280109
rect 254216 280143 254268 280152
rect 254216 280109 254225 280143
rect 254225 280109 254259 280143
rect 254259 280109 254268 280143
rect 254216 280100 254268 280109
rect 287336 280143 287388 280152
rect 287336 280109 287345 280143
rect 287345 280109 287379 280143
rect 287379 280109 287388 280143
rect 287336 280100 287388 280109
rect 290096 280143 290148 280152
rect 290096 280109 290105 280143
rect 290105 280109 290139 280143
rect 290139 280109 290148 280143
rect 290096 280100 290148 280109
rect 291476 280100 291528 280152
rect 291568 280100 291620 280152
rect 298560 280100 298612 280152
rect 305460 280100 305512 280152
rect 324504 280100 324556 280152
rect 324780 280100 324832 280152
rect 327540 280100 327592 280152
rect 342536 280143 342588 280152
rect 342536 280109 342545 280143
rect 342545 280109 342579 280143
rect 342579 280109 342588 280143
rect 342536 280100 342588 280109
rect 347964 280100 348016 280152
rect 348056 280100 348108 280152
rect 363144 280143 363196 280152
rect 363144 280109 363153 280143
rect 363153 280109 363187 280143
rect 363187 280109 363196 280143
rect 363144 280100 363196 280109
rect 305276 280032 305328 280084
rect 327356 280032 327408 280084
rect 239128 278740 239180 278792
rect 239312 278740 239364 278792
rect 251180 278740 251232 278792
rect 251456 278740 251508 278792
rect 255504 278740 255556 278792
rect 255872 278740 255924 278792
rect 262404 278876 262456 278928
rect 262496 278851 262548 278860
rect 262496 278817 262505 278851
rect 262505 278817 262539 278851
rect 262539 278817 262548 278851
rect 262496 278808 262548 278817
rect 262404 278740 262456 278792
rect 307944 278740 307996 278792
rect 308220 278740 308272 278792
rect 316224 278740 316276 278792
rect 316316 278740 316368 278792
rect 235080 278715 235132 278724
rect 235080 278681 235089 278715
rect 235089 278681 235123 278715
rect 235123 278681 235132 278715
rect 235080 278672 235132 278681
rect 262496 278715 262548 278724
rect 262496 278681 262505 278715
rect 262505 278681 262539 278715
rect 262539 278681 262548 278715
rect 262496 278672 262548 278681
rect 324504 278715 324556 278724
rect 324504 278681 324513 278715
rect 324513 278681 324547 278715
rect 324547 278681 324556 278715
rect 324504 278672 324556 278681
rect 435364 278060 435416 278112
rect 435548 278060 435600 278112
rect 310704 277380 310756 277432
rect 310796 277380 310848 277432
rect 239128 274048 239180 274100
rect 251456 273887 251508 273896
rect 251456 273853 251465 273887
rect 251465 273853 251499 273887
rect 251499 273853 251508 273887
rect 251456 273844 251508 273853
rect 310704 273411 310756 273420
rect 310704 273377 310713 273411
rect 310713 273377 310747 273411
rect 310747 273377 310756 273411
rect 310704 273368 310756 273377
rect 261208 273164 261260 273216
rect 299848 273164 299900 273216
rect 309416 273207 309468 273216
rect 309416 273173 309425 273207
rect 309425 273173 309459 273207
rect 309459 273173 309468 273207
rect 309416 273164 309468 273173
rect 325976 273164 326028 273216
rect 229376 273139 229428 273148
rect 229376 273105 229385 273139
rect 229385 273105 229419 273139
rect 229419 273105 229428 273139
rect 229376 273096 229428 273105
rect 261208 273028 261260 273080
rect 299848 273028 299900 273080
rect 325976 273028 326028 273080
rect 290096 273003 290148 273012
rect 290096 272969 290105 273003
rect 290105 272969 290139 273003
rect 290139 272969 290148 273003
rect 290096 272960 290148 272969
rect 298468 270623 298520 270632
rect 298468 270589 298477 270623
rect 298477 270589 298511 270623
rect 298511 270589 298520 270623
rect 298468 270580 298520 270589
rect 254216 270555 254268 270564
rect 254216 270521 254225 270555
rect 254225 270521 254259 270555
rect 254259 270521 254268 270555
rect 254216 270512 254268 270521
rect 255596 270512 255648 270564
rect 255872 270512 255924 270564
rect 287336 270555 287388 270564
rect 287336 270521 287345 270555
rect 287345 270521 287379 270555
rect 287379 270521 287388 270555
rect 287336 270512 287388 270521
rect 288624 270512 288676 270564
rect 288716 270512 288768 270564
rect 342536 270555 342588 270564
rect 342536 270521 342545 270555
rect 342545 270521 342579 270555
rect 342579 270521 342588 270555
rect 342536 270512 342588 270521
rect 363236 270512 363288 270564
rect 229376 270487 229428 270496
rect 229376 270453 229385 270487
rect 229385 270453 229419 270487
rect 229419 270453 229428 270487
rect 229376 270444 229428 270453
rect 244280 270487 244332 270496
rect 244280 270453 244289 270487
rect 244289 270453 244323 270487
rect 244323 270453 244332 270487
rect 244280 270444 244332 270453
rect 245936 270487 245988 270496
rect 245936 270453 245945 270487
rect 245945 270453 245979 270487
rect 245979 270453 245988 270487
rect 245936 270444 245988 270453
rect 307944 270487 307996 270496
rect 307944 270453 307953 270487
rect 307953 270453 307987 270487
rect 307987 270453 307996 270487
rect 307944 270444 307996 270453
rect 345204 270487 345256 270496
rect 345204 270453 345213 270487
rect 345213 270453 345247 270487
rect 345247 270453 345256 270487
rect 345204 270444 345256 270453
rect 347964 270487 348016 270496
rect 347964 270453 347973 270487
rect 347973 270453 348007 270487
rect 348007 270453 348016 270487
rect 347964 270444 348016 270453
rect 434352 270444 434404 270496
rect 255596 270419 255648 270428
rect 255596 270385 255605 270419
rect 255605 270385 255639 270419
rect 255639 270385 255648 270419
rect 255596 270376 255648 270385
rect 288716 270419 288768 270428
rect 288716 270385 288725 270419
rect 288725 270385 288759 270419
rect 288759 270385 288768 270419
rect 288716 270376 288768 270385
rect 240232 269084 240284 269136
rect 240416 269084 240468 269136
rect 241888 269084 241940 269136
rect 242072 269084 242124 269136
rect 291476 269084 291528 269136
rect 291660 269084 291712 269136
rect 310796 267792 310848 267844
rect 239312 267767 239364 267776
rect 239312 267733 239321 267767
rect 239321 267733 239355 267767
rect 239355 267733 239364 267767
rect 309416 267767 309468 267776
rect 239312 267724 239364 267733
rect 309416 267733 309425 267767
rect 309425 267733 309459 267767
rect 309459 267733 309468 267767
rect 309416 267724 309468 267733
rect 310796 263644 310848 263696
rect 233332 263576 233384 263628
rect 233516 263576 233568 263628
rect 280436 263576 280488 263628
rect 280620 263576 280672 263628
rect 291476 263576 291528 263628
rect 298468 263576 298520 263628
rect 288716 263551 288768 263560
rect 288716 263517 288725 263551
rect 288725 263517 288759 263551
rect 288759 263517 288768 263551
rect 288716 263508 288768 263517
rect 229376 263483 229428 263492
rect 229376 263449 229385 263483
rect 229385 263449 229419 263483
rect 229419 263449 229428 263483
rect 229376 263440 229428 263449
rect 262680 263440 262732 263492
rect 291568 263440 291620 263492
rect 435364 263576 435416 263628
rect 435548 263576 435600 263628
rect 444012 263576 444064 263628
rect 444196 263576 444248 263628
rect 310796 263508 310848 263560
rect 298560 263440 298612 263492
rect 324688 263440 324740 263492
rect 345204 260967 345256 260976
rect 345204 260933 345213 260967
rect 345213 260933 345247 260967
rect 345247 260933 345256 260967
rect 345204 260924 345256 260933
rect 347964 260967 348016 260976
rect 347964 260933 347973 260967
rect 347973 260933 348007 260967
rect 348007 260933 348016 260967
rect 347964 260924 348016 260933
rect 235080 260899 235132 260908
rect 235080 260865 235089 260899
rect 235089 260865 235123 260899
rect 235123 260865 235132 260899
rect 235080 260856 235132 260865
rect 244280 260899 244332 260908
rect 244280 260865 244289 260899
rect 244289 260865 244323 260899
rect 244323 260865 244332 260899
rect 244280 260856 244332 260865
rect 245936 260899 245988 260908
rect 245936 260865 245945 260899
rect 245945 260865 245979 260899
rect 245979 260865 245988 260899
rect 245936 260856 245988 260865
rect 251456 260899 251508 260908
rect 251456 260865 251465 260899
rect 251465 260865 251499 260899
rect 251499 260865 251508 260899
rect 251456 260856 251508 260865
rect 255688 260856 255740 260908
rect 434260 260899 434312 260908
rect 434260 260865 434269 260899
rect 434269 260865 434303 260899
rect 434303 260865 434312 260899
rect 434260 260856 434312 260865
rect 229376 260831 229428 260840
rect 229376 260797 229385 260831
rect 229385 260797 229419 260831
rect 229419 260797 229428 260831
rect 229376 260788 229428 260797
rect 254216 260831 254268 260840
rect 254216 260797 254225 260831
rect 254225 260797 254259 260831
rect 254259 260797 254268 260831
rect 254216 260788 254268 260797
rect 262680 260788 262732 260840
rect 287336 260831 287388 260840
rect 287336 260797 287345 260831
rect 287345 260797 287379 260831
rect 287379 260797 287388 260831
rect 287336 260788 287388 260797
rect 290096 260831 290148 260840
rect 290096 260797 290105 260831
rect 290105 260797 290139 260831
rect 290139 260797 290148 260831
rect 290096 260788 290148 260797
rect 291568 260788 291620 260840
rect 298560 260788 298612 260840
rect 324688 260788 324740 260840
rect 342536 260831 342588 260840
rect 342536 260797 342545 260831
rect 342545 260797 342579 260831
rect 342579 260797 342588 260831
rect 342536 260788 342588 260797
rect 347964 260788 348016 260840
rect 363144 260831 363196 260840
rect 363144 260797 363153 260831
rect 363153 260797 363187 260831
rect 363187 260797 363196 260831
rect 363144 260788 363196 260797
rect 435272 260831 435324 260840
rect 435272 260797 435281 260831
rect 435281 260797 435315 260831
rect 435315 260797 435324 260831
rect 435272 260788 435324 260797
rect 255688 260720 255740 260772
rect 348056 260720 348108 260772
rect 234620 259428 234672 259480
rect 234896 259428 234948 259480
rect 239128 259428 239180 259480
rect 239312 259428 239364 259480
rect 267188 259428 267240 259480
rect 267280 259428 267332 259480
rect 235080 259403 235132 259412
rect 235080 259369 235089 259403
rect 235089 259369 235123 259403
rect 235123 259369 235132 259403
rect 235080 259360 235132 259369
rect 251456 259403 251508 259412
rect 251456 259369 251465 259403
rect 251465 259369 251499 259403
rect 251499 259369 251508 259403
rect 251456 259360 251508 259369
rect 307944 258111 307996 258120
rect 307944 258077 307953 258111
rect 307953 258077 307987 258111
rect 307987 258077 307996 258111
rect 307944 258068 307996 258077
rect 310888 256640 310940 256692
rect 261208 253852 261260 253904
rect 299848 253852 299900 253904
rect 325976 253852 326028 253904
rect 229376 253827 229428 253836
rect 229376 253793 229385 253827
rect 229385 253793 229419 253827
rect 229419 253793 229428 253827
rect 229376 253784 229428 253793
rect 261208 253716 261260 253768
rect 299848 253716 299900 253768
rect 325976 253716 326028 253768
rect 290096 252875 290148 252884
rect 290096 252841 290105 252875
rect 290105 252841 290139 252875
rect 290139 252841 290148 252875
rect 290096 252832 290148 252841
rect 291476 251311 291528 251320
rect 291476 251277 291485 251311
rect 291485 251277 291519 251311
rect 291519 251277 291528 251311
rect 291476 251268 291528 251277
rect 298468 251311 298520 251320
rect 298468 251277 298477 251311
rect 298477 251277 298511 251311
rect 298511 251277 298520 251311
rect 298468 251268 298520 251277
rect 435272 251311 435324 251320
rect 435272 251277 435281 251311
rect 435281 251277 435315 251311
rect 435315 251277 435324 251311
rect 435272 251268 435324 251277
rect 234896 251200 234948 251252
rect 254216 251243 254268 251252
rect 254216 251209 254225 251243
rect 254225 251209 254259 251243
rect 254259 251209 254268 251243
rect 254216 251200 254268 251209
rect 255596 251243 255648 251252
rect 255596 251209 255605 251243
rect 255605 251209 255639 251243
rect 255639 251209 255648 251243
rect 255596 251200 255648 251209
rect 262588 251243 262640 251252
rect 262588 251209 262597 251243
rect 262597 251209 262631 251243
rect 262631 251209 262640 251243
rect 262588 251200 262640 251209
rect 287336 251243 287388 251252
rect 287336 251209 287345 251243
rect 287345 251209 287379 251243
rect 287379 251209 287388 251243
rect 287336 251200 287388 251209
rect 288624 251200 288676 251252
rect 288716 251200 288768 251252
rect 324596 251243 324648 251252
rect 324596 251209 324605 251243
rect 324605 251209 324639 251243
rect 324639 251209 324648 251243
rect 324596 251200 324648 251209
rect 342536 251243 342588 251252
rect 342536 251209 342545 251243
rect 342545 251209 342579 251243
rect 342579 251209 342588 251243
rect 342536 251200 342588 251209
rect 363236 251200 363288 251252
rect 244280 251175 244332 251184
rect 244280 251141 244289 251175
rect 244289 251141 244323 251175
rect 244323 251141 244332 251175
rect 244280 251132 244332 251141
rect 245936 251175 245988 251184
rect 245936 251141 245945 251175
rect 245945 251141 245979 251175
rect 245979 251141 245988 251175
rect 245936 251132 245988 251141
rect 291476 251175 291528 251184
rect 291476 251141 291485 251175
rect 291485 251141 291519 251175
rect 291519 251141 291528 251175
rect 291476 251132 291528 251141
rect 298468 251175 298520 251184
rect 298468 251141 298477 251175
rect 298477 251141 298511 251175
rect 298511 251141 298520 251175
rect 298468 251132 298520 251141
rect 305276 251132 305328 251184
rect 307944 251175 307996 251184
rect 307944 251141 307953 251175
rect 307953 251141 307987 251175
rect 307987 251141 307996 251175
rect 307944 251132 307996 251141
rect 327356 251132 327408 251184
rect 345204 251175 345256 251184
rect 345204 251141 345213 251175
rect 345213 251141 345247 251175
rect 345247 251141 345256 251175
rect 345204 251132 345256 251141
rect 347964 251175 348016 251184
rect 347964 251141 347973 251175
rect 347973 251141 348007 251175
rect 348007 251141 348016 251175
rect 347964 251132 348016 251141
rect 434352 251132 434404 251184
rect 435180 251132 435232 251184
rect 234988 251064 235040 251116
rect 251548 251064 251600 251116
rect 239220 249840 239272 249892
rect 240232 249772 240284 249824
rect 240416 249772 240468 249824
rect 241888 249772 241940 249824
rect 242072 249772 242124 249824
rect 267004 249772 267056 249824
rect 267280 249772 267332 249824
rect 229376 244332 229428 244384
rect 233332 244264 233384 244316
rect 233516 244264 233568 244316
rect 288716 244264 288768 244316
rect 444012 244264 444064 244316
rect 444196 244264 444248 244316
rect 229284 244196 229336 244248
rect 308036 244196 308088 244248
rect 288808 244128 288860 244180
rect 327264 242675 327316 242684
rect 327264 242641 327273 242675
rect 327273 242641 327307 242675
rect 327307 242641 327316 242675
rect 327264 242632 327316 242641
rect 234896 241476 234948 241528
rect 234988 241476 235040 241528
rect 235080 241519 235132 241528
rect 235080 241485 235089 241519
rect 235089 241485 235123 241519
rect 235123 241485 235132 241519
rect 244280 241519 244332 241528
rect 235080 241476 235132 241485
rect 244280 241485 244289 241519
rect 244289 241485 244323 241519
rect 244323 241485 244332 241519
rect 244280 241476 244332 241485
rect 245936 241519 245988 241528
rect 245936 241485 245945 241519
rect 245945 241485 245979 241519
rect 245979 241485 245988 241519
rect 245936 241476 245988 241485
rect 251456 241519 251508 241528
rect 251456 241485 251465 241519
rect 251465 241485 251499 241519
rect 251499 241485 251508 241519
rect 251456 241476 251508 241485
rect 255780 241476 255832 241528
rect 255872 241476 255924 241528
rect 262772 241476 262824 241528
rect 262864 241476 262916 241528
rect 267004 241476 267056 241528
rect 291568 241476 291620 241528
rect 298560 241476 298612 241528
rect 305184 241519 305236 241528
rect 305184 241485 305193 241519
rect 305193 241485 305227 241519
rect 305227 241485 305236 241519
rect 305184 241476 305236 241485
rect 324780 241476 324832 241528
rect 324872 241476 324924 241528
rect 345204 241519 345256 241528
rect 345204 241485 345213 241519
rect 345213 241485 345247 241519
rect 345247 241485 345256 241519
rect 345204 241476 345256 241485
rect 347964 241519 348016 241528
rect 347964 241485 347973 241519
rect 347973 241485 348007 241519
rect 348007 241485 348016 241519
rect 347964 241476 348016 241485
rect 434260 241519 434312 241528
rect 434260 241485 434269 241519
rect 434269 241485 434303 241519
rect 434303 241485 434312 241519
rect 434260 241476 434312 241485
rect 435088 241519 435140 241528
rect 435088 241485 435097 241519
rect 435097 241485 435131 241519
rect 435131 241485 435140 241519
rect 435088 241476 435140 241485
rect 267004 241340 267056 241392
rect 239128 240159 239180 240168
rect 239128 240125 239137 240159
rect 239137 240125 239171 240159
rect 239171 240125 239180 240159
rect 239128 240116 239180 240125
rect 251456 240159 251508 240168
rect 251456 240125 251465 240159
rect 251465 240125 251499 240159
rect 251499 240125 251508 240159
rect 251456 240116 251508 240125
rect 234896 240091 234948 240100
rect 234896 240057 234905 240091
rect 234905 240057 234939 240091
rect 234939 240057 234948 240091
rect 234896 240048 234948 240057
rect 288716 240091 288768 240100
rect 288716 240057 288725 240091
rect 288725 240057 288759 240091
rect 288759 240057 288768 240091
rect 288716 240048 288768 240057
rect 327264 240048 327316 240100
rect 327356 240048 327408 240100
rect 251456 240023 251508 240032
rect 251456 239989 251465 240023
rect 251465 239989 251499 240023
rect 251499 239989 251508 240023
rect 251456 239980 251508 239989
rect 310796 240023 310848 240032
rect 310796 239989 310805 240023
rect 310805 239989 310839 240023
rect 310839 239989 310848 240023
rect 310796 239980 310848 239989
rect 310704 238688 310756 238740
rect 310796 238688 310848 238740
rect 280620 234676 280672 234728
rect 434260 234608 434312 234660
rect 435088 234608 435140 234660
rect 261208 234540 261260 234592
rect 280528 234540 280580 234592
rect 287336 234540 287388 234592
rect 299848 234540 299900 234592
rect 325976 234540 326028 234592
rect 434352 234472 434404 234524
rect 435180 234472 435232 234524
rect 261208 234404 261260 234456
rect 287336 234404 287388 234456
rect 299848 234404 299900 234456
rect 325976 234404 326028 234456
rect 308036 231956 308088 232008
rect 345388 231888 345440 231940
rect 254216 231820 254268 231872
rect 254400 231820 254452 231872
rect 262588 231820 262640 231872
rect 262864 231820 262916 231872
rect 288808 231820 288860 231872
rect 298560 231820 298612 231872
rect 305184 231820 305236 231872
rect 305276 231820 305328 231872
rect 308036 231820 308088 231872
rect 324596 231820 324648 231872
rect 324872 231820 324924 231872
rect 342352 231820 342404 231872
rect 342536 231820 342588 231872
rect 345296 231820 345348 231872
rect 362960 231820 363012 231872
rect 363236 231820 363288 231872
rect 244464 231752 244516 231804
rect 244556 231752 244608 231804
rect 298560 231684 298612 231736
rect 229376 230460 229428 230512
rect 229560 230460 229612 230512
rect 234896 230503 234948 230512
rect 234896 230469 234905 230503
rect 234905 230469 234939 230503
rect 234939 230469 234948 230503
rect 234896 230460 234948 230469
rect 235080 230460 235132 230512
rect 235264 230460 235316 230512
rect 240232 230460 240284 230512
rect 240416 230460 240468 230512
rect 241888 230460 241940 230512
rect 242072 230460 242124 230512
rect 251456 230503 251508 230512
rect 251456 230469 251465 230503
rect 251465 230469 251499 230503
rect 251499 230469 251508 230503
rect 251456 230460 251508 230469
rect 255780 230460 255832 230512
rect 255872 230460 255924 230512
rect 266820 230460 266872 230512
rect 267004 230460 267056 230512
rect 291568 230460 291620 230512
rect 291660 230460 291712 230512
rect 298560 229032 298612 229084
rect 298652 229032 298704 229084
rect 229376 225020 229428 225072
rect 233332 224952 233384 225004
rect 233516 224952 233568 225004
rect 288808 224952 288860 225004
rect 229284 224884 229336 224936
rect 434352 225020 434404 225072
rect 435088 224995 435140 225004
rect 435088 224961 435097 224995
rect 435097 224961 435131 224995
rect 435131 224961 435140 224995
rect 435088 224952 435140 224961
rect 444012 224952 444064 225004
rect 444196 224952 444248 225004
rect 434260 224884 434312 224936
rect 288808 224816 288860 224868
rect 251180 224204 251232 224256
rect 251456 224204 251508 224256
rect 235080 222300 235132 222352
rect 235080 222164 235132 222216
rect 244188 222164 244240 222216
rect 244280 222164 244332 222216
rect 245752 222164 245804 222216
rect 245936 222164 245988 222216
rect 262496 222164 262548 222216
rect 262864 222164 262916 222216
rect 345204 222164 345256 222216
rect 345296 222164 345348 222216
rect 347964 222164 348016 222216
rect 348148 222164 348200 222216
rect 435088 222207 435140 222216
rect 435088 222173 435097 222207
rect 435097 222173 435131 222207
rect 435131 222173 435140 222207
rect 435088 222164 435140 222173
rect 291384 220872 291436 220924
rect 291752 220872 291804 220924
rect 239128 220804 239180 220856
rect 239220 220804 239272 220856
rect 266912 220804 266964 220856
rect 267004 220804 267056 220856
rect 316224 220804 316276 220856
rect 316316 220804 316368 220856
rect 327356 220804 327408 220856
rect 327540 220804 327592 220856
rect 229284 220779 229336 220788
rect 229284 220745 229293 220779
rect 229293 220745 229327 220779
rect 229327 220745 229336 220779
rect 229284 220736 229336 220745
rect 235080 220779 235132 220788
rect 235080 220745 235089 220779
rect 235089 220745 235123 220779
rect 235123 220745 235132 220779
rect 235080 220736 235132 220745
rect 291384 220779 291436 220788
rect 291384 220745 291393 220779
rect 291393 220745 291427 220779
rect 291427 220745 291436 220779
rect 291384 220736 291436 220745
rect 434260 220779 434312 220788
rect 434260 220745 434269 220779
rect 434269 220745 434303 220779
rect 434303 220745 434312 220779
rect 434260 220736 434312 220745
rect 310888 219419 310940 219428
rect 310888 219385 310897 219419
rect 310897 219385 310931 219419
rect 310931 219385 310940 219419
rect 310888 219376 310940 219385
rect 308036 217447 308088 217456
rect 308036 217413 308045 217447
rect 308045 217413 308079 217447
rect 308079 217413 308088 217447
rect 308036 217404 308088 217413
rect 261208 215976 261260 216028
rect 261392 215976 261444 216028
rect 327356 215364 327408 215416
rect 267004 215339 267056 215348
rect 267004 215305 267013 215339
rect 267013 215305 267047 215339
rect 267047 215305 267056 215339
rect 267004 215296 267056 215305
rect 288716 215339 288768 215348
rect 288716 215305 288725 215339
rect 288725 215305 288759 215339
rect 288759 215305 288768 215339
rect 288716 215296 288768 215305
rect 305368 215296 305420 215348
rect 435088 215296 435140 215348
rect 229284 215271 229336 215280
rect 229284 215237 229293 215271
rect 229293 215237 229327 215271
rect 229327 215237 229336 215271
rect 229284 215228 229336 215237
rect 273352 215228 273404 215280
rect 273536 215228 273588 215280
rect 299848 215228 299900 215280
rect 305276 215228 305328 215280
rect 325976 215228 326028 215280
rect 327356 215228 327408 215280
rect 434260 215271 434312 215280
rect 434260 215237 434269 215271
rect 434269 215237 434303 215271
rect 434303 215237 434312 215271
rect 434260 215228 434312 215237
rect 435180 215160 435232 215212
rect 299848 215092 299900 215144
rect 325976 215092 326028 215144
rect 310888 214591 310940 214600
rect 310888 214557 310897 214591
rect 310897 214557 310931 214591
rect 310931 214557 310940 214591
rect 310888 214548 310940 214557
rect 345388 212576 345440 212628
rect 254216 212508 254268 212560
rect 254400 212508 254452 212560
rect 262588 212508 262640 212560
rect 262864 212508 262916 212560
rect 267004 212551 267056 212560
rect 267004 212517 267013 212551
rect 267013 212517 267047 212551
rect 267047 212517 267056 212551
rect 267004 212508 267056 212517
rect 287336 212508 287388 212560
rect 287520 212508 287572 212560
rect 288808 212508 288860 212560
rect 308036 212551 308088 212560
rect 308036 212517 308045 212551
rect 308045 212517 308079 212551
rect 308079 212517 308088 212551
rect 308036 212508 308088 212517
rect 324596 212508 324648 212560
rect 324872 212508 324924 212560
rect 342352 212508 342404 212560
rect 342536 212508 342588 212560
rect 343824 212508 343876 212560
rect 345296 212508 345348 212560
rect 362960 212508 363012 212560
rect 363236 212508 363288 212560
rect 343732 212440 343784 212492
rect 239036 211216 239088 211268
rect 239128 211216 239180 211268
rect 235080 211191 235132 211200
rect 235080 211157 235089 211191
rect 235089 211157 235123 211191
rect 235123 211157 235132 211191
rect 235080 211148 235132 211157
rect 239128 211123 239180 211132
rect 239128 211089 239137 211123
rect 239137 211089 239171 211123
rect 239171 211089 239180 211123
rect 239128 211080 239180 211089
rect 267004 211123 267056 211132
rect 267004 211089 267013 211123
rect 267013 211089 267047 211123
rect 267047 211089 267056 211123
rect 267004 211080 267056 211089
rect 316316 211080 316368 211132
rect 316500 211080 316552 211132
rect 327356 211080 327408 211132
rect 327540 211080 327592 211132
rect 343732 211123 343784 211132
rect 343732 211089 343741 211123
rect 343741 211089 343775 211123
rect 343775 211089 343784 211123
rect 343732 211080 343784 211089
rect 251364 209720 251416 209772
rect 251732 209720 251784 209772
rect 2780 208156 2832 208208
rect 5172 208156 5224 208208
rect 233332 205640 233384 205692
rect 233516 205640 233568 205692
rect 288808 205683 288860 205692
rect 288808 205649 288817 205683
rect 288817 205649 288851 205683
rect 288851 205649 288860 205683
rect 288808 205640 288860 205649
rect 305276 205683 305328 205692
rect 305276 205649 305285 205683
rect 305285 205649 305319 205683
rect 305319 205649 305328 205683
rect 305276 205640 305328 205649
rect 444012 205640 444064 205692
rect 444196 205640 444248 205692
rect 308036 205504 308088 205556
rect 308220 205504 308272 205556
rect 238760 204552 238812 204604
rect 238944 204552 238996 204604
rect 255596 202920 255648 202972
rect 255688 202920 255740 202972
rect 291384 202963 291436 202972
rect 291384 202929 291393 202963
rect 291393 202929 291427 202963
rect 291427 202929 291436 202963
rect 291384 202920 291436 202929
rect 229284 202852 229336 202904
rect 229376 202852 229428 202904
rect 234804 202852 234856 202904
rect 234896 202852 234948 202904
rect 288808 202895 288860 202904
rect 288808 202861 288817 202895
rect 288817 202861 288851 202895
rect 288851 202861 288860 202895
rect 288808 202852 288860 202861
rect 305276 202895 305328 202904
rect 305276 202861 305285 202895
rect 305285 202861 305319 202895
rect 305319 202861 305328 202895
rect 305276 202852 305328 202861
rect 347964 202852 348016 202904
rect 348148 202852 348200 202904
rect 434352 202852 434404 202904
rect 434536 202852 434588 202904
rect 239128 202827 239180 202836
rect 239128 202793 239137 202827
rect 239137 202793 239171 202827
rect 239171 202793 239180 202827
rect 239128 202784 239180 202793
rect 267096 202784 267148 202836
rect 343732 202827 343784 202836
rect 343732 202793 343741 202827
rect 343741 202793 343775 202827
rect 343775 202793 343784 202827
rect 343732 202784 343784 202793
rect 298560 201492 298612 201544
rect 298652 201492 298704 201544
rect 234804 201467 234856 201476
rect 234804 201433 234813 201467
rect 234813 201433 234847 201467
rect 234847 201433 234856 201467
rect 234804 201424 234856 201433
rect 240416 201467 240468 201476
rect 240416 201433 240425 201467
rect 240425 201433 240459 201467
rect 240459 201433 240468 201467
rect 240416 201424 240468 201433
rect 291384 201424 291436 201476
rect 291660 201424 291712 201476
rect 305276 201467 305328 201476
rect 305276 201433 305285 201467
rect 305285 201433 305319 201467
rect 305319 201433 305328 201467
rect 305276 201424 305328 201433
rect 309324 201424 309376 201476
rect 310796 201424 310848 201476
rect 310888 201424 310940 201476
rect 313556 201424 313608 201476
rect 313648 201424 313700 201476
rect 345204 201424 345256 201476
rect 309416 201356 309468 201408
rect 267096 200064 267148 200116
rect 310796 200107 310848 200116
rect 310796 200073 310805 200107
rect 310805 200073 310839 200107
rect 310839 200073 310848 200107
rect 310796 200064 310848 200073
rect 238852 198475 238904 198484
rect 238852 198441 238861 198475
rect 238861 198441 238895 198475
rect 238895 198441 238904 198475
rect 238852 198432 238904 198441
rect 238852 198067 238904 198076
rect 238852 198033 238861 198067
rect 238861 198033 238895 198067
rect 238895 198033 238904 198067
rect 238852 198024 238904 198033
rect 254216 196596 254268 196648
rect 254400 196596 254452 196648
rect 298560 196052 298612 196104
rect 327356 196052 327408 196104
rect 273352 195984 273404 196036
rect 273536 195984 273588 196036
rect 288716 196027 288768 196036
rect 288716 195993 288725 196027
rect 288725 195993 288759 196027
rect 288759 195993 288768 196027
rect 288716 195984 288768 195993
rect 308036 196027 308088 196036
rect 308036 195993 308045 196027
rect 308045 195993 308079 196027
rect 308079 195993 308088 196027
rect 308036 195984 308088 195993
rect 434444 196027 434496 196036
rect 434444 195993 434453 196027
rect 434453 195993 434487 196027
rect 434487 195993 434496 196027
rect 434444 195984 434496 195993
rect 299848 195916 299900 195968
rect 305276 195959 305328 195968
rect 305276 195925 305285 195959
rect 305285 195925 305319 195959
rect 305319 195925 305328 195959
rect 305276 195916 305328 195925
rect 325976 195916 326028 195968
rect 327356 195916 327408 195968
rect 435180 195848 435232 195900
rect 435364 195848 435416 195900
rect 299848 195780 299900 195832
rect 325976 195780 326028 195832
rect 262588 193332 262640 193384
rect 345112 193264 345164 193316
rect 229376 193196 229428 193248
rect 229560 193196 229612 193248
rect 235080 193196 235132 193248
rect 239128 193196 239180 193248
rect 244096 193196 244148 193248
rect 244280 193196 244332 193248
rect 262588 193196 262640 193248
rect 287336 193196 287388 193248
rect 287520 193196 287572 193248
rect 288808 193196 288860 193248
rect 298468 193239 298520 193248
rect 298468 193205 298477 193239
rect 298477 193205 298511 193239
rect 298511 193205 298520 193239
rect 298468 193196 298520 193205
rect 308036 193239 308088 193248
rect 308036 193205 308045 193239
rect 308045 193205 308079 193239
rect 308079 193205 308088 193239
rect 308036 193196 308088 193205
rect 324596 193196 324648 193248
rect 324688 193196 324740 193248
rect 235264 193128 235316 193180
rect 362960 193196 363012 193248
rect 363236 193196 363288 193248
rect 434444 193239 434496 193248
rect 434444 193205 434453 193239
rect 434453 193205 434487 193239
rect 434487 193205 434496 193239
rect 434444 193196 434496 193205
rect 239220 193128 239272 193180
rect 240508 193128 240560 193180
rect 345112 193128 345164 193180
rect 345020 192763 345072 192772
rect 345020 192729 345029 192763
rect 345029 192729 345063 192763
rect 345063 192729 345072 192763
rect 345020 192720 345072 192729
rect 234804 192287 234856 192296
rect 234804 192253 234813 192287
rect 234813 192253 234847 192287
rect 234847 192253 234856 192287
rect 234804 192244 234856 192253
rect 251456 191836 251508 191888
rect 251548 191836 251600 191888
rect 316316 191836 316368 191888
rect 255596 191811 255648 191820
rect 255596 191777 255605 191811
rect 255605 191777 255639 191811
rect 255639 191777 255648 191811
rect 255596 191768 255648 191777
rect 262588 191811 262640 191820
rect 262588 191777 262597 191811
rect 262597 191777 262631 191811
rect 262631 191777 262640 191811
rect 262588 191768 262640 191777
rect 345020 190612 345072 190664
rect 345296 190612 345348 190664
rect 267004 190519 267056 190528
rect 267004 190485 267013 190519
rect 267013 190485 267047 190519
rect 267047 190485 267056 190519
rect 267004 190476 267056 190485
rect 316224 190519 316276 190528
rect 316224 190485 316233 190519
rect 316233 190485 316267 190519
rect 316267 190485 316276 190519
rect 316224 190476 316276 190485
rect 244280 189388 244332 189440
rect 244464 189388 244516 189440
rect 261208 186396 261260 186448
rect 233332 186328 233384 186380
rect 233516 186328 233568 186380
rect 238760 186328 238812 186380
rect 238944 186328 238996 186380
rect 276296 186396 276348 186448
rect 276112 186328 276164 186380
rect 288808 186371 288860 186380
rect 288808 186337 288817 186371
rect 288817 186337 288851 186371
rect 288851 186337 288860 186371
rect 288808 186328 288860 186337
rect 327356 186328 327408 186380
rect 346584 186328 346636 186380
rect 444012 186328 444064 186380
rect 444196 186328 444248 186380
rect 255596 186303 255648 186312
rect 255596 186269 255605 186303
rect 255605 186269 255639 186303
rect 255639 186269 255648 186303
rect 255596 186260 255648 186269
rect 261208 186260 261260 186312
rect 280436 186260 280488 186312
rect 280620 186260 280672 186312
rect 327448 186192 327500 186244
rect 346676 186192 346728 186244
rect 310428 185580 310480 185632
rect 241888 183608 241940 183660
rect 434444 183608 434496 183660
rect 234988 183540 235040 183592
rect 235264 183540 235316 183592
rect 239128 183540 239180 183592
rect 239220 183540 239272 183592
rect 241796 183540 241848 183592
rect 288808 183583 288860 183592
rect 288808 183549 288817 183583
rect 288817 183549 288851 183583
rect 288851 183549 288860 183583
rect 288808 183540 288860 183549
rect 305184 183540 305236 183592
rect 305460 183540 305512 183592
rect 308128 183540 308180 183592
rect 308312 183540 308364 183592
rect 342352 183540 342404 183592
rect 342536 183540 342588 183592
rect 347964 183540 348016 183592
rect 348148 183540 348200 183592
rect 434260 183540 434312 183592
rect 262588 183515 262640 183524
rect 262588 183481 262597 183515
rect 262597 183481 262631 183515
rect 262631 183481 262640 183515
rect 262588 183472 262640 183481
rect 343824 183472 343876 183524
rect 343916 183472 343968 183524
rect 316224 182180 316276 182232
rect 316316 182180 316368 182232
rect 239128 182155 239180 182164
rect 239128 182121 239137 182155
rect 239137 182121 239171 182155
rect 239171 182121 239180 182155
rect 239128 182112 239180 182121
rect 255688 182112 255740 182164
rect 324504 182112 324556 182164
rect 324688 182112 324740 182164
rect 343916 182112 343968 182164
rect 344100 182112 344152 182164
rect 309048 181024 309100 181076
rect 312084 181024 312136 181076
rect 398472 180956 398524 181008
rect 399024 180956 399076 181008
rect 417884 180956 417936 181008
rect 418344 180956 418396 181008
rect 338028 180888 338080 180940
rect 454408 180888 454460 180940
rect 458364 180888 458416 180940
rect 270500 180820 270552 180872
rect 275376 180820 275428 180872
rect 313648 180752 313700 180804
rect 313740 180752 313792 180804
rect 327448 180752 327500 180804
rect 338028 180752 338080 180804
rect 2780 179800 2832 179852
rect 5080 179800 5132 179852
rect 234988 179324 235040 179376
rect 235172 179324 235224 179376
rect 310796 179367 310848 179376
rect 310796 179333 310805 179367
rect 310805 179333 310839 179367
rect 310839 179333 310848 179367
rect 310796 179324 310848 179333
rect 241796 178823 241848 178832
rect 241796 178789 241805 178823
rect 241805 178789 241839 178823
rect 241839 178789 241848 178823
rect 241796 178780 241848 178789
rect 248788 176740 248840 176792
rect 288808 176740 288860 176792
rect 287244 176672 287296 176724
rect 238760 176604 238812 176656
rect 238944 176604 238996 176656
rect 248696 176604 248748 176656
rect 276112 176604 276164 176656
rect 287336 176604 287388 176656
rect 288808 176604 288860 176656
rect 276296 176536 276348 176588
rect 267096 173952 267148 174004
rect 299848 173952 299900 174004
rect 229376 173884 229428 173936
rect 229560 173884 229612 173936
rect 234804 173884 234856 173936
rect 234896 173884 234948 173936
rect 240416 173884 240468 173936
rect 240508 173884 240560 173936
rect 241796 173927 241848 173936
rect 241796 173893 241805 173927
rect 241805 173893 241839 173927
rect 241839 173893 241848 173927
rect 241796 173884 241848 173893
rect 244280 173884 244332 173936
rect 244464 173884 244516 173936
rect 261208 173884 261260 173936
rect 261300 173884 261352 173936
rect 262680 173884 262732 173936
rect 267004 173884 267056 173936
rect 291384 173884 291436 173936
rect 291476 173884 291528 173936
rect 299756 173884 299808 173936
rect 305368 173884 305420 173936
rect 305460 173884 305512 173936
rect 308036 173884 308088 173936
rect 308220 173884 308272 173936
rect 362960 173884 363012 173936
rect 363236 173884 363288 173936
rect 443920 173884 443972 173936
rect 444104 173884 444156 173936
rect 239128 173859 239180 173868
rect 239128 173825 239137 173859
rect 239137 173825 239171 173859
rect 239171 173825 239180 173859
rect 239128 173816 239180 173825
rect 262772 173748 262824 173800
rect 255596 172567 255648 172576
rect 255596 172533 255605 172567
rect 255605 172533 255639 172567
rect 255639 172533 255648 172567
rect 255596 172524 255648 172533
rect 251364 172456 251416 172508
rect 251456 172456 251508 172508
rect 299756 172456 299808 172508
rect 300032 172456 300084 172508
rect 327356 171139 327408 171148
rect 327356 171105 327365 171139
rect 327365 171105 327399 171139
rect 327399 171105 327408 171139
rect 327356 171096 327408 171105
rect 251364 171071 251416 171080
rect 251364 171037 251373 171071
rect 251373 171037 251407 171071
rect 251407 171037 251416 171071
rect 251364 171028 251416 171037
rect 313556 171071 313608 171080
rect 313556 171037 313565 171071
rect 313565 171037 313599 171071
rect 313599 171037 313608 171071
rect 313556 171028 313608 171037
rect 345020 171028 345072 171080
rect 345204 171028 345256 171080
rect 310888 169736 310940 169788
rect 239128 169056 239180 169108
rect 239312 169056 239364 169108
rect 233332 167016 233384 167068
rect 233516 167016 233568 167068
rect 238760 167016 238812 167068
rect 238944 167016 238996 167068
rect 346492 167016 346544 167068
rect 346676 167016 346728 167068
rect 435180 167016 435232 167068
rect 435364 167016 435416 167068
rect 2780 165452 2832 165504
rect 4988 165452 5040 165504
rect 435180 165044 435232 165096
rect 435548 165044 435600 165096
rect 255596 164228 255648 164280
rect 262680 164228 262732 164280
rect 262772 164228 262824 164280
rect 254216 164160 254268 164212
rect 254400 164160 254452 164212
rect 287336 164203 287388 164212
rect 287336 164169 287345 164203
rect 287345 164169 287379 164203
rect 287379 164169 287388 164203
rect 287336 164160 287388 164169
rect 324688 164160 324740 164212
rect 362960 164160 363012 164212
rect 363144 164160 363196 164212
rect 444104 164203 444156 164212
rect 444104 164169 444113 164203
rect 444113 164169 444147 164203
rect 444147 164169 444156 164203
rect 444104 164160 444156 164169
rect 255688 164092 255740 164144
rect 234988 162936 235040 162988
rect 235172 162936 235224 162988
rect 241888 162843 241940 162852
rect 241888 162809 241897 162843
rect 241897 162809 241931 162843
rect 241931 162809 241940 162843
rect 241888 162800 241940 162809
rect 261392 162800 261444 162852
rect 262680 162800 262732 162852
rect 288716 162800 288768 162852
rect 288808 162800 288860 162852
rect 305368 162800 305420 162852
rect 342536 162800 342588 162852
rect 342628 162800 342680 162852
rect 343916 162843 343968 162852
rect 343916 162809 343925 162843
rect 343925 162809 343959 162843
rect 343959 162809 343968 162843
rect 343916 162800 343968 162809
rect 345204 162843 345256 162852
rect 345204 162809 345213 162843
rect 345213 162809 345247 162843
rect 345247 162809 345256 162843
rect 345204 162800 345256 162809
rect 251456 161440 251508 161492
rect 313832 161440 313884 161492
rect 234988 161415 235040 161424
rect 234988 161381 234997 161415
rect 234997 161381 235031 161415
rect 235031 161381 235040 161415
rect 234988 161372 235040 161381
rect 288716 161415 288768 161424
rect 288716 161381 288725 161415
rect 288725 161381 288759 161415
rect 288759 161381 288768 161415
rect 288716 161372 288768 161381
rect 308128 161372 308180 161424
rect 310888 161372 310940 161424
rect 310980 161372 311032 161424
rect 234896 161347 234948 161356
rect 234896 161313 234905 161347
rect 234905 161313 234939 161347
rect 234939 161313 234948 161347
rect 234896 161304 234948 161313
rect 238852 159715 238904 159724
rect 238852 159681 238861 159715
rect 238861 159681 238895 159715
rect 238895 159681 238904 159715
rect 238852 159672 238904 159681
rect 238852 159375 238904 159384
rect 238852 159341 238861 159375
rect 238861 159341 238895 159375
rect 238895 159341 238904 159375
rect 238852 159332 238904 159341
rect 434444 159171 434496 159180
rect 434444 159137 434453 159171
rect 434453 159137 434487 159171
rect 434487 159137 434496 159171
rect 434444 159128 434496 159137
rect 229284 157360 229336 157412
rect 280528 157360 280580 157412
rect 229376 157292 229428 157344
rect 325976 157292 326028 157344
rect 444104 157335 444156 157344
rect 444104 157301 444113 157335
rect 444113 157301 444147 157335
rect 444147 157301 444156 157335
rect 444104 157292 444156 157301
rect 280620 157224 280672 157276
rect 325976 157156 326028 157208
rect 239128 154640 239180 154692
rect 255596 154640 255648 154692
rect 255688 154640 255740 154692
rect 240508 154572 240560 154624
rect 287336 154615 287388 154624
rect 287336 154581 287345 154615
rect 287345 154581 287379 154615
rect 287379 154581 287388 154615
rect 287336 154572 287388 154581
rect 324596 154615 324648 154624
rect 324596 154581 324605 154615
rect 324605 154581 324639 154615
rect 324639 154581 324648 154615
rect 324596 154572 324648 154581
rect 434444 154615 434496 154624
rect 434444 154581 434453 154615
rect 434453 154581 434487 154615
rect 434487 154581 434496 154615
rect 434444 154572 434496 154581
rect 229376 154504 229428 154556
rect 229560 154504 229612 154556
rect 245752 154504 245804 154556
rect 245936 154504 245988 154556
rect 290096 154504 290148 154556
rect 290188 154504 290240 154556
rect 316316 154504 316368 154556
rect 316408 154504 316460 154556
rect 347964 154504 348016 154556
rect 348148 154504 348200 154556
rect 444196 154504 444248 154556
rect 288808 153824 288860 153876
rect 327356 153527 327408 153536
rect 327356 153493 327365 153527
rect 327365 153493 327399 153527
rect 327399 153493 327408 153527
rect 327356 153484 327408 153493
rect 240416 153323 240468 153332
rect 240416 153289 240425 153323
rect 240425 153289 240459 153323
rect 240459 153289 240468 153323
rect 240416 153280 240468 153289
rect 241888 153255 241940 153264
rect 241888 153221 241897 153255
rect 241897 153221 241931 153255
rect 241931 153221 241940 153255
rect 241888 153212 241940 153221
rect 261300 153255 261352 153264
rect 261300 153221 261309 153255
rect 261309 153221 261343 153255
rect 261343 153221 261352 153255
rect 261300 153212 261352 153221
rect 262496 153255 262548 153264
rect 262496 153221 262505 153255
rect 262505 153221 262539 153255
rect 262539 153221 262548 153255
rect 262496 153212 262548 153221
rect 305276 153255 305328 153264
rect 305276 153221 305285 153255
rect 305285 153221 305319 153255
rect 305319 153221 305328 153255
rect 305276 153212 305328 153221
rect 343916 153255 343968 153264
rect 343916 153221 343925 153255
rect 343925 153221 343959 153255
rect 343959 153221 343968 153255
rect 343916 153212 343968 153221
rect 240416 153144 240468 153196
rect 255320 153144 255372 153196
rect 255596 153144 255648 153196
rect 305276 153119 305328 153128
rect 305276 153085 305285 153119
rect 305285 153085 305319 153119
rect 305319 153085 305328 153119
rect 305276 153076 305328 153085
rect 235080 151784 235132 151836
rect 239036 151827 239088 151836
rect 239036 151793 239045 151827
rect 239045 151793 239079 151827
rect 239079 151793 239088 151827
rect 239036 151784 239088 151793
rect 251180 151784 251232 151836
rect 251364 151784 251416 151836
rect 308036 151827 308088 151836
rect 308036 151793 308045 151827
rect 308045 151793 308079 151827
rect 308079 151793 308088 151827
rect 308036 151784 308088 151793
rect 313832 150560 313884 150612
rect 313648 150467 313700 150476
rect 313648 150433 313657 150467
rect 313657 150433 313691 150467
rect 313691 150433 313700 150467
rect 313648 150424 313700 150433
rect 288808 149039 288860 149048
rect 288808 149005 288817 149039
rect 288817 149005 288851 149039
rect 288851 149005 288860 149039
rect 288808 148996 288860 149005
rect 309508 149039 309560 149048
rect 309508 149005 309517 149039
rect 309517 149005 309551 149039
rect 309551 149005 309560 149039
rect 309508 148996 309560 149005
rect 343916 148316 343968 148368
rect 238944 147772 238996 147824
rect 435548 147772 435600 147824
rect 238852 147704 238904 147756
rect 233332 147636 233384 147688
rect 233516 147636 233568 147688
rect 324596 147704 324648 147756
rect 435456 147704 435508 147756
rect 280436 147636 280488 147688
rect 280620 147636 280672 147688
rect 238852 147568 238904 147620
rect 238944 147568 238996 147620
rect 324596 147568 324648 147620
rect 327356 147611 327408 147620
rect 327356 147577 327365 147611
rect 327365 147577 327399 147611
rect 327399 147577 327408 147611
rect 327356 147568 327408 147577
rect 434444 147568 434496 147620
rect 434720 147568 434772 147620
rect 435456 147568 435508 147620
rect 435548 147568 435600 147620
rect 287244 144984 287296 145036
rect 287336 144984 287388 145036
rect 444104 145027 444156 145036
rect 444104 144993 444113 145027
rect 444113 144993 444147 145027
rect 444147 144993 444156 145027
rect 444104 144984 444156 144993
rect 345296 144916 345348 144968
rect 241796 144848 241848 144900
rect 241980 144848 242032 144900
rect 244096 144848 244148 144900
rect 244280 144848 244332 144900
rect 254216 144848 254268 144900
rect 254400 144848 254452 144900
rect 240324 143599 240376 143608
rect 240324 143565 240333 143599
rect 240333 143565 240367 143599
rect 240367 143565 240376 143599
rect 240324 143556 240376 143565
rect 238760 143488 238812 143540
rect 238944 143488 238996 143540
rect 239036 143488 239088 143540
rect 239128 143488 239180 143540
rect 251364 143488 251416 143540
rect 287244 143531 287296 143540
rect 287244 143497 287253 143531
rect 287253 143497 287287 143531
rect 287287 143497 287296 143531
rect 287244 143488 287296 143497
rect 345204 143488 345256 143540
rect 345388 143488 345440 143540
rect 434444 143531 434496 143540
rect 434444 143497 434453 143531
rect 434453 143497 434487 143531
rect 434487 143497 434496 143531
rect 434444 143488 434496 143497
rect 444104 143531 444156 143540
rect 444104 143497 444113 143531
rect 444113 143497 444147 143531
rect 444147 143497 444156 143531
rect 444104 143488 444156 143497
rect 305368 142128 305420 142180
rect 239128 142103 239180 142112
rect 239128 142069 239137 142103
rect 239137 142069 239171 142103
rect 239171 142069 239180 142103
rect 239128 142060 239180 142069
rect 240324 142103 240376 142112
rect 240324 142069 240333 142103
rect 240333 142069 240367 142103
rect 240367 142069 240376 142103
rect 240324 142060 240376 142069
rect 316316 142103 316368 142112
rect 316316 142069 316325 142103
rect 316325 142069 316359 142103
rect 316359 142069 316368 142103
rect 316316 142060 316368 142069
rect 234804 140836 234856 140888
rect 234804 140743 234856 140752
rect 234804 140709 234813 140743
rect 234813 140709 234847 140743
rect 234847 140709 234856 140743
rect 234804 140700 234856 140709
rect 288808 139519 288860 139528
rect 288808 139485 288817 139519
rect 288817 139485 288851 139519
rect 288851 139485 288860 139519
rect 288808 139476 288860 139485
rect 309508 139451 309560 139460
rect 309508 139417 309517 139451
rect 309517 139417 309551 139451
rect 309551 139417 309560 139451
rect 309508 139408 309560 139417
rect 262680 139383 262732 139392
rect 262680 139349 262689 139383
rect 262689 139349 262723 139383
rect 262723 139349 262732 139383
rect 262680 139340 262732 139349
rect 288808 139340 288860 139392
rect 288900 139340 288952 139392
rect 229284 137980 229336 138032
rect 267188 138048 267240 138100
rect 435364 137980 435416 138032
rect 435548 137980 435600 138032
rect 229376 137912 229428 137964
rect 267096 137912 267148 137964
rect 434536 137912 434588 137964
rect 287428 137776 287480 137828
rect 2780 136348 2832 136400
rect 4896 136348 4948 136400
rect 343824 135303 343876 135312
rect 343824 135269 343833 135303
rect 343833 135269 343867 135303
rect 343867 135269 343876 135303
rect 343824 135260 343876 135269
rect 346584 135260 346636 135312
rect 346676 135260 346728 135312
rect 229376 135192 229428 135244
rect 229560 135192 229612 135244
rect 241888 135235 241940 135244
rect 241888 135201 241897 135235
rect 241897 135201 241931 135235
rect 241931 135201 241940 135235
rect 241888 135192 241940 135201
rect 245752 135192 245804 135244
rect 245936 135192 245988 135244
rect 251548 135235 251600 135244
rect 251548 135201 251557 135235
rect 251557 135201 251591 135235
rect 251591 135201 251600 135235
rect 251548 135192 251600 135201
rect 267096 135235 267148 135244
rect 267096 135201 267105 135235
rect 267105 135201 267139 135235
rect 267139 135201 267148 135235
rect 267096 135192 267148 135201
rect 327356 135235 327408 135244
rect 327356 135201 327365 135235
rect 327365 135201 327399 135235
rect 327399 135201 327408 135235
rect 327356 135192 327408 135201
rect 328552 135192 328604 135244
rect 328736 135192 328788 135244
rect 347964 135192 348016 135244
rect 348148 135192 348200 135244
rect 234988 134580 235040 134632
rect 309508 134512 309560 134564
rect 309692 134512 309744 134564
rect 269120 134104 269172 134156
rect 275376 134104 275428 134156
rect 357440 134036 357492 134088
rect 361120 134036 361172 134088
rect 398472 134036 398524 134088
rect 399024 134036 399076 134088
rect 417884 134036 417936 134088
rect 418344 134036 418396 134088
rect 317512 133968 317564 134020
rect 326896 133968 326948 134020
rect 251180 133900 251232 133952
rect 260748 133900 260800 133952
rect 308128 133900 308180 133952
rect 308220 133900 308272 133952
rect 327264 133900 327316 133952
rect 336648 133900 336700 133952
rect 251548 133832 251600 133884
rect 287336 133832 287388 133884
rect 287520 133832 287572 133884
rect 310796 133875 310848 133884
rect 310796 133841 310805 133875
rect 310805 133841 310839 133875
rect 310839 133841 310848 133875
rect 310796 133832 310848 133841
rect 233424 132515 233476 132524
rect 233424 132481 233433 132515
rect 233433 132481 233467 132515
rect 233467 132481 233476 132515
rect 233424 132472 233476 132481
rect 239128 132515 239180 132524
rect 239128 132481 239137 132515
rect 239137 132481 239171 132515
rect 239171 132481 239180 132515
rect 239128 132472 239180 132481
rect 240416 132472 240468 132524
rect 316316 132515 316368 132524
rect 316316 132481 316325 132515
rect 316325 132481 316359 132515
rect 316359 132481 316368 132515
rect 316316 132472 316368 132481
rect 305368 132447 305420 132456
rect 305368 132413 305377 132447
rect 305377 132413 305411 132447
rect 305411 132413 305420 132447
rect 305368 132404 305420 132413
rect 233424 131155 233476 131164
rect 233424 131121 233433 131155
rect 233433 131121 233467 131155
rect 233467 131121 233476 131155
rect 233424 131112 233476 131121
rect 324596 131044 324648 131096
rect 324872 131044 324924 131096
rect 255504 130432 255556 130484
rect 255780 130432 255832 130484
rect 262864 129752 262916 129804
rect 235080 128367 235132 128376
rect 235080 128333 235089 128367
rect 235089 128333 235123 128367
rect 235123 128333 235132 128367
rect 235080 128324 235132 128333
rect 238760 128256 238812 128308
rect 238944 128256 238996 128308
rect 267096 128299 267148 128308
rect 267096 128265 267105 128299
rect 267105 128265 267139 128299
rect 267139 128265 267148 128299
rect 267096 128256 267148 128265
rect 327356 128299 327408 128308
rect 327356 128265 327365 128299
rect 327365 128265 327399 128299
rect 327399 128265 327408 128299
rect 327356 128256 327408 128265
rect 444104 128299 444156 128308
rect 444104 128265 444113 128299
rect 444113 128265 444147 128299
rect 444147 128265 444156 128299
rect 444104 128256 444156 128265
rect 241888 125647 241940 125656
rect 241888 125613 241897 125647
rect 241897 125613 241931 125647
rect 241931 125613 241940 125647
rect 241888 125604 241940 125613
rect 345204 125604 345256 125656
rect 345388 125604 345440 125656
rect 254216 125579 254268 125588
rect 254216 125545 254225 125579
rect 254225 125545 254259 125579
rect 254259 125545 254268 125579
rect 254216 125536 254268 125545
rect 328460 125579 328512 125588
rect 328460 125545 328469 125579
rect 328469 125545 328503 125579
rect 328503 125545 328512 125579
rect 347964 125579 348016 125588
rect 328460 125536 328512 125545
rect 347964 125545 347973 125579
rect 347973 125545 348007 125579
rect 348007 125545 348016 125579
rect 347964 125536 348016 125545
rect 435364 125536 435416 125588
rect 435548 125536 435600 125588
rect 444104 125536 444156 125588
rect 233424 125511 233476 125520
rect 233424 125477 233433 125511
rect 233433 125477 233467 125511
rect 233467 125477 233476 125511
rect 233424 125468 233476 125477
rect 316316 124244 316368 124296
rect 251456 124219 251508 124228
rect 251456 124185 251465 124219
rect 251465 124185 251499 124219
rect 251499 124185 251508 124219
rect 251456 124176 251508 124185
rect 291568 124219 291620 124228
rect 291568 124185 291577 124219
rect 291577 124185 291611 124219
rect 291611 124185 291620 124219
rect 291568 124176 291620 124185
rect 310796 124219 310848 124228
rect 310796 124185 310805 124219
rect 310805 124185 310839 124219
rect 310839 124185 310848 124219
rect 310796 124176 310848 124185
rect 316224 124176 316276 124228
rect 241888 124151 241940 124160
rect 241888 124117 241897 124151
rect 241897 124117 241931 124151
rect 241931 124117 241940 124151
rect 241888 124108 241940 124117
rect 261300 124108 261352 124160
rect 287244 124108 287296 124160
rect 345204 124151 345256 124160
rect 345204 124117 345213 124151
rect 345213 124117 345247 124151
rect 345247 124117 345256 124151
rect 345204 124108 345256 124117
rect 287428 124040 287480 124092
rect 252836 123564 252888 123616
rect 252744 123496 252796 123548
rect 235080 122859 235132 122868
rect 235080 122825 235089 122859
rect 235089 122825 235123 122859
rect 235123 122825 235132 122859
rect 235080 122816 235132 122825
rect 305368 122859 305420 122868
rect 305368 122825 305377 122859
rect 305377 122825 305411 122859
rect 305411 122825 305420 122859
rect 305368 122816 305420 122825
rect 240416 122748 240468 122800
rect 2780 122068 2832 122120
rect 4804 122068 4856 122120
rect 233424 121499 233476 121508
rect 233424 121465 233433 121499
rect 233433 121465 233467 121499
rect 233467 121465 233476 121499
rect 233424 121456 233476 121465
rect 291568 121499 291620 121508
rect 291568 121465 291577 121499
rect 291577 121465 291611 121499
rect 291611 121465 291620 121499
rect 291568 121456 291620 121465
rect 309416 120096 309468 120148
rect 309692 120096 309744 120148
rect 234896 120071 234948 120080
rect 234896 120037 234905 120071
rect 234905 120037 234939 120071
rect 234939 120037 234948 120071
rect 234896 120028 234948 120037
rect 262864 120028 262916 120080
rect 292856 118736 292908 118788
rect 305000 118736 305052 118788
rect 305368 118736 305420 118788
rect 229284 118668 229336 118720
rect 267004 118668 267056 118720
rect 267188 118668 267240 118720
rect 280528 118668 280580 118720
rect 229376 118600 229428 118652
rect 261208 118643 261260 118652
rect 261208 118609 261217 118643
rect 261217 118609 261251 118643
rect 261251 118609 261260 118643
rect 261208 118600 261260 118609
rect 280620 118600 280672 118652
rect 292856 118600 292908 118652
rect 328552 118600 328604 118652
rect 444196 118643 444248 118652
rect 444196 118609 444205 118643
rect 444205 118609 444239 118643
rect 444239 118609 444248 118643
rect 444196 118600 444248 118609
rect 347964 116059 348016 116068
rect 347964 116025 347973 116059
rect 347973 116025 348007 116059
rect 348007 116025 348016 116059
rect 347964 116016 348016 116025
rect 254216 115991 254268 116000
rect 254216 115957 254225 115991
rect 254225 115957 254259 115991
rect 254259 115957 254268 115991
rect 254216 115948 254268 115957
rect 229376 115880 229428 115932
rect 245936 115923 245988 115932
rect 245936 115889 245945 115923
rect 245945 115889 245979 115923
rect 245979 115889 245988 115923
rect 245936 115880 245988 115889
rect 267004 115880 267056 115932
rect 267188 115880 267240 115932
rect 298468 115923 298520 115932
rect 298468 115889 298477 115923
rect 298477 115889 298511 115923
rect 298511 115889 298520 115923
rect 298468 115880 298520 115889
rect 347964 115880 348016 115932
rect 348148 115880 348200 115932
rect 309324 115243 309376 115252
rect 309324 115209 309333 115243
rect 309333 115209 309367 115243
rect 309367 115209 309376 115243
rect 309324 115200 309376 115209
rect 310796 114588 310848 114640
rect 241888 114563 241940 114572
rect 241888 114529 241897 114563
rect 241897 114529 241931 114563
rect 241931 114529 241940 114563
rect 241888 114520 241940 114529
rect 234988 114452 235040 114504
rect 235080 114452 235132 114504
rect 255596 114495 255648 114504
rect 255596 114461 255605 114495
rect 255605 114461 255639 114495
rect 255639 114461 255648 114495
rect 255596 114452 255648 114461
rect 287336 114495 287388 114504
rect 287336 114461 287345 114495
rect 287345 114461 287379 114495
rect 287379 114461 287388 114495
rect 287336 114452 287388 114461
rect 288716 114495 288768 114504
rect 288716 114461 288725 114495
rect 288725 114461 288759 114495
rect 288759 114461 288768 114495
rect 288716 114452 288768 114461
rect 316224 114520 316276 114572
rect 316316 114520 316368 114572
rect 345204 114563 345256 114572
rect 345204 114529 345213 114563
rect 345213 114529 345247 114563
rect 345247 114529 345256 114563
rect 345204 114520 345256 114529
rect 310888 114452 310940 114504
rect 342536 114495 342588 114504
rect 342536 114461 342545 114495
rect 342545 114461 342579 114495
rect 342579 114461 342588 114495
rect 342536 114452 342588 114461
rect 313648 113135 313700 113144
rect 313648 113101 313657 113135
rect 313657 113101 313691 113135
rect 313691 113101 313700 113135
rect 313648 113092 313700 113101
rect 241612 111052 241664 111104
rect 241888 111052 241940 111104
rect 239128 109080 239180 109132
rect 238760 109012 238812 109064
rect 238944 109012 238996 109064
rect 238944 108876 238996 108928
rect 280436 109012 280488 109064
rect 280620 109012 280672 109064
rect 434352 109012 434404 109064
rect 435364 109012 435416 109064
rect 435548 109012 435600 109064
rect 444012 109012 444064 109064
rect 444196 109012 444248 109064
rect 434444 108944 434496 108996
rect 298560 108808 298612 108860
rect 229284 106335 229336 106344
rect 229284 106301 229293 106335
rect 229293 106301 229327 106335
rect 229327 106301 229336 106335
rect 229284 106292 229336 106301
rect 245936 106335 245988 106344
rect 245936 106301 245945 106335
rect 245945 106301 245979 106335
rect 245979 106301 245988 106335
rect 245936 106292 245988 106301
rect 324688 106335 324740 106344
rect 324688 106301 324697 106335
rect 324697 106301 324731 106335
rect 324731 106301 324740 106335
rect 324688 106292 324740 106301
rect 305276 106267 305328 106276
rect 305276 106233 305285 106267
rect 305285 106233 305319 106267
rect 305319 106233 305328 106267
rect 305276 106224 305328 106233
rect 347964 106267 348016 106276
rect 347964 106233 347973 106267
rect 347973 106233 348007 106267
rect 348007 106233 348016 106267
rect 347964 106224 348016 106233
rect 444104 106267 444156 106276
rect 444104 106233 444113 106267
rect 444113 106233 444147 106267
rect 444147 106233 444156 106267
rect 444104 106224 444156 106233
rect 342536 104975 342588 104984
rect 342536 104941 342545 104975
rect 342545 104941 342579 104975
rect 342579 104941 342588 104975
rect 342536 104932 342588 104941
rect 240324 104907 240376 104916
rect 240324 104873 240333 104907
rect 240333 104873 240367 104907
rect 240367 104873 240376 104907
rect 240324 104864 240376 104873
rect 255596 104907 255648 104916
rect 255596 104873 255605 104907
rect 255605 104873 255639 104907
rect 255639 104873 255648 104907
rect 255596 104864 255648 104873
rect 287336 104907 287388 104916
rect 287336 104873 287345 104907
rect 287345 104873 287379 104907
rect 287379 104873 287388 104907
rect 287336 104864 287388 104873
rect 288808 104864 288860 104916
rect 324688 104907 324740 104916
rect 324688 104873 324697 104907
rect 324697 104873 324731 104907
rect 324731 104873 324740 104907
rect 324688 104864 324740 104873
rect 234988 104796 235040 104848
rect 235080 104796 235132 104848
rect 241796 104839 241848 104848
rect 241796 104805 241805 104839
rect 241805 104805 241839 104839
rect 241839 104805 241848 104839
rect 241796 104796 241848 104805
rect 251456 104839 251508 104848
rect 251456 104805 251465 104839
rect 251465 104805 251499 104839
rect 251499 104805 251508 104839
rect 251456 104796 251508 104805
rect 280528 104839 280580 104848
rect 280528 104805 280537 104839
rect 280537 104805 280571 104839
rect 280571 104805 280580 104839
rect 280528 104796 280580 104805
rect 327448 104796 327500 104848
rect 342536 104839 342588 104848
rect 342536 104805 342545 104839
rect 342545 104805 342579 104839
rect 342579 104805 342588 104839
rect 342536 104796 342588 104805
rect 345204 104839 345256 104848
rect 345204 104805 345213 104839
rect 345213 104805 345247 104839
rect 345247 104805 345256 104839
rect 345204 104796 345256 104805
rect 434444 104796 434496 104848
rect 305092 103572 305144 103624
rect 305092 103436 305144 103488
rect 308036 103436 308088 103488
rect 308128 103436 308180 103488
rect 310888 103436 310940 103488
rect 311072 103436 311124 103488
rect 309324 102459 309376 102468
rect 309324 102425 309333 102459
rect 309333 102425 309367 102459
rect 309367 102425 309376 102459
rect 309324 102416 309376 102425
rect 313464 102416 313516 102468
rect 262680 102187 262732 102196
rect 262680 102153 262689 102187
rect 262689 102153 262723 102187
rect 262723 102153 262732 102187
rect 262680 102144 262732 102153
rect 305276 102187 305328 102196
rect 305276 102153 305285 102187
rect 305285 102153 305319 102187
rect 305319 102153 305328 102187
rect 305276 102144 305328 102153
rect 267096 102076 267148 102128
rect 238944 100036 238996 100088
rect 239128 100036 239180 100088
rect 262680 99424 262732 99476
rect 288808 99424 288860 99476
rect 290096 99424 290148 99476
rect 229284 99356 229336 99408
rect 298560 99424 298612 99476
rect 324688 99424 324740 99476
rect 229376 99288 229428 99340
rect 290096 99288 290148 99340
rect 298468 99288 298520 99340
rect 324596 99288 324648 99340
rect 444104 99331 444156 99340
rect 444104 99297 444113 99331
rect 444113 99297 444147 99331
rect 444147 99297 444156 99331
rect 444104 99288 444156 99297
rect 255596 98676 255648 98728
rect 345388 98676 345440 98728
rect 347964 96747 348016 96756
rect 347964 96713 347973 96747
rect 347973 96713 348007 96747
rect 348007 96713 348016 96747
rect 347964 96704 348016 96713
rect 229376 96568 229428 96620
rect 347964 96568 348016 96620
rect 348056 96568 348108 96620
rect 251456 95319 251508 95328
rect 251456 95285 251465 95319
rect 251465 95285 251499 95319
rect 251499 95285 251508 95319
rect 251456 95276 251508 95285
rect 241888 95208 241940 95260
rect 280620 95208 280672 95260
rect 327356 95251 327408 95260
rect 327356 95217 327365 95251
rect 327365 95217 327399 95251
rect 327399 95217 327408 95251
rect 327356 95208 327408 95217
rect 342536 95251 342588 95260
rect 342536 95217 342545 95251
rect 342545 95217 342579 95251
rect 342579 95217 342588 95251
rect 342536 95208 342588 95217
rect 434352 95251 434404 95260
rect 434352 95217 434361 95251
rect 434361 95217 434395 95251
rect 434395 95217 434404 95251
rect 434352 95208 434404 95217
rect 240416 95140 240468 95192
rect 240508 95140 240560 95192
rect 251180 95140 251232 95192
rect 251456 95140 251508 95192
rect 244464 94639 244516 94648
rect 244464 94605 244473 94639
rect 244473 94605 244507 94639
rect 244507 94605 244516 94639
rect 244464 94596 244516 94605
rect 248696 94639 248748 94648
rect 248696 94605 248705 94639
rect 248705 94605 248739 94639
rect 248739 94605 248748 94639
rect 248696 94596 248748 94605
rect 255688 93891 255740 93900
rect 255688 93857 255697 93891
rect 255697 93857 255731 93891
rect 255731 93857 255740 93891
rect 255688 93848 255740 93857
rect 240508 93823 240560 93832
rect 240508 93789 240517 93823
rect 240517 93789 240551 93823
rect 240551 93789 240560 93823
rect 240508 93780 240560 93789
rect 345388 93780 345440 93832
rect 255688 93755 255740 93764
rect 255688 93721 255697 93755
rect 255697 93721 255731 93755
rect 255731 93721 255740 93755
rect 255688 93712 255740 93721
rect 234804 92055 234856 92064
rect 234804 92021 234813 92055
rect 234813 92021 234847 92055
rect 234847 92021 234856 92055
rect 234804 92012 234856 92021
rect 434352 91783 434404 91792
rect 434352 91749 434361 91783
rect 434361 91749 434395 91783
rect 434395 91749 434404 91783
rect 434352 91740 434404 91749
rect 309416 89811 309468 89820
rect 309416 89777 309425 89811
rect 309425 89777 309459 89811
rect 309459 89777 309468 89811
rect 309416 89768 309468 89777
rect 233332 89700 233384 89752
rect 233516 89700 233568 89752
rect 280436 89700 280488 89752
rect 280620 89700 280672 89752
rect 444012 89700 444064 89752
rect 444196 89700 444248 89752
rect 434628 87320 434680 87372
rect 282828 87184 282880 87236
rect 292764 87184 292816 87236
rect 356060 87116 356112 87168
rect 365628 87116 365680 87168
rect 417884 87116 417936 87168
rect 418344 87116 418396 87168
rect 434536 87116 434588 87168
rect 434628 87116 434680 87168
rect 398472 87048 398524 87100
rect 398840 87048 398892 87100
rect 229284 87023 229336 87032
rect 229284 86989 229293 87023
rect 229293 86989 229327 87023
rect 229327 86989 229336 87023
rect 229284 86980 229336 86989
rect 305552 86980 305604 87032
rect 444380 86980 444432 87032
rect 449256 86980 449308 87032
rect 463792 86980 463844 87032
rect 466552 86980 466604 87032
rect 262496 86955 262548 86964
rect 262496 86921 262505 86955
rect 262505 86921 262539 86955
rect 262539 86921 262548 86955
rect 262496 86912 262548 86921
rect 298468 86912 298520 86964
rect 298560 86912 298612 86964
rect 305460 86912 305512 86964
rect 343732 86912 343784 86964
rect 343824 86912 343876 86964
rect 363052 86912 363104 86964
rect 444104 86955 444156 86964
rect 444104 86921 444113 86955
rect 444113 86921 444147 86955
rect 444147 86921 444156 86955
rect 444104 86912 444156 86921
rect 327356 86887 327408 86896
rect 327356 86853 327365 86887
rect 327365 86853 327399 86887
rect 327399 86853 327408 86887
rect 327356 86844 327408 86853
rect 288624 86139 288676 86148
rect 288624 86105 288633 86139
rect 288633 86105 288667 86139
rect 288667 86105 288676 86139
rect 288624 86096 288676 86105
rect 244464 85595 244516 85604
rect 244464 85561 244473 85595
rect 244473 85561 244507 85595
rect 244507 85561 244516 85595
rect 244464 85552 244516 85561
rect 248788 85552 248840 85604
rect 287336 85552 287388 85604
rect 287428 85552 287480 85604
rect 309416 85595 309468 85604
rect 309416 85561 309425 85595
rect 309425 85561 309459 85595
rect 309459 85561 309468 85595
rect 309416 85552 309468 85561
rect 313464 85552 313516 85604
rect 313648 85552 313700 85604
rect 343732 85527 343784 85536
rect 343732 85493 343741 85527
rect 343741 85493 343775 85527
rect 343775 85493 343784 85527
rect 343732 85484 343784 85493
rect 435180 85527 435232 85536
rect 435180 85493 435189 85527
rect 435189 85493 435223 85527
rect 435223 85493 435232 85527
rect 435180 85484 435232 85493
rect 240416 84192 240468 84244
rect 255780 84192 255832 84244
rect 291476 84192 291528 84244
rect 291568 84192 291620 84244
rect 234804 84167 234856 84176
rect 234804 84133 234813 84167
rect 234813 84133 234847 84167
rect 234847 84133 234856 84167
rect 234804 84124 234856 84133
rect 307944 84167 307996 84176
rect 307944 84133 307953 84167
rect 307953 84133 307987 84167
rect 307987 84133 307996 84167
rect 307944 84124 307996 84133
rect 313648 84167 313700 84176
rect 313648 84133 313657 84167
rect 313657 84133 313691 84167
rect 313691 84133 313700 84167
rect 313648 84124 313700 84133
rect 267096 82832 267148 82884
rect 324596 82356 324648 82408
rect 324596 82220 324648 82272
rect 287336 80112 287388 80164
rect 342536 80112 342588 80164
rect 229284 80044 229336 80096
rect 254216 80044 254268 80096
rect 299848 80044 299900 80096
rect 325976 80044 326028 80096
rect 287336 79976 287388 80028
rect 342536 79976 342588 80028
rect 229376 79908 229428 79960
rect 254216 79908 254268 79960
rect 299848 79908 299900 79960
rect 325976 79908 326028 79960
rect 2780 79432 2832 79484
rect 6184 79432 6236 79484
rect 291568 79296 291620 79348
rect 267096 77979 267148 77988
rect 267096 77945 267105 77979
rect 267105 77945 267139 77979
rect 267139 77945 267148 77979
rect 267096 77936 267148 77945
rect 255596 77528 255648 77580
rect 255780 77528 255832 77580
rect 233424 77256 233476 77308
rect 233516 77256 233568 77308
rect 234988 77256 235040 77308
rect 235080 77256 235132 77308
rect 244464 77256 244516 77308
rect 244556 77256 244608 77308
rect 327356 77299 327408 77308
rect 327356 77265 327365 77299
rect 327365 77265 327399 77299
rect 327399 77265 327408 77299
rect 327356 77256 327408 77265
rect 362960 77299 363012 77308
rect 362960 77265 362969 77299
rect 362969 77265 363003 77299
rect 363003 77265 363012 77299
rect 362960 77256 363012 77265
rect 444196 77256 444248 77308
rect 261116 77188 261168 77240
rect 262496 77188 262548 77240
rect 262864 77188 262916 77240
rect 261300 77120 261352 77172
rect 362960 77163 363012 77172
rect 362960 77129 362969 77163
rect 362969 77129 363003 77163
rect 363003 77129 363012 77163
rect 362960 77120 363012 77129
rect 343732 76007 343784 76016
rect 343732 75973 343741 76007
rect 343741 75973 343775 76007
rect 343775 75973 343784 76007
rect 343732 75964 343784 75973
rect 290096 75896 290148 75948
rect 345204 75939 345256 75948
rect 345204 75905 345213 75939
rect 345213 75905 345247 75939
rect 345247 75905 345256 75939
rect 345204 75896 345256 75905
rect 435180 75939 435232 75948
rect 435180 75905 435189 75939
rect 435189 75905 435223 75939
rect 435223 75905 435232 75939
rect 435180 75896 435232 75905
rect 240416 75828 240468 75880
rect 244464 75828 244516 75880
rect 244556 75828 244608 75880
rect 248788 75871 248840 75880
rect 248788 75837 248797 75871
rect 248797 75837 248831 75871
rect 248831 75837 248840 75871
rect 248788 75828 248840 75837
rect 262864 75828 262916 75880
rect 343732 75871 343784 75880
rect 343732 75837 343741 75871
rect 343741 75837 343775 75871
rect 343775 75837 343784 75871
rect 343732 75828 343784 75837
rect 434352 75828 434404 75880
rect 290188 75760 290240 75812
rect 234804 74579 234856 74588
rect 234804 74545 234813 74579
rect 234813 74545 234847 74579
rect 234847 74545 234856 74579
rect 234804 74536 234856 74545
rect 305276 74536 305328 74588
rect 305460 74536 305512 74588
rect 308128 74536 308180 74588
rect 313740 74536 313792 74588
rect 229376 74468 229428 74520
rect 348056 74468 348108 74520
rect 305276 74443 305328 74452
rect 305276 74409 305285 74443
rect 305285 74409 305319 74443
rect 305319 74409 305328 74443
rect 305276 74400 305328 74409
rect 288624 73788 288676 73840
rect 280528 73176 280580 73228
rect 280620 73176 280672 73228
rect 290004 70864 290056 70916
rect 290188 70864 290240 70916
rect 276296 70456 276348 70508
rect 287336 70456 287388 70508
rect 328552 70456 328604 70508
rect 346584 70456 346636 70508
rect 276112 70388 276164 70440
rect 287336 70320 287388 70372
rect 328552 70320 328604 70372
rect 346584 70320 346636 70372
rect 363052 70252 363104 70304
rect 324596 67736 324648 67788
rect 435180 67736 435232 67788
rect 325976 67668 326028 67720
rect 267096 67643 267148 67652
rect 267096 67609 267105 67643
rect 267105 67609 267139 67643
rect 267139 67609 267148 67643
rect 267096 67600 267148 67609
rect 324596 67600 324648 67652
rect 325884 67600 325936 67652
rect 327356 67643 327408 67652
rect 327356 67609 327365 67643
rect 327365 67609 327399 67643
rect 327399 67609 327408 67643
rect 327356 67600 327408 67609
rect 435180 67600 435232 67652
rect 444104 67600 444156 67652
rect 444196 67600 444248 67652
rect 244280 67575 244332 67584
rect 244280 67541 244289 67575
rect 244289 67541 244323 67575
rect 244323 67541 244332 67575
rect 244280 67532 244332 67541
rect 252744 67532 252796 67584
rect 252836 67532 252888 67584
rect 240416 66308 240468 66360
rect 434260 66351 434312 66360
rect 434260 66317 434269 66351
rect 434269 66317 434303 66351
rect 434303 66317 434312 66351
rect 434260 66308 434312 66317
rect 248788 66283 248840 66292
rect 248788 66249 248797 66283
rect 248797 66249 248831 66283
rect 248831 66249 248840 66283
rect 248788 66240 248840 66249
rect 262772 66283 262824 66292
rect 262772 66249 262781 66283
rect 262781 66249 262815 66283
rect 262815 66249 262824 66283
rect 262772 66240 262824 66249
rect 308036 66283 308088 66292
rect 255596 66215 255648 66224
rect 255596 66181 255605 66215
rect 255605 66181 255639 66215
rect 255639 66181 255648 66215
rect 255596 66172 255648 66181
rect 291476 66104 291528 66156
rect 308036 66249 308045 66283
rect 308045 66249 308079 66283
rect 308079 66249 308088 66283
rect 308036 66240 308088 66249
rect 327356 66283 327408 66292
rect 327356 66249 327365 66283
rect 327365 66249 327399 66283
rect 327399 66249 327408 66283
rect 327356 66240 327408 66249
rect 343916 66240 343968 66292
rect 309324 66172 309376 66224
rect 309416 66172 309468 66224
rect 324596 66215 324648 66224
rect 324596 66181 324605 66215
rect 324605 66181 324639 66215
rect 324639 66181 324648 66215
rect 324596 66172 324648 66181
rect 345204 66215 345256 66224
rect 345204 66181 345213 66215
rect 345213 66181 345247 66215
rect 345247 66181 345256 66215
rect 345204 66172 345256 66181
rect 434260 66172 434312 66224
rect 435180 66215 435232 66224
rect 435180 66181 435189 66215
rect 435189 66181 435223 66215
rect 435223 66181 435232 66215
rect 435180 66172 435232 66181
rect 434444 66104 434496 66156
rect 229284 64991 229336 65000
rect 229284 64957 229293 64991
rect 229293 64957 229327 64991
rect 229327 64957 229336 64991
rect 229284 64948 229336 64957
rect 233424 64880 233476 64932
rect 233516 64880 233568 64932
rect 305368 64880 305420 64932
rect 308036 64923 308088 64932
rect 308036 64889 308045 64923
rect 308045 64889 308079 64923
rect 308079 64889 308088 64923
rect 308036 64880 308088 64889
rect 310888 64880 310940 64932
rect 310980 64880 311032 64932
rect 347964 64923 348016 64932
rect 347964 64889 347973 64923
rect 347973 64889 348007 64923
rect 348007 64889 348016 64923
rect 347964 64880 348016 64889
rect 229284 64812 229336 64864
rect 229468 64812 229520 64864
rect 234804 64855 234856 64864
rect 234804 64821 234813 64855
rect 234813 64821 234847 64855
rect 234847 64821 234856 64855
rect 234804 64812 234856 64821
rect 240416 64812 240468 64864
rect 292764 64812 292816 64864
rect 292856 64812 292908 64864
rect 255780 64676 255832 64728
rect 326804 63724 326856 63776
rect 335268 63724 335320 63776
rect 398472 63724 398524 63776
rect 399024 63724 399076 63776
rect 359556 63656 359608 63708
rect 365628 63656 365680 63708
rect 417884 63656 417936 63708
rect 419632 63656 419684 63708
rect 280252 63452 280304 63504
rect 280528 63452 280580 63504
rect 267096 61072 267148 61124
rect 261300 60800 261352 60852
rect 444104 60800 444156 60852
rect 261208 60664 261260 60716
rect 273352 60664 273404 60716
rect 336924 60664 336976 60716
rect 337108 60664 337160 60716
rect 363052 60664 363104 60716
rect 363236 60664 363288 60716
rect 444012 60664 444064 60716
rect 273536 60596 273588 60648
rect 310796 58760 310848 58812
rect 310980 58760 311032 58812
rect 325884 58012 325936 58064
rect 244280 57987 244332 57996
rect 244280 57953 244289 57987
rect 244289 57953 244323 57987
rect 244323 57953 244332 57987
rect 244280 57944 244332 57953
rect 287336 57944 287388 57996
rect 287428 57944 287480 57996
rect 288716 57987 288768 57996
rect 288716 57953 288725 57987
rect 288725 57953 288759 57987
rect 288759 57953 288768 57987
rect 288716 57944 288768 57953
rect 239128 57876 239180 57928
rect 245936 57919 245988 57928
rect 245936 57885 245945 57919
rect 245945 57885 245979 57919
rect 245979 57885 245988 57919
rect 245936 57876 245988 57885
rect 325884 57876 325936 57928
rect 337108 57876 337160 57928
rect 363236 57876 363288 57928
rect 313740 56652 313792 56704
rect 249984 56584 250036 56636
rect 250076 56584 250128 56636
rect 262680 56584 262732 56636
rect 262864 56584 262916 56636
rect 267004 56627 267056 56636
rect 267004 56593 267013 56627
rect 267013 56593 267047 56627
rect 267047 56593 267056 56627
rect 267004 56584 267056 56593
rect 309416 56584 309468 56636
rect 254124 56559 254176 56568
rect 254124 56525 254133 56559
rect 254133 56525 254167 56559
rect 254167 56525 254176 56559
rect 254124 56516 254176 56525
rect 262680 56448 262732 56500
rect 262864 56448 262916 56500
rect 345204 56627 345256 56636
rect 345204 56593 345213 56627
rect 345213 56593 345247 56627
rect 345247 56593 345256 56627
rect 345204 56584 345256 56593
rect 313740 56516 313792 56568
rect 309508 56448 309560 56500
rect 290096 55292 290148 55344
rect 234804 55267 234856 55276
rect 234804 55233 234813 55267
rect 234813 55233 234847 55267
rect 234847 55233 234856 55267
rect 234804 55224 234856 55233
rect 240324 55267 240376 55276
rect 240324 55233 240333 55267
rect 240333 55233 240367 55267
rect 240367 55233 240376 55267
rect 240324 55224 240376 55233
rect 290004 55224 290056 55276
rect 255780 55156 255832 55208
rect 347964 55156 348016 55208
rect 290004 55131 290056 55140
rect 290004 55097 290013 55131
rect 290013 55097 290047 55131
rect 290047 55097 290056 55131
rect 290004 55088 290056 55097
rect 252744 53116 252796 53168
rect 261208 53159 261260 53168
rect 261208 53125 261217 53159
rect 261217 53125 261251 53159
rect 261251 53125 261260 53159
rect 261208 53116 261260 53125
rect 327356 53116 327408 53168
rect 252836 53048 252888 53100
rect 324780 53048 324832 53100
rect 327264 53048 327316 53100
rect 229376 51076 229428 51128
rect 287336 51212 287388 51264
rect 299848 51187 299900 51196
rect 299848 51153 299857 51187
rect 299857 51153 299891 51187
rect 299891 51153 299900 51187
rect 299848 51144 299900 51153
rect 342536 51187 342588 51196
rect 342536 51153 342545 51187
rect 342545 51153 342579 51187
rect 342579 51153 342588 51187
rect 342536 51144 342588 51153
rect 346584 51187 346636 51196
rect 346584 51153 346593 51187
rect 346593 51153 346627 51187
rect 346627 51153 346636 51187
rect 346584 51144 346636 51153
rect 434352 51076 434404 51128
rect 229284 51008 229336 51060
rect 239036 51051 239088 51060
rect 239036 51017 239045 51051
rect 239045 51017 239079 51051
rect 239079 51017 239088 51051
rect 239036 51008 239088 51017
rect 287244 51008 287296 51060
rect 434260 51008 434312 51060
rect 435180 51051 435232 51060
rect 435180 51017 435189 51051
rect 435189 51017 435223 51051
rect 435223 51017 435232 51051
rect 435180 51008 435232 51017
rect 444012 51008 444064 51060
rect 444196 51008 444248 51060
rect 240324 48288 240376 48340
rect 240416 48288 240468 48340
rect 245936 48331 245988 48340
rect 245936 48297 245945 48331
rect 245945 48297 245979 48331
rect 245979 48297 245988 48331
rect 245936 48288 245988 48297
rect 261300 48288 261352 48340
rect 299848 48331 299900 48340
rect 299848 48297 299857 48331
rect 299857 48297 299891 48331
rect 299891 48297 299900 48331
rect 299848 48288 299900 48297
rect 336924 48331 336976 48340
rect 336924 48297 336933 48331
rect 336933 48297 336967 48331
rect 336967 48297 336976 48331
rect 336924 48288 336976 48297
rect 363144 48331 363196 48340
rect 363144 48297 363153 48331
rect 363153 48297 363187 48331
rect 363187 48297 363196 48331
rect 363144 48288 363196 48297
rect 239036 48220 239088 48272
rect 239128 48220 239180 48272
rect 267188 48220 267240 48272
rect 288624 48220 288676 48272
rect 288808 48220 288860 48272
rect 435272 48263 435324 48272
rect 435272 48229 435281 48263
rect 435281 48229 435315 48263
rect 435315 48229 435324 48263
rect 435272 48220 435324 48229
rect 444196 48220 444248 48272
rect 254124 46971 254176 46980
rect 254124 46937 254133 46971
rect 254133 46937 254167 46971
rect 254167 46937 254176 46971
rect 254124 46928 254176 46937
rect 291476 46928 291528 46980
rect 291568 46928 291620 46980
rect 342536 46971 342588 46980
rect 342536 46937 342545 46971
rect 342545 46937 342579 46971
rect 342579 46937 342588 46971
rect 342536 46928 342588 46937
rect 251364 46860 251416 46912
rect 251456 46860 251508 46912
rect 262864 46903 262916 46912
rect 262864 46869 262873 46903
rect 262873 46869 262907 46903
rect 262907 46869 262916 46903
rect 345204 46903 345256 46912
rect 262864 46860 262916 46869
rect 345204 46869 345213 46903
rect 345213 46869 345247 46903
rect 345247 46869 345256 46903
rect 345204 46860 345256 46869
rect 325884 46792 325936 46844
rect 326160 46792 326212 46844
rect 255596 45679 255648 45688
rect 255596 45645 255605 45679
rect 255605 45645 255639 45679
rect 255639 45645 255648 45679
rect 255596 45636 255648 45645
rect 347964 45636 348016 45688
rect 290004 45611 290056 45620
rect 290004 45577 290013 45611
rect 290013 45577 290047 45611
rect 290047 45577 290056 45611
rect 290004 45568 290056 45577
rect 346584 45611 346636 45620
rect 346584 45577 346593 45611
rect 346593 45577 346627 45611
rect 346627 45577 346636 45611
rect 346584 45568 346636 45577
rect 234804 45543 234856 45552
rect 234804 45509 234813 45543
rect 234813 45509 234847 45543
rect 234847 45509 234856 45543
rect 234804 45500 234856 45509
rect 234988 45500 235040 45552
rect 235172 45500 235224 45552
rect 255596 45500 255648 45552
rect 255688 45500 255740 45552
rect 299848 45500 299900 45552
rect 299940 45500 299992 45552
rect 280252 44480 280304 44532
rect 241796 44115 241848 44124
rect 241796 44081 241805 44115
rect 241805 44081 241839 44115
rect 241839 44081 241848 44115
rect 241796 44072 241848 44081
rect 229284 41463 229336 41472
rect 229284 41429 229293 41463
rect 229293 41429 229327 41463
rect 229327 41429 229336 41463
rect 229284 41420 229336 41429
rect 313556 41420 313608 41472
rect 313740 41420 313792 41472
rect 363052 41352 363104 41404
rect 363236 41352 363288 41404
rect 270500 40332 270552 40384
rect 280528 40332 280580 40384
rect 398472 40196 398524 40248
rect 399024 40196 399076 40248
rect 417884 40196 417936 40248
rect 418344 40196 418396 40248
rect 356060 40060 356112 40112
rect 365628 40060 365680 40112
rect 229376 38700 229428 38752
rect 287244 38700 287296 38752
rect 267096 38675 267148 38684
rect 267096 38641 267105 38675
rect 267105 38641 267139 38675
rect 267139 38641 267148 38675
rect 267096 38632 267148 38641
rect 273260 38632 273312 38684
rect 273536 38632 273588 38684
rect 435364 38632 435416 38684
rect 444104 38675 444156 38684
rect 444104 38641 444113 38675
rect 444113 38641 444147 38675
rect 444147 38641 444156 38675
rect 444104 38632 444156 38641
rect 245936 38607 245988 38616
rect 245936 38573 245945 38607
rect 245945 38573 245979 38607
rect 245979 38573 245988 38607
rect 245936 38564 245988 38573
rect 287244 38564 287296 38616
rect 324780 38564 324832 38616
rect 363236 38564 363288 38616
rect 324780 38428 324832 38480
rect 254124 37272 254176 37324
rect 254216 37272 254268 37324
rect 262680 37272 262732 37324
rect 267096 37204 267148 37256
rect 234804 35955 234856 35964
rect 234804 35921 234813 35955
rect 234813 35921 234847 35955
rect 234847 35921 234856 35955
rect 234804 35912 234856 35921
rect 290004 35887 290056 35896
rect 290004 35853 290013 35887
rect 290013 35853 290047 35887
rect 290047 35853 290056 35887
rect 290004 35844 290056 35853
rect 299756 35844 299808 35896
rect 300032 35844 300084 35896
rect 305368 35887 305420 35896
rect 305368 35853 305377 35887
rect 305377 35853 305411 35887
rect 305411 35853 305420 35887
rect 305368 35844 305420 35853
rect 434444 35071 434496 35080
rect 434444 35037 434453 35071
rect 434453 35037 434487 35071
rect 434487 35037 434496 35071
rect 434444 35028 434496 35037
rect 307944 34484 307996 34536
rect 308128 34484 308180 34536
rect 253940 32376 253992 32428
rect 254216 32376 254268 32428
rect 328552 31875 328604 31884
rect 328552 31841 328561 31875
rect 328561 31841 328595 31875
rect 328595 31841 328604 31875
rect 328552 31832 328604 31841
rect 444104 31875 444156 31884
rect 444104 31841 444113 31875
rect 444113 31841 444147 31875
rect 444147 31841 444156 31875
rect 444104 31832 444156 31841
rect 229284 31764 229336 31816
rect 261208 31807 261260 31816
rect 261208 31773 261217 31807
rect 261217 31773 261251 31807
rect 261251 31773 261260 31807
rect 261208 31764 261260 31773
rect 229376 31628 229428 31680
rect 292856 30676 292908 30728
rect 270500 29180 270552 29232
rect 273996 29180 274048 29232
rect 398472 29180 398524 29232
rect 399024 29180 399076 29232
rect 476028 29180 476080 29232
rect 482928 29180 482980 29232
rect 417884 29112 417936 29164
rect 418160 29112 418212 29164
rect 342444 29044 342496 29096
rect 434536 29044 434588 29096
rect 444380 29044 444432 29096
rect 449256 29044 449308 29096
rect 241796 29019 241848 29028
rect 241796 28985 241805 29019
rect 241805 28985 241839 29019
rect 241839 28985 241848 29019
rect 241796 28976 241848 28985
rect 245936 29019 245988 29028
rect 245936 28985 245945 29019
rect 245945 28985 245979 29019
rect 245979 28985 245988 29019
rect 245936 28976 245988 28985
rect 342536 28976 342588 29028
rect 345296 28976 345348 29028
rect 363144 29019 363196 29028
rect 363144 28985 363153 29019
rect 363153 28985 363187 29019
rect 363187 28985 363196 29019
rect 363144 28976 363196 28985
rect 444104 29019 444156 29028
rect 444104 28985 444113 29019
rect 444113 28985 444147 29019
rect 444147 28985 444156 29019
rect 444104 28976 444156 28985
rect 298560 28908 298612 28960
rect 298652 28908 298704 28960
rect 324596 28951 324648 28960
rect 324596 28917 324605 28951
rect 324605 28917 324639 28951
rect 324639 28917 324648 28951
rect 324596 28908 324648 28917
rect 327264 28908 327316 28960
rect 327448 28908 327500 28960
rect 435364 28908 435416 28960
rect 280528 28883 280580 28892
rect 280528 28849 280537 28883
rect 280537 28849 280571 28883
rect 280571 28849 280580 28883
rect 280528 28840 280580 28849
rect 261208 27659 261260 27668
rect 261208 27625 261217 27659
rect 261217 27625 261251 27659
rect 261251 27625 261260 27659
rect 261208 27616 261260 27625
rect 267004 27659 267056 27668
rect 267004 27625 267013 27659
rect 267013 27625 267047 27659
rect 267047 27625 267056 27659
rect 267004 27616 267056 27625
rect 328552 27659 328604 27668
rect 328552 27625 328561 27659
rect 328561 27625 328595 27659
rect 328595 27625 328604 27659
rect 328552 27616 328604 27625
rect 251456 27548 251508 27600
rect 342536 27548 342588 27600
rect 345296 27548 345348 27600
rect 434536 27548 434588 27600
rect 290188 26256 290240 26308
rect 292764 26299 292816 26308
rect 292764 26265 292773 26299
rect 292773 26265 292807 26299
rect 292807 26265 292816 26299
rect 292764 26256 292816 26265
rect 234804 26231 234856 26240
rect 234804 26197 234813 26231
rect 234813 26197 234847 26231
rect 234847 26197 234856 26231
rect 234804 26188 234856 26197
rect 235080 26188 235132 26240
rect 239128 26188 239180 26240
rect 346584 26188 346636 26240
rect 305368 24871 305420 24880
rect 305368 24837 305377 24871
rect 305377 24837 305411 24871
rect 305411 24837 305420 24871
rect 305368 24828 305420 24837
rect 262680 24148 262732 24200
rect 252836 22720 252888 22772
rect 253940 22720 253992 22772
rect 255320 22720 255372 22772
rect 255688 22720 255740 22772
rect 328552 22720 328604 22772
rect 245936 22108 245988 22160
rect 245752 22040 245804 22092
rect 363052 22040 363104 22092
rect 363236 22040 363288 22092
rect 308128 19499 308180 19508
rect 308128 19465 308137 19499
rect 308137 19465 308171 19499
rect 308171 19465 308180 19499
rect 308128 19456 308180 19465
rect 244556 19388 244608 19440
rect 248788 19388 248840 19440
rect 244464 19320 244516 19372
rect 248696 19320 248748 19372
rect 249984 19320 250036 19372
rect 250076 19320 250128 19372
rect 261116 19320 261168 19372
rect 261208 19320 261260 19372
rect 262588 19363 262640 19372
rect 262588 19329 262597 19363
rect 262597 19329 262631 19363
rect 262631 19329 262640 19363
rect 262588 19320 262640 19329
rect 288716 19320 288768 19372
rect 288992 19320 289044 19372
rect 292764 19320 292816 19372
rect 292856 19320 292908 19372
rect 324596 19363 324648 19372
rect 324596 19329 324605 19363
rect 324605 19329 324639 19363
rect 324639 19329 324648 19363
rect 324596 19320 324648 19329
rect 435272 19363 435324 19372
rect 435272 19329 435281 19363
rect 435281 19329 435315 19363
rect 435315 19329 435324 19363
rect 435272 19320 435324 19329
rect 327356 19252 327408 19304
rect 363236 19295 363288 19304
rect 363236 19261 363245 19295
rect 363245 19261 363279 19295
rect 363279 19261 363288 19295
rect 363236 19252 363288 19261
rect 310796 18028 310848 18080
rect 229376 17892 229428 17944
rect 240324 17892 240376 17944
rect 241612 17935 241664 17944
rect 241612 17901 241621 17935
rect 241621 17901 241655 17935
rect 241655 17901 241664 17935
rect 241612 17892 241664 17901
rect 280436 17960 280488 18012
rect 280528 17960 280580 18012
rect 310704 17960 310756 18012
rect 434536 17960 434588 18012
rect 251548 17892 251600 17944
rect 434536 17008 434588 17060
rect 434628 17008 434680 17060
rect 398472 16804 398524 16856
rect 399024 16804 399076 16856
rect 434536 16804 434588 16856
rect 434628 16804 434680 16856
rect 476028 16804 476080 16856
rect 482928 16804 482980 16856
rect 360016 16736 360068 16788
rect 361120 16736 361172 16788
rect 300032 16668 300084 16720
rect 425060 16668 425112 16720
rect 434444 16668 434496 16720
rect 444380 16668 444432 16720
rect 447232 16668 447284 16720
rect 234896 16643 234948 16652
rect 234896 16609 234905 16643
rect 234905 16609 234939 16643
rect 234939 16609 234948 16643
rect 234896 16600 234948 16609
rect 346400 16643 346452 16652
rect 346400 16609 346409 16643
rect 346409 16609 346443 16643
rect 346443 16609 346452 16643
rect 346400 16600 346452 16609
rect 299848 15215 299900 15224
rect 299848 15181 299857 15215
rect 299857 15181 299891 15215
rect 299891 15181 299900 15215
rect 299848 15172 299900 15181
rect 107476 15104 107528 15156
rect 269212 15104 269264 15156
rect 103428 15036 103480 15088
rect 267832 15036 267884 15088
rect 99288 14968 99340 15020
rect 266452 14968 266504 15020
rect 96528 14900 96580 14952
rect 265072 14900 265124 14952
rect 92388 14832 92440 14884
rect 263692 14832 263744 14884
rect 89628 14764 89680 14816
rect 262588 14764 262640 14816
rect 85488 14696 85540 14748
rect 261116 14696 261168 14748
rect 82728 14628 82780 14680
rect 259552 14628 259604 14680
rect 78588 14560 78640 14612
rect 258172 14560 258224 14612
rect 74448 14492 74500 14544
rect 256792 14492 256844 14544
rect 31668 14424 31720 14476
rect 241704 14424 241756 14476
rect 110328 14356 110380 14408
rect 270592 14356 270644 14408
rect 114468 14288 114520 14340
rect 271972 14288 272024 14340
rect 117228 14220 117280 14272
rect 273352 14220 273404 14272
rect 121368 14152 121420 14204
rect 274732 14152 274784 14204
rect 125416 14084 125468 14136
rect 276112 14084 276164 14136
rect 197268 14016 197320 14068
rect 303896 14016 303948 14068
rect 190368 13744 190420 13796
rect 301044 13744 301096 13796
rect 186228 13676 186280 13728
rect 299664 13676 299716 13728
rect 183468 13608 183520 13660
rect 298284 13608 298336 13660
rect 179328 13540 179380 13592
rect 296996 13540 297048 13592
rect 176568 13472 176620 13524
rect 295616 13472 295668 13524
rect 172428 13404 172480 13456
rect 294236 13404 294288 13456
rect 160008 13336 160060 13388
rect 288716 13336 288768 13388
rect 155868 13268 155920 13320
rect 287336 13268 287388 13320
rect 135168 13200 135220 13252
rect 280344 13200 280396 13252
rect 71688 13132 71740 13184
rect 255412 13132 255464 13184
rect 23388 13064 23440 13116
rect 237472 13064 237524 13116
rect 194508 12996 194560 13048
rect 302424 12996 302476 13048
rect 211068 12928 211120 12980
rect 213828 12860 213880 12912
rect 309324 12860 309376 12912
rect 217968 12792 218020 12844
rect 310704 12792 310756 12844
rect 220728 12724 220780 12776
rect 312176 12724 312228 12776
rect 224868 12656 224920 12708
rect 313556 12656 313608 12708
rect 229008 12588 229060 12640
rect 314936 12588 314988 12640
rect 316224 12520 316276 12572
rect 234712 12495 234764 12504
rect 234712 12461 234721 12495
rect 234721 12461 234755 12495
rect 234755 12461 234764 12495
rect 234712 12452 234764 12461
rect 290096 12495 290148 12504
rect 290096 12461 290105 12495
rect 290105 12461 290139 12495
rect 290139 12461 290148 12495
rect 290096 12452 290148 12461
rect 325976 12452 326028 12504
rect 173808 12384 173860 12436
rect 294052 12384 294104 12436
rect 325884 12384 325936 12436
rect 169392 12316 169444 12368
rect 292948 12316 293000 12368
rect 328552 12316 328604 12368
rect 165896 12248 165948 12300
rect 291660 12248 291712 12300
rect 162308 12180 162360 12232
rect 151728 12112 151780 12164
rect 285864 12112 285916 12164
rect 148968 12044 149020 12096
rect 285956 12044 286008 12096
rect 144828 11976 144880 12028
rect 284484 11976 284536 12028
rect 140872 11908 140924 11960
rect 283104 11908 283156 11960
rect 128268 11840 128320 11892
rect 277492 11840 277544 11892
rect 126888 11772 126940 11824
rect 277584 11772 277636 11824
rect 18328 11704 18380 11756
rect 236092 11704 236144 11756
rect 176384 11636 176436 11688
rect 295432 11636 295484 11688
rect 180708 11568 180760 11620
rect 296812 11568 296864 11620
rect 184756 11500 184808 11552
rect 298652 11500 298704 11552
rect 187608 11432 187660 11484
rect 299848 11432 299900 11484
rect 191748 11364 191800 11416
rect 300952 11364 301004 11416
rect 194416 11296 194468 11348
rect 302332 11296 302384 11348
rect 198648 11228 198700 11280
rect 303804 11228 303856 11280
rect 234712 11203 234764 11212
rect 234712 11169 234721 11203
rect 234721 11169 234755 11203
rect 234755 11169 234764 11203
rect 234712 11160 234764 11169
rect 108948 10956 109000 11008
rect 270684 10956 270736 11008
rect 106188 10888 106240 10940
rect 269304 10888 269356 10940
rect 102048 10820 102100 10872
rect 267924 10820 267976 10872
rect 99196 10752 99248 10804
rect 266544 10752 266596 10804
rect 95148 10684 95200 10736
rect 265164 10684 265216 10736
rect 91008 10616 91060 10668
rect 263784 10616 263836 10668
rect 63592 10548 63644 10600
rect 252652 10548 252704 10600
rect 60004 10480 60056 10532
rect 251272 10480 251324 10532
rect 56416 10412 56468 10464
rect 249892 10412 249944 10464
rect 52828 10344 52880 10396
rect 248604 10344 248656 10396
rect 49332 10276 49384 10328
rect 248512 10276 248564 10328
rect 113088 10208 113140 10260
rect 272064 10208 272116 10260
rect 117136 10140 117188 10192
rect 273444 10140 273496 10192
rect 119988 10072 120040 10124
rect 274824 10072 274876 10124
rect 124128 10004 124180 10056
rect 276204 10004 276256 10056
rect 154488 9936 154540 9988
rect 287152 9936 287204 9988
rect 158628 9868 158680 9920
rect 288532 9868 288584 9920
rect 161388 9800 161440 9852
rect 289912 9800 289964 9852
rect 231308 9707 231360 9716
rect 231308 9673 231317 9707
rect 231317 9673 231351 9707
rect 231351 9673 231360 9707
rect 231308 9664 231360 9673
rect 252744 9707 252796 9716
rect 252744 9673 252753 9707
rect 252753 9673 252787 9707
rect 252787 9673 252796 9707
rect 252744 9664 252796 9673
rect 254124 9707 254176 9716
rect 254124 9673 254133 9707
rect 254133 9673 254167 9707
rect 254167 9673 254176 9707
rect 254124 9664 254176 9673
rect 327264 9707 327316 9716
rect 327264 9673 327273 9707
rect 327273 9673 327307 9707
rect 327307 9673 327316 9707
rect 327264 9664 327316 9673
rect 342444 9707 342496 9716
rect 342444 9673 342453 9707
rect 342453 9673 342487 9707
rect 342487 9673 342496 9707
rect 342444 9664 342496 9673
rect 345204 9707 345256 9716
rect 345204 9673 345213 9707
rect 345213 9673 345247 9707
rect 345247 9673 345256 9707
rect 345204 9664 345256 9673
rect 363236 9707 363288 9716
rect 363236 9673 363245 9707
rect 363245 9673 363279 9707
rect 363279 9673 363288 9707
rect 363236 9664 363288 9673
rect 203892 9596 203944 9648
rect 306564 9596 306616 9648
rect 405556 9596 405608 9648
rect 463240 9596 463292 9648
rect 200396 9528 200448 9580
rect 305092 9528 305144 9580
rect 406936 9528 406988 9580
rect 466828 9528 466880 9580
rect 150440 9460 150492 9512
rect 285772 9460 285824 9512
rect 408316 9460 408368 9512
rect 470324 9460 470376 9512
rect 146852 9392 146904 9444
rect 284392 9392 284444 9444
rect 439964 9392 440016 9444
rect 555976 9392 556028 9444
rect 143264 9324 143316 9376
rect 283012 9324 283064 9376
rect 441436 9324 441488 9376
rect 559564 9324 559616 9376
rect 139676 9256 139728 9308
rect 281724 9256 281776 9308
rect 442724 9256 442776 9308
rect 563152 9256 563204 9308
rect 136088 9188 136140 9240
rect 280436 9188 280488 9240
rect 444012 9188 444064 9240
rect 566740 9188 566792 9240
rect 44548 9120 44600 9172
rect 245752 9120 245804 9172
rect 250352 9120 250404 9172
rect 323216 9120 323268 9172
rect 445484 9120 445536 9172
rect 570236 9120 570288 9172
rect 40960 9052 41012 9104
rect 244464 9052 244516 9104
rect 246764 9052 246816 9104
rect 323124 9052 323176 9104
rect 446956 9052 447008 9104
rect 573824 9052 573876 9104
rect 27896 8984 27948 9036
rect 233884 8984 233936 9036
rect 239588 8984 239640 9036
rect 320364 8984 320416 9036
rect 448336 8984 448388 9036
rect 577412 8984 577464 9036
rect 13636 8916 13688 8968
rect 236000 8916 236052 8968
rect 318984 8916 319036 8968
rect 400036 8916 400088 8968
rect 448980 8916 449032 8968
rect 449716 8916 449768 8968
rect 581000 8916 581052 8968
rect 207480 8848 207532 8900
rect 307852 8848 307904 8900
rect 404176 8848 404228 8900
rect 459652 8848 459704 8900
rect 210884 8780 210936 8832
rect 309232 8780 309284 8832
rect 402796 8780 402848 8832
rect 456064 8780 456116 8832
rect 214656 8712 214708 8764
rect 310612 8712 310664 8764
rect 401416 8712 401468 8764
rect 452476 8712 452528 8764
rect 218152 8644 218204 8696
rect 311992 8644 312044 8696
rect 221740 8576 221792 8628
rect 313372 8576 313424 8628
rect 225328 8508 225380 8560
rect 314752 8508 314804 8560
rect 228916 8440 228968 8492
rect 316132 8440 316184 8492
rect 232504 8372 232556 8424
rect 317604 8372 317656 8424
rect 229192 8347 229244 8356
rect 229192 8313 229201 8347
rect 229201 8313 229235 8347
rect 229235 8313 229244 8347
rect 229192 8304 229244 8313
rect 234896 8304 234948 8356
rect 235080 8304 235132 8356
rect 239036 8304 239088 8356
rect 240232 8347 240284 8356
rect 240232 8313 240241 8347
rect 240241 8313 240275 8347
rect 240275 8313 240284 8347
rect 240232 8304 240284 8313
rect 241704 8304 241756 8356
rect 243176 8304 243228 8356
rect 321744 8304 321796 8356
rect 129004 8236 129056 8288
rect 277400 8236 277452 8288
rect 420736 8236 420788 8288
rect 504824 8236 504876 8288
rect 87328 8168 87380 8220
rect 262404 8168 262456 8220
rect 267004 8168 267056 8220
rect 329932 8168 329984 8220
rect 391480 8168 391532 8220
rect 391756 8168 391808 8220
rect 422116 8168 422168 8220
rect 508412 8168 508464 8220
rect 83832 8100 83884 8152
rect 261024 8100 261076 8152
rect 263416 8100 263468 8152
rect 328460 8100 328512 8152
rect 427636 8100 427688 8152
rect 523868 8100 523920 8152
rect 80244 8032 80296 8084
rect 259736 8032 259788 8084
rect 259828 8032 259880 8084
rect 327264 8032 327316 8084
rect 429016 8032 429068 8084
rect 527456 8032 527508 8084
rect 37372 7964 37424 8016
rect 243084 7964 243136 8016
rect 256240 7964 256292 8016
rect 325884 7964 325936 8016
rect 430396 7964 430448 8016
rect 531044 7964 531096 8016
rect 33876 7896 33928 7948
rect 241704 7896 241756 7948
rect 252652 7896 252704 7948
rect 324596 7896 324648 7948
rect 431776 7896 431828 7948
rect 534540 7896 534592 7948
rect 30288 7828 30340 7880
rect 240232 7828 240284 7880
rect 249156 7828 249208 7880
rect 323032 7828 323084 7880
rect 433156 7828 433208 7880
rect 538128 7828 538180 7880
rect 26700 7760 26752 7812
rect 239036 7760 239088 7812
rect 245568 7760 245620 7812
rect 321652 7760 321704 7812
rect 434536 7760 434588 7812
rect 541716 7760 541768 7812
rect 21916 7692 21968 7744
rect 237656 7692 237708 7744
rect 241980 7692 242032 7744
rect 320272 7692 320324 7744
rect 435916 7692 435968 7744
rect 545304 7692 545356 7744
rect 17224 7624 17276 7676
rect 236184 7624 236236 7676
rect 238392 7624 238444 7676
rect 319168 7624 319220 7676
rect 437296 7624 437348 7676
rect 548892 7624 548944 7676
rect 8852 7556 8904 7608
rect 227720 7556 227772 7608
rect 229008 7556 229060 7608
rect 234804 7556 234856 7608
rect 317788 7556 317840 7608
rect 438676 7556 438728 7608
rect 552388 7556 552440 7608
rect 138480 7488 138532 7540
rect 281816 7488 281868 7540
rect 419356 7488 419408 7540
rect 501236 7488 501288 7540
rect 142068 7420 142120 7472
rect 283196 7420 283248 7472
rect 417976 7420 418028 7472
rect 497740 7420 497792 7472
rect 145656 7352 145708 7404
rect 284576 7352 284628 7404
rect 416504 7352 416556 7404
rect 494152 7352 494204 7404
rect 149244 7284 149296 7336
rect 286048 7284 286100 7336
rect 415216 7284 415268 7336
rect 490564 7284 490616 7336
rect 152740 7216 152792 7268
rect 287060 7216 287112 7268
rect 413836 7216 413888 7268
rect 486976 7216 487028 7268
rect 156328 7148 156380 7200
rect 288440 7148 288492 7200
rect 412548 7148 412600 7200
rect 483480 7148 483532 7200
rect 158720 7080 158772 7132
rect 160008 7080 160060 7132
rect 159916 7012 159968 7064
rect 289820 7080 289872 7132
rect 398564 7080 398616 7132
rect 445392 7080 445444 7132
rect 164700 7012 164752 7064
rect 291292 7012 291344 7064
rect 168196 6944 168248 6996
rect 292672 6944 292724 6996
rect 175372 6876 175424 6928
rect 176568 6876 176620 6928
rect 193220 6876 193272 6928
rect 194508 6876 194560 6928
rect 209872 6876 209924 6928
rect 211068 6876 211120 6928
rect 232044 6876 232096 6928
rect 348056 6876 348108 6928
rect 348240 6876 348292 6928
rect 174176 6808 174228 6860
rect 295340 6808 295392 6860
rect 413928 6808 413980 6860
rect 484584 6808 484636 6860
rect 170588 6740 170640 6792
rect 293960 6740 294012 6792
rect 415308 6740 415360 6792
rect 488172 6740 488224 6792
rect 167092 6672 167144 6724
rect 292580 6672 292632 6724
rect 416596 6672 416648 6724
rect 491760 6672 491812 6724
rect 163504 6604 163556 6656
rect 291200 6604 291252 6656
rect 416688 6604 416740 6656
rect 495348 6604 495400 6656
rect 131396 6536 131448 6588
rect 279056 6536 279108 6588
rect 418068 6536 418120 6588
rect 498936 6536 498988 6588
rect 76656 6468 76708 6520
rect 258356 6468 258408 6520
rect 419448 6468 419500 6520
rect 502432 6468 502484 6520
rect 73068 6400 73120 6452
rect 256976 6400 257028 6452
rect 305000 6400 305052 6452
rect 343732 6400 343784 6452
rect 420828 6400 420880 6452
rect 506020 6400 506072 6452
rect 69480 6332 69532 6384
rect 255412 6332 255464 6384
rect 284208 6332 284260 6384
rect 334164 6332 334216 6384
rect 422208 6332 422260 6384
rect 509608 6332 509660 6384
rect 65984 6264 66036 6316
rect 254032 6264 254084 6316
rect 261024 6264 261076 6316
rect 327172 6264 327224 6316
rect 423496 6264 423548 6316
rect 513196 6264 513248 6316
rect 62396 6196 62448 6248
rect 252744 6196 252796 6248
rect 257436 6196 257488 6248
rect 325792 6196 325844 6248
rect 424876 6196 424928 6248
rect 516784 6196 516836 6248
rect 58808 6128 58860 6180
rect 251272 6128 251324 6180
rect 253848 6128 253900 6180
rect 324412 6128 324464 6180
rect 426256 6128 426308 6180
rect 520280 6128 520332 6180
rect 177764 6060 177816 6112
rect 296720 6060 296772 6112
rect 411168 6060 411220 6112
rect 479892 6060 479944 6112
rect 181352 5992 181404 6044
rect 298100 5992 298152 6044
rect 409788 5992 409840 6044
rect 476304 5992 476356 6044
rect 184848 5924 184900 5976
rect 299480 5924 299532 5976
rect 408408 5924 408460 5976
rect 472716 5924 472768 5976
rect 188436 5856 188488 5908
rect 300860 5856 300912 5908
rect 407028 5856 407080 5908
rect 469128 5856 469180 5908
rect 192024 5788 192076 5840
rect 302240 5788 302292 5840
rect 405648 5788 405700 5840
rect 465632 5788 465684 5840
rect 195612 5720 195664 5772
rect 303620 5720 303672 5772
rect 404268 5720 404320 5772
rect 462044 5720 462096 5772
rect 199200 5652 199252 5704
rect 303712 5652 303764 5704
rect 402888 5652 402940 5704
rect 458456 5652 458508 5704
rect 202696 5584 202748 5636
rect 305184 5584 305236 5636
rect 401508 5584 401560 5636
rect 454868 5584 454920 5636
rect 206284 5516 206336 5568
rect 306472 5516 306524 5568
rect 137284 5448 137336 5500
rect 281540 5448 281592 5500
rect 290740 5448 290792 5500
rect 339592 5448 339644 5500
rect 390376 5448 390428 5500
rect 423956 5448 424008 5500
rect 434628 5448 434680 5500
rect 540520 5448 540572 5500
rect 133788 5380 133840 5432
rect 280160 5380 280212 5432
rect 287152 5380 287204 5432
rect 338212 5380 338264 5432
rect 391664 5380 391716 5432
rect 426348 5380 426400 5432
rect 436008 5380 436060 5432
rect 544108 5380 544160 5432
rect 130200 5312 130252 5364
rect 278780 5312 278832 5364
rect 283656 5312 283708 5364
rect 336832 5312 336884 5364
rect 393044 5312 393096 5364
rect 429936 5312 429988 5364
rect 437388 5312 437440 5364
rect 547696 5312 547748 5364
rect 67180 5244 67232 5296
rect 254124 5244 254176 5296
rect 280068 5244 280120 5296
rect 335544 5244 335596 5296
rect 394516 5244 394568 5296
rect 433524 5244 433576 5296
rect 438768 5244 438820 5296
rect 551192 5244 551244 5296
rect 51632 5176 51684 5228
rect 248696 5176 248748 5228
rect 251456 5176 251508 5228
rect 324320 5176 324372 5228
rect 394424 5176 394476 5228
rect 434628 5176 434680 5228
rect 440056 5176 440108 5228
rect 554780 5176 554832 5228
rect 48136 5108 48188 5160
rect 247132 5108 247184 5160
rect 247960 5108 248012 5160
rect 323308 5108 323360 5160
rect 395804 5108 395856 5160
rect 437020 5108 437072 5160
rect 441528 5108 441580 5160
rect 558368 5108 558420 5160
rect 12440 5040 12492 5092
rect 233240 5040 233292 5092
rect 244372 5040 244424 5092
rect 321836 5040 321888 5092
rect 395896 5040 395948 5092
rect 438216 5040 438268 5092
rect 442816 5040 442868 5092
rect 561956 5040 562008 5092
rect 7656 4972 7708 5024
rect 231952 4972 232004 5024
rect 240784 4972 240836 5024
rect 320456 4972 320508 5024
rect 397368 4972 397420 5024
rect 440608 4972 440660 5024
rect 444288 4972 444340 5024
rect 565544 4972 565596 5024
rect 2872 4904 2924 4956
rect 237196 4904 237248 4956
rect 318708 4904 318760 4956
rect 318800 4904 318852 4956
rect 346400 4904 346452 4956
rect 398656 4904 398708 4956
rect 444196 4904 444248 4956
rect 445576 4904 445628 4956
rect 569040 4904 569092 4956
rect 229192 4836 229244 4888
rect 572 4768 624 4820
rect 230480 4836 230532 4888
rect 233700 4836 233752 4888
rect 317420 4836 317472 4888
rect 320180 4836 320232 4888
rect 347872 4836 347924 4888
rect 397276 4836 397328 4888
rect 441804 4836 441856 4888
rect 447048 4836 447100 4888
rect 572628 4836 572680 4888
rect 230112 4768 230164 4820
rect 316040 4768 316092 4820
rect 316684 4768 316736 4820
rect 345112 4768 345164 4820
rect 398748 4768 398800 4820
rect 447784 4768 447836 4820
rect 448428 4768 448480 4820
rect 576216 4768 576268 4820
rect 1676 4700 1728 4752
rect 208676 4700 208728 4752
rect 212264 4632 212316 4684
rect 314660 4700 314712 4752
rect 315948 4700 316000 4752
rect 331404 4700 331456 4752
rect 390468 4700 390520 4752
rect 422760 4700 422812 4752
rect 433248 4700 433300 4752
rect 536932 4700 536984 4752
rect 215852 4564 215904 4616
rect 307760 4632 307812 4684
rect 310520 4632 310572 4684
rect 327080 4632 327132 4684
rect 387524 4632 387576 4684
rect 415676 4632 415728 4684
rect 431868 4632 431920 4684
rect 533436 4632 533488 4684
rect 309048 4564 309100 4616
rect 309140 4564 309192 4616
rect 325700 4564 325752 4616
rect 386236 4564 386288 4616
rect 413284 4564 413336 4616
rect 430488 4564 430540 4616
rect 529848 4564 529900 4616
rect 219348 4496 219400 4548
rect 311808 4496 311860 4548
rect 314568 4496 314620 4548
rect 330024 4496 330076 4548
rect 429108 4496 429160 4548
rect 526260 4496 526312 4548
rect 222936 4428 222988 4480
rect 226524 4360 226576 4412
rect 310612 4428 310664 4480
rect 313188 4428 313240 4480
rect 328644 4428 328696 4480
rect 427728 4428 427780 4480
rect 522672 4428 522724 4480
rect 313280 4360 313332 4412
rect 317420 4360 317472 4412
rect 332784 4360 332836 4412
rect 426256 4360 426308 4412
rect 519084 4360 519136 4412
rect 201500 4292 201552 4344
rect 267280 4292 267332 4344
rect 294328 4292 294380 4344
rect 340972 4292 341024 4344
rect 424968 4292 425020 4344
rect 515588 4292 515640 4344
rect 229100 4224 229152 4276
rect 298008 4224 298060 4276
rect 341064 4224 341116 4276
rect 423588 4224 423640 4276
rect 512000 4224 512052 4276
rect 124220 4156 124272 4208
rect 125416 4156 125468 4208
rect 301412 4156 301464 4208
rect 342444 4156 342496 4208
rect 5264 4088 5316 4140
rect 10324 4088 10376 4140
rect 36176 4088 36228 4140
rect 39304 4088 39356 4140
rect 57612 4088 57664 4140
rect 249064 4088 249116 4140
rect 268108 4088 268160 4140
rect 269028 4088 269080 4140
rect 274088 4088 274140 4140
rect 274548 4088 274600 4140
rect 275284 4088 275336 4140
rect 276664 4088 276716 4140
rect 278872 4088 278924 4140
rect 279976 4088 280028 4140
rect 281264 4088 281316 4140
rect 284760 4088 284812 4140
rect 285588 4088 285640 4140
rect 291936 4088 291988 4140
rect 292488 4088 292540 4140
rect 296720 4088 296772 4140
rect 297916 4088 297968 4140
rect 307392 4088 307444 4140
rect 344284 4088 344336 4140
rect 344928 4088 344980 4140
rect 400128 4156 400180 4208
rect 451280 4156 451332 4208
rect 477500 4156 477552 4208
rect 478696 4156 478748 4208
rect 345204 4088 345256 4140
rect 345480 4088 345532 4140
rect 349804 4088 349856 4140
rect 355324 4088 355376 4140
rect 362132 4088 362184 4140
rect 362868 4088 362920 4140
rect 364524 4088 364576 4140
rect 366364 4088 366416 4140
rect 368020 4088 368072 4140
rect 368480 4088 368532 4140
rect 368572 4088 368624 4140
rect 369216 4088 369268 4140
rect 371148 4088 371200 4140
rect 374000 4088 374052 4140
rect 381544 4088 381596 4140
rect 384672 4088 384724 4140
rect 387708 4088 387760 4140
rect 417976 4088 418028 4140
rect 421564 4088 421616 4140
rect 503628 4088 503680 4140
rect 507124 4088 507176 4140
rect 521476 4088 521528 4140
rect 525064 4088 525116 4140
rect 560760 4088 560812 4140
rect 50528 4020 50580 4072
rect 247684 4020 247736 4072
rect 269304 4020 269356 4072
rect 315948 4020 316000 4072
rect 319260 4020 319312 4072
rect 344376 4020 344428 4072
rect 346676 4020 346728 4072
rect 356704 4020 356756 4072
rect 387616 4020 387668 4072
rect 46940 3952 46992 4004
rect 247224 3952 247276 4004
rect 265808 3952 265860 4004
rect 20720 3884 20772 3936
rect 42064 3884 42116 3936
rect 45744 3884 45796 3936
rect 246304 3884 246356 3936
rect 39764 3816 39816 3868
rect 244280 3816 244332 3868
rect 270500 3816 270552 3868
rect 271788 3816 271840 3868
rect 272892 3952 272944 4004
rect 317420 3952 317472 4004
rect 320456 3952 320508 4004
rect 321468 3952 321520 4004
rect 327816 3952 327868 4004
rect 330024 3952 330076 4004
rect 331128 3952 331180 4004
rect 352012 3952 352064 4004
rect 360936 3952 360988 4004
rect 362224 3952 362276 4004
rect 389088 3952 389140 4004
rect 414480 4020 414532 4072
rect 428464 4020 428516 4072
rect 510804 4020 510856 4072
rect 527824 4020 527876 4072
rect 567844 4020 567896 4072
rect 290464 3884 290516 3936
rect 293132 3884 293184 3936
rect 339684 3884 339736 3936
rect 343088 3884 343140 3936
rect 314568 3816 314620 3868
rect 316960 3816 317012 3868
rect 344192 3816 344244 3868
rect 352104 3884 352156 3936
rect 384948 3884 385000 3936
rect 388996 3884 389048 3936
rect 376024 3816 376076 3868
rect 383476 3816 383528 3868
rect 387064 3816 387116 3868
rect 393044 3816 393096 3868
rect 416872 3952 416924 4004
rect 429844 3952 429896 4004
rect 517888 3952 517940 4004
rect 529204 3952 529256 4004
rect 575020 3952 575072 4004
rect 420368 3884 420420 3936
rect 434076 3884 434128 3936
rect 525064 3884 525116 3936
rect 530584 3884 530636 3936
rect 582196 3884 582248 3936
rect 421564 3816 421616 3868
rect 436744 3816 436796 3868
rect 532240 3816 532292 3868
rect 38568 3748 38620 3800
rect 244464 3748 244516 3800
rect 262220 3748 262272 3800
rect 313188 3748 313240 3800
rect 315764 3748 315816 3800
rect 320180 3748 320232 3800
rect 325240 3748 325292 3800
rect 330484 3748 330536 3800
rect 350816 3748 350868 3800
rect 374644 3748 374696 3800
rect 381176 3748 381228 3800
rect 384856 3748 384908 3800
rect 427544 3748 427596 3800
rect 435180 3748 435232 3800
rect 539324 3748 539376 3800
rect 32680 3680 32732 3732
rect 241520 3680 241572 3732
rect 264612 3680 264664 3732
rect 276388 3680 276440 3732
rect 276480 3680 276532 3732
rect 284208 3680 284260 3732
rect 285956 3680 286008 3732
rect 328828 3680 328880 3732
rect 334624 3680 334676 3732
rect 337108 3680 337160 3732
rect 338028 3680 338080 3732
rect 339500 3680 339552 3732
rect 357624 3680 357676 3732
rect 376668 3680 376720 3732
rect 385868 3680 385920 3732
rect 386328 3680 386380 3732
rect 25504 3612 25556 3664
rect 238760 3612 238812 3664
rect 277676 3612 277728 3664
rect 287704 3612 287756 3664
rect 288348 3612 288400 3664
rect 338304 3612 338356 3664
rect 341892 3612 341944 3664
rect 358820 3612 358872 3664
rect 377404 3612 377456 3664
rect 387064 3612 387116 3664
rect 393136 3680 393188 3732
rect 428740 3680 428792 3732
rect 436836 3680 436888 3732
rect 546500 3680 546552 3732
rect 431132 3612 431184 3664
rect 440148 3612 440200 3664
rect 557172 3612 557224 3664
rect 11244 3544 11296 3596
rect 19984 3544 20036 3596
rect 24308 3544 24360 3596
rect 238852 3544 238904 3596
rect 258632 3544 258684 3596
rect 310520 3544 310572 3596
rect 312176 3544 312228 3596
rect 318800 3544 318852 3596
rect 324044 3544 324096 3596
rect 347872 3544 347924 3596
rect 349068 3544 349120 3596
rect 353760 3544 353812 3596
rect 358084 3544 358136 3596
rect 378048 3544 378100 3596
rect 389456 3544 389508 3596
rect 391756 3544 391808 3596
rect 16028 3476 16080 3528
rect 235080 3476 235132 3528
rect 14832 3408 14884 3460
rect 234712 3408 234764 3460
rect 255044 3408 255096 3460
rect 326436 3476 326488 3528
rect 19524 3340 19576 3392
rect 28264 3340 28316 3392
rect 34980 3340 35032 3392
rect 57244 3340 57296 3392
rect 64696 3340 64748 3392
rect 250444 3340 250496 3392
rect 10048 3272 10100 3324
rect 13084 3272 13136 3324
rect 29092 3272 29144 3324
rect 35164 3272 35216 3324
rect 42156 3272 42208 3324
rect 66904 3272 66956 3324
rect 70676 3272 70728 3324
rect 71688 3272 71740 3324
rect 71872 3272 71924 3324
rect 251824 3272 251876 3324
rect 43352 3204 43404 3256
rect 61384 3204 61436 3256
rect 77852 3204 77904 3256
rect 78588 3204 78640 3256
rect 81440 3204 81492 3256
rect 82728 3204 82780 3256
rect 54024 3136 54076 3188
rect 71044 3136 71096 3188
rect 75460 3136 75512 3188
rect 79324 3136 79376 3188
rect 82636 3136 82688 3188
rect 84844 3204 84896 3256
rect 84936 3204 84988 3256
rect 85488 3204 85540 3256
rect 88524 3204 88576 3256
rect 89628 3204 89680 3256
rect 253204 3204 253256 3256
rect 61200 3068 61252 3120
rect 77944 3068 77996 3120
rect 89720 3068 89772 3120
rect 254584 3136 254636 3188
rect 282460 3136 282512 3188
rect 299112 3272 299164 3324
rect 314568 3408 314620 3460
rect 321652 3340 321704 3392
rect 326252 3340 326304 3392
rect 334808 3476 334860 3528
rect 351368 3476 351420 3528
rect 351828 3476 351880 3528
rect 352564 3476 352616 3528
rect 353208 3476 353260 3528
rect 354956 3476 355008 3528
rect 355968 3476 356020 3528
rect 348056 3408 348108 3460
rect 350264 3408 350316 3460
rect 361764 3476 361816 3528
rect 363328 3476 363380 3528
rect 364248 3476 364300 3528
rect 371056 3476 371108 3528
rect 371608 3476 371660 3528
rect 373264 3476 373316 3528
rect 377588 3476 377640 3528
rect 377956 3476 378008 3528
rect 388444 3476 388496 3528
rect 391848 3476 391900 3528
rect 393228 3544 393280 3596
rect 432328 3544 432380 3596
rect 435456 3544 435508 3596
rect 442908 3544 442960 3596
rect 564348 3544 564400 3596
rect 394608 3476 394660 3528
rect 435824 3476 435876 3528
rect 438124 3476 438176 3528
rect 449164 3476 449216 3528
rect 373908 3408 373960 3460
rect 378784 3408 378836 3460
rect 380164 3408 380216 3460
rect 394240 3408 394292 3460
rect 332416 3340 332468 3392
rect 354864 3340 354916 3392
rect 390652 3340 390704 3392
rect 391480 3340 391532 3392
rect 395344 3408 395396 3460
rect 400220 3408 400272 3460
rect 439412 3408 439464 3460
rect 453672 3408 453724 3460
rect 571432 3476 571484 3528
rect 578608 3408 578660 3460
rect 405004 3340 405056 3392
rect 406108 3340 406160 3392
rect 431224 3340 431276 3392
rect 496544 3340 496596 3392
rect 500224 3340 500276 3392
rect 507216 3340 507268 3392
rect 309784 3272 309836 3324
rect 338764 3272 338816 3324
rect 349068 3272 349120 3324
rect 351184 3272 351236 3324
rect 356152 3272 356204 3324
rect 363236 3272 363288 3324
rect 365720 3272 365772 3324
rect 366916 3272 366968 3324
rect 375288 3272 375340 3324
rect 382372 3272 382424 3324
rect 383568 3272 383620 3324
rect 407304 3272 407356 3324
rect 407764 3272 407816 3324
rect 419172 3272 419224 3324
rect 420184 3272 420236 3324
rect 475108 3272 475160 3324
rect 306196 3204 306248 3256
rect 336924 3204 336976 3256
rect 338304 3204 338356 3256
rect 348424 3204 348476 3256
rect 384304 3204 384356 3256
rect 388260 3204 388312 3256
rect 408500 3204 408552 3256
rect 409144 3204 409196 3256
rect 412548 3204 412600 3256
rect 489368 3204 489420 3256
rect 502984 3204 503036 3256
rect 514392 3340 514444 3392
rect 523684 3340 523736 3392
rect 553584 3340 553636 3392
rect 520924 3272 520976 3324
rect 550088 3272 550140 3324
rect 518164 3204 518216 3256
rect 542912 3204 542964 3256
rect 289544 3136 289596 3188
rect 316592 3136 316644 3188
rect 327632 3136 327684 3188
rect 352472 3136 352524 3188
rect 382096 3136 382148 3188
rect 403716 3136 403768 3188
rect 409696 3136 409748 3188
rect 411904 3136 411956 3188
rect 94504 3068 94556 3120
rect 95148 3068 95200 3120
rect 95700 3068 95752 3120
rect 96528 3068 96580 3120
rect 98092 3068 98144 3120
rect 99196 3068 99248 3120
rect 101588 3068 101640 3120
rect 102048 3068 102100 3120
rect 102784 3068 102836 3120
rect 103428 3068 103480 3120
rect 105176 3068 105228 3120
rect 106188 3068 106240 3120
rect 106372 3068 106424 3120
rect 107476 3068 107528 3120
rect 68284 3000 68336 3052
rect 102600 3000 102652 3052
rect 79048 2932 79100 2984
rect 86132 2932 86184 2984
rect 93308 2864 93360 2916
rect 97264 2864 97316 2916
rect 96896 2796 96948 2848
rect 254676 3068 254728 3120
rect 295524 3068 295576 3120
rect 312544 3068 312596 3120
rect 103980 2864 104032 2916
rect 255964 3000 256016 3052
rect 300308 3000 300360 3052
rect 319444 3068 319496 3120
rect 313372 3000 313424 3052
rect 341524 3068 341576 3120
rect 357348 3068 357400 3120
rect 359464 3068 359516 3120
rect 382188 3068 382240 3120
rect 401324 3068 401376 3120
rect 405096 3068 405148 3120
rect 412088 3068 412140 3120
rect 417424 3136 417476 3188
rect 467932 3136 467984 3188
rect 496084 3136 496136 3188
rect 500132 3136 500184 3188
rect 514024 3136 514076 3188
rect 535736 3136 535788 3188
rect 460848 3068 460900 3120
rect 511264 3068 511316 3120
rect 528652 3068 528704 3120
rect 345756 3000 345808 3052
rect 380808 3000 380860 3052
rect 397828 3000 397880 3052
rect 402612 3000 402664 3052
rect 425152 3000 425204 3052
rect 433984 3000 434036 3052
rect 481088 3000 481140 3052
rect 112352 2932 112404 2984
rect 113088 2932 113140 2984
rect 113548 2932 113600 2984
rect 114468 2932 114520 2984
rect 115940 2932 115992 2984
rect 116952 2932 117004 2984
rect 119436 2932 119488 2984
rect 119988 2932 120040 2984
rect 120632 2932 120684 2984
rect 121368 2932 121420 2984
rect 111156 2864 111208 2916
rect 257344 2932 257396 2984
rect 271696 2932 271748 2984
rect 273904 2932 273956 2984
rect 105544 2796 105596 2848
rect 114744 2796 114796 2848
rect 258724 2864 258776 2916
rect 302608 2864 302660 2916
rect 303528 2864 303580 2916
rect 303804 2932 303856 2984
rect 322204 2932 322256 2984
rect 309140 2864 309192 2916
rect 310980 2864 311032 2916
rect 326160 2932 326212 2984
rect 334624 2932 334676 2984
rect 334716 2932 334768 2984
rect 356428 2932 356480 2984
rect 381636 2932 381688 2984
rect 395436 2932 395488 2984
rect 395988 2932 396040 2984
rect 410524 2932 410576 2984
rect 322848 2864 322900 2916
rect 327724 2864 327776 2916
rect 331220 2864 331272 2916
rect 345664 2864 345716 2916
rect 392584 2864 392636 2916
rect 396632 2864 396684 2916
rect 399484 2864 399536 2916
rect 410892 2864 410944 2916
rect 412548 2932 412600 2984
rect 446588 2932 446640 2984
rect 482284 2932 482336 2984
rect 442264 2864 442316 2916
rect 121828 2796 121880 2848
rect 258816 2796 258868 2848
rect 308588 2796 308640 2848
rect 316684 2796 316736 2848
rect 318064 2796 318116 2848
rect 326436 2796 326488 2848
rect 335912 2796 335964 2848
rect 356520 2796 356572 2848
rect 393964 2796 394016 2848
rect 404912 2796 404964 2848
rect 406384 2796 406436 2848
rect 443000 2796 443052 2848
rect 445668 2796 445720 2848
rect 473912 2796 473964 2848
rect 23112 552 23164 604
rect 23388 552 23440 604
rect 148048 552 148100 604
rect 148968 552 149020 604
rect 151544 552 151596 604
rect 151728 552 151780 604
rect 153936 552 153988 604
rect 154488 552 154540 604
rect 155132 552 155184 604
rect 155868 552 155920 604
rect 157524 552 157576 604
rect 158628 552 158680 604
rect 161112 552 161164 604
rect 161388 552 161440 604
rect 171784 552 171836 604
rect 172428 552 172480 604
rect 172980 552 173032 604
rect 173808 552 173860 604
rect 178960 552 179012 604
rect 179328 552 179380 604
rect 180156 552 180208 604
rect 180708 552 180760 604
rect 182548 552 182600 604
rect 183468 552 183520 604
rect 183744 552 183796 604
rect 184756 552 184808 604
rect 189632 552 189684 604
rect 190368 552 190420 604
rect 190828 552 190880 604
rect 191748 552 191800 604
rect 196808 552 196860 604
rect 197268 552 197320 604
rect 198004 552 198056 604
rect 198648 552 198700 604
rect 217048 552 217100 604
rect 217968 552 218020 604
rect 220544 552 220596 604
rect 220728 552 220780 604
rect 224132 552 224184 604
rect 224868 552 224920 604
rect 358544 552 358596 604
rect 358728 552 358780 604
rect 379612 552 379664 604
rect 379980 552 380032 604
rect 492680 552 492732 604
rect 492956 552 493008 604
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 700369 8156 703520
rect 8114 700360 8170 700369
rect 24320 700330 24348 703520
rect 40512 700398 40540 703520
rect 72988 700466 73016 703520
rect 89180 700534 89208 703520
rect 105464 700602 105492 703520
rect 137848 700738 137876 703520
rect 154132 700874 154160 703520
rect 170324 700942 170352 703520
rect 170312 700936 170364 700942
rect 170312 700878 170364 700884
rect 154120 700868 154172 700874
rect 154120 700810 154172 700816
rect 137836 700732 137888 700738
rect 137836 700674 137888 700680
rect 105452 700596 105504 700602
rect 105452 700538 105504 700544
rect 89168 700528 89220 700534
rect 89168 700470 89220 700476
rect 72976 700460 73028 700466
rect 72976 700402 73028 700408
rect 40500 700392 40552 700398
rect 40500 700334 40552 700340
rect 8114 700295 8170 700304
rect 24308 700324 24360 700330
rect 24308 700266 24360 700272
rect 202800 700262 202828 703520
rect 202788 700256 202840 700262
rect 202788 700198 202840 700204
rect 218992 700126 219020 703520
rect 218980 700120 219032 700126
rect 218980 700062 219032 700068
rect 235184 700058 235212 703520
rect 235172 700052 235224 700058
rect 235172 699994 235224 700000
rect 267660 699922 267688 703520
rect 267648 699916 267700 699922
rect 267648 699858 267700 699864
rect 283852 699786 283880 703520
rect 283840 699780 283892 699786
rect 283840 699722 283892 699728
rect 300136 699718 300164 703520
rect 328368 701004 328420 701010
rect 328368 700946 328420 700952
rect 320088 700800 320140 700806
rect 320088 700742 320140 700748
rect 300124 699712 300176 699718
rect 300124 699654 300176 699660
rect 300768 699712 300820 699718
rect 300768 699654 300820 699660
rect 3514 682272 3570 682281
rect 3514 682207 3570 682216
rect 3528 681766 3556 682207
rect 3516 681760 3568 681766
rect 3516 681702 3568 681708
rect 3422 667992 3478 668001
rect 3422 667927 3424 667936
rect 3476 667927 3478 667936
rect 3424 667898 3476 667904
rect 3054 653576 3110 653585
rect 3054 653511 3110 653520
rect 3068 652798 3096 653511
rect 3056 652792 3108 652798
rect 3056 652734 3108 652740
rect 3422 624880 3478 624889
rect 3422 624815 3478 624824
rect 3436 623830 3464 624815
rect 3424 623824 3476 623830
rect 3424 623766 3476 623772
rect 3422 610464 3478 610473
rect 3422 610399 3478 610408
rect 3436 610026 3464 610399
rect 3424 610020 3476 610026
rect 3424 609962 3476 609968
rect 3238 596048 3294 596057
rect 3238 595983 3294 595992
rect 3252 594862 3280 595983
rect 3240 594856 3292 594862
rect 3240 594798 3292 594804
rect 300676 579692 300728 579698
rect 300676 579634 300728 579640
rect 3422 567352 3478 567361
rect 3422 567287 3478 567296
rect 3436 567254 3464 567287
rect 3424 567248 3476 567254
rect 3424 567190 3476 567196
rect 289820 563032 289872 563038
rect 249982 563000 250038 563009
rect 249982 562935 250038 562944
rect 288622 563000 288678 563009
rect 289820 562974 289872 562980
rect 288622 562935 288678 562944
rect 4158 562728 4214 562737
rect 4158 562663 4214 562672
rect 3974 562592 4030 562601
rect 3974 562527 4030 562536
rect 3056 562352 3108 562358
rect 3056 562294 3108 562300
rect 3790 562320 3846 562329
rect 2962 558240 3018 558249
rect 2962 558175 3018 558184
rect 2780 553104 2832 553110
rect 2778 553072 2780 553081
rect 2832 553072 2834 553081
rect 2778 553007 2834 553016
rect 2976 538665 3004 558175
rect 2962 538656 3018 538665
rect 2962 538591 3018 538600
rect 3068 509969 3096 562294
rect 3790 562255 3846 562264
rect 3148 562216 3200 562222
rect 3148 562158 3200 562164
rect 3054 509960 3110 509969
rect 3054 509895 3110 509904
rect 3056 495576 3108 495582
rect 3054 495544 3056 495553
rect 3108 495544 3110 495553
rect 3054 495479 3110 495488
rect 3056 481160 3108 481166
rect 3054 481128 3056 481137
rect 3108 481128 3110 481137
rect 3054 481063 3110 481072
rect 3160 452441 3188 562158
rect 3240 562012 3292 562018
rect 3240 561954 3292 561960
rect 3146 452432 3202 452441
rect 3146 452367 3202 452376
rect 3148 438728 3200 438734
rect 3148 438670 3200 438676
rect 3160 438025 3188 438670
rect 3146 438016 3202 438025
rect 3146 437951 3202 437960
rect 2780 424720 2832 424726
rect 2780 424662 2832 424668
rect 2792 423745 2820 424662
rect 2778 423736 2834 423745
rect 2778 423671 2834 423680
rect 3252 395049 3280 561954
rect 3332 561808 3384 561814
rect 3332 561750 3384 561756
rect 3606 561776 3662 561785
rect 3238 395040 3294 395049
rect 3238 394975 3294 394984
rect 3148 380656 3200 380662
rect 3146 380624 3148 380633
rect 3200 380624 3202 380633
rect 3146 380559 3202 380568
rect 2780 366988 2832 366994
rect 2780 366930 2832 366936
rect 2792 366217 2820 366930
rect 2778 366208 2834 366217
rect 2778 366143 2834 366152
rect 3344 323105 3372 561750
rect 3606 561711 3662 561720
rect 3516 559156 3568 559162
rect 3516 559098 3568 559104
rect 3422 559056 3478 559065
rect 3422 558991 3478 559000
rect 3330 323096 3386 323105
rect 3330 323031 3386 323040
rect 2780 295248 2832 295254
rect 2780 295190 2832 295196
rect 2792 294409 2820 295190
rect 2778 294400 2834 294409
rect 2778 294335 2834 294344
rect 3148 280152 3200 280158
rect 3146 280120 3148 280129
rect 3200 280120 3202 280129
rect 3146 280055 3202 280064
rect 3146 252512 3202 252521
rect 3146 252447 3202 252456
rect 3160 251297 3188 252447
rect 3146 251288 3202 251297
rect 3146 251223 3202 251232
rect 2780 208208 2832 208214
rect 2778 208176 2780 208185
rect 2832 208176 2834 208185
rect 2778 208111 2834 208120
rect 2780 179852 2832 179858
rect 2780 179794 2832 179800
rect 2792 179489 2820 179794
rect 2778 179480 2834 179489
rect 2778 179415 2834 179424
rect 2780 165504 2832 165510
rect 2780 165446 2832 165452
rect 2792 165073 2820 165446
rect 2778 165064 2834 165073
rect 2778 164999 2834 165008
rect 2780 136400 2832 136406
rect 2778 136368 2780 136377
rect 2832 136368 2834 136377
rect 2778 136303 2834 136312
rect 2780 122120 2832 122126
rect 2778 122088 2780 122097
rect 2832 122088 2834 122097
rect 2778 122023 2834 122032
rect 2780 79484 2832 79490
rect 2780 79426 2832 79432
rect 2792 78985 2820 79426
rect 2778 78976 2834 78985
rect 2778 78911 2834 78920
rect 3436 64569 3464 558991
rect 3528 93265 3556 559098
rect 3620 107681 3648 561711
rect 3700 559360 3752 559366
rect 3700 559302 3752 559308
rect 3712 150793 3740 559302
rect 3804 193905 3832 562255
rect 3884 559768 3936 559774
rect 3884 559710 3936 559716
rect 3896 222601 3924 559710
rect 3988 237017 4016 562527
rect 4068 560992 4120 560998
rect 4068 560934 4120 560940
rect 4080 265713 4108 560934
rect 4066 265704 4122 265713
rect 4066 265639 4122 265648
rect 3974 237008 4030 237017
rect 3974 236943 4030 236952
rect 3882 222592 3938 222601
rect 3882 222527 3938 222536
rect 3790 193896 3846 193905
rect 3790 193831 3846 193840
rect 3698 150784 3754 150793
rect 3698 150719 3754 150728
rect 3606 107672 3662 107681
rect 3606 107607 3662 107616
rect 3514 93256 3570 93265
rect 3514 93191 3570 93200
rect 3422 64560 3478 64569
rect 3422 64495 3478 64504
rect 4066 50144 4122 50153
rect 4172 50130 4200 562663
rect 242254 562592 242310 562601
rect 242254 562527 242310 562536
rect 248050 562592 248106 562601
rect 248050 562527 248106 562536
rect 6552 562420 6604 562426
rect 6552 562362 6604 562368
rect 5354 562320 5410 562329
rect 5354 562255 5410 562264
rect 5078 562184 5134 562193
rect 5078 562119 5134 562128
rect 4894 561912 4950 561921
rect 4894 561847 4950 561856
rect 4804 560380 4856 560386
rect 4804 560322 4856 560328
rect 4816 122126 4844 560322
rect 4908 136406 4936 561847
rect 4988 560448 5040 560454
rect 4988 560390 5040 560396
rect 5000 165510 5028 560390
rect 5092 179858 5120 562119
rect 5368 562057 5396 562255
rect 5448 562148 5500 562154
rect 5448 562090 5500 562096
rect 5354 562048 5410 562057
rect 5354 561983 5410 561992
rect 5356 561944 5408 561950
rect 5356 561886 5408 561892
rect 5264 560584 5316 560590
rect 5264 560526 5316 560532
rect 5172 560516 5224 560522
rect 5172 560458 5224 560464
rect 5184 208214 5212 560458
rect 5276 295254 5304 560526
rect 5368 366994 5396 561886
rect 5460 424726 5488 562090
rect 6460 562080 6512 562086
rect 6460 562022 6512 562028
rect 6368 561876 6420 561882
rect 6368 561818 6420 561824
rect 6276 561740 6328 561746
rect 6276 561682 6328 561688
rect 6184 560312 6236 560318
rect 6184 560254 6236 560260
rect 5540 559428 5592 559434
rect 5540 559370 5592 559376
rect 5552 553110 5580 559370
rect 5540 553104 5592 553110
rect 5540 553046 5592 553052
rect 5448 424720 5500 424726
rect 5448 424662 5500 424668
rect 5356 366988 5408 366994
rect 5356 366930 5408 366936
rect 5264 295248 5316 295254
rect 5264 295190 5316 295196
rect 5172 208208 5224 208214
rect 5172 208150 5224 208156
rect 5080 179852 5132 179858
rect 5080 179794 5132 179800
rect 4988 165504 5040 165510
rect 4988 165446 5040 165452
rect 4896 136400 4948 136406
rect 4896 136342 4948 136348
rect 4804 122120 4856 122126
rect 4804 122062 4856 122068
rect 6196 79490 6224 560254
rect 6288 280158 6316 561682
rect 6380 380662 6408 561818
rect 6472 438734 6500 562022
rect 6564 481166 6592 562362
rect 6644 562284 6696 562290
rect 6644 562226 6696 562232
rect 6656 495582 6684 562226
rect 242268 559980 242296 562527
rect 243818 562456 243874 562465
rect 243818 562391 243874 562400
rect 243832 559994 243860 562391
rect 243832 559966 244214 559994
rect 248064 559980 248092 562527
rect 249996 559980 250024 562935
rect 255780 562896 255832 562902
rect 255780 562838 255832 562844
rect 286968 562896 287020 562902
rect 286968 562838 287020 562844
rect 253846 560416 253902 560425
rect 253846 560351 253902 560360
rect 253860 559980 253888 560351
rect 255792 559980 255820 562838
rect 284760 562828 284812 562834
rect 284760 562770 284812 562776
rect 280896 562760 280948 562766
rect 280896 562702 280948 562708
rect 278964 562692 279016 562698
rect 278964 562634 279016 562640
rect 261576 562624 261628 562630
rect 261576 562566 261628 562572
rect 278780 562624 278832 562630
rect 278780 562566 278832 562572
rect 259644 562488 259696 562494
rect 259644 562430 259696 562436
rect 259656 559980 259684 562430
rect 261588 559980 261616 562566
rect 273168 562556 273220 562562
rect 273168 562498 273220 562504
rect 271236 560720 271288 560726
rect 271236 560662 271288 560668
rect 269672 560040 269724 560046
rect 267398 559978 267688 559994
rect 269330 559988 269672 559994
rect 269330 559982 269724 559988
rect 267398 559972 267700 559978
rect 267398 559966 267648 559972
rect 269330 559966 269712 559982
rect 271248 559980 271276 560662
rect 273180 559980 273208 562498
rect 277032 560788 277084 560794
rect 277032 560730 277084 560736
rect 275100 560108 275152 560114
rect 275100 560050 275152 560056
rect 275112 559980 275140 560050
rect 277044 559980 277072 560730
rect 278792 560182 278820 562566
rect 278780 560176 278832 560182
rect 278780 560118 278832 560124
rect 278976 559980 279004 562634
rect 280908 559980 280936 562702
rect 282828 560856 282880 560862
rect 282828 560798 282880 560804
rect 282840 559980 282868 560798
rect 284772 559980 284800 562770
rect 286692 562624 286744 562630
rect 286692 562566 286744 562572
rect 286704 559980 286732 562566
rect 286980 560658 287008 562838
rect 286968 560652 287020 560658
rect 286968 560594 287020 560600
rect 288636 559980 288664 562935
rect 289832 560998 289860 562974
rect 298284 562964 298336 562970
rect 298284 562906 298336 562912
rect 292488 562896 292540 562902
rect 292488 562838 292540 562844
rect 289820 560992 289872 560998
rect 289820 560934 289872 560940
rect 290556 560924 290608 560930
rect 290556 560866 290608 560872
rect 290568 559980 290596 560866
rect 292500 559980 292528 562838
rect 296352 560992 296404 560998
rect 296352 560934 296404 560940
rect 294420 560652 294472 560658
rect 294420 560594 294472 560600
rect 294432 559980 294460 560594
rect 296364 559980 296392 560934
rect 298296 559980 298324 562906
rect 300688 559994 300716 579634
rect 300780 563922 300808 699654
rect 314568 696992 314620 696998
rect 314568 696934 314620 696940
rect 311808 673532 311860 673538
rect 311808 673474 311860 673480
rect 309048 650072 309100 650078
rect 309048 650014 309100 650020
rect 306288 626612 306340 626618
rect 306288 626554 306340 626560
rect 302148 603152 302200 603158
rect 302148 603094 302200 603100
rect 300768 563916 300820 563922
rect 300768 563858 300820 563864
rect 300242 559966 300716 559994
rect 302160 559980 302188 603094
rect 304908 592068 304960 592074
rect 304908 592010 304960 592016
rect 304920 560266 304948 592010
rect 304552 560238 304948 560266
rect 304552 559994 304580 560238
rect 306300 559994 306328 626554
rect 309060 565146 309088 650014
rect 310428 638988 310480 638994
rect 310428 638930 310480 638936
rect 310440 565146 310468 638930
rect 311820 565146 311848 673474
rect 314580 565146 314608 696934
rect 315948 685908 316000 685914
rect 315948 685850 316000 685856
rect 315960 565146 315988 685850
rect 307760 565140 307812 565146
rect 307760 565082 307812 565088
rect 309048 565140 309100 565146
rect 309048 565082 309100 565088
rect 309140 565140 309192 565146
rect 309140 565082 309192 565088
rect 310428 565140 310480 565146
rect 310428 565082 310480 565088
rect 310520 565140 310572 565146
rect 310520 565082 310572 565088
rect 311808 565140 311860 565146
rect 311808 565082 311860 565088
rect 313280 565140 313332 565146
rect 313280 565082 313332 565088
rect 314568 565140 314620 565146
rect 314568 565082 314620 565088
rect 314660 565140 314712 565146
rect 314660 565082 314712 565088
rect 315948 565140 316000 565146
rect 315948 565082 316000 565088
rect 304106 559966 304580 559994
rect 305946 559966 306328 559994
rect 307772 559994 307800 565082
rect 309152 560130 309180 565082
rect 310532 562970 310560 565082
rect 310520 562964 310572 562970
rect 310520 562906 310572 562912
rect 311716 562964 311768 562970
rect 311716 562906 311768 562912
rect 309152 560102 309456 560130
rect 309428 559994 309456 560102
rect 307772 559966 307878 559994
rect 309428 559966 309810 559994
rect 311728 559980 311756 562906
rect 313292 559994 313320 565082
rect 314672 560130 314700 565082
rect 317512 563712 317564 563718
rect 317512 563654 317564 563660
rect 314672 560102 315252 560130
rect 315224 559994 315252 560102
rect 313292 559966 313674 559994
rect 315224 559966 315606 559994
rect 317524 559980 317552 563654
rect 320100 560130 320128 700742
rect 321468 700664 321520 700670
rect 321468 700606 321520 700612
rect 319732 560102 320128 560130
rect 319732 559994 319760 560102
rect 321480 559994 321508 700606
rect 325608 700188 325660 700194
rect 325608 700130 325660 700136
rect 323308 563780 323360 563786
rect 323308 563722 323360 563728
rect 319470 559966 319760 559994
rect 321402 559966 321508 559994
rect 323320 559980 323348 563722
rect 325620 559994 325648 700130
rect 328380 565146 328408 700946
rect 331128 699848 331180 699854
rect 331128 699790 331180 699796
rect 331140 565146 331168 699790
rect 332520 699718 332548 703520
rect 347872 700256 347924 700262
rect 347872 700198 347924 700204
rect 348424 700256 348476 700262
rect 348424 700198 348476 700204
rect 346400 700052 346452 700058
rect 346400 699994 346452 700000
rect 333888 699984 333940 699990
rect 333888 699926 333940 699932
rect 332508 699712 332560 699718
rect 332508 699654 332560 699660
rect 333900 565146 333928 699926
rect 342260 699916 342312 699922
rect 342260 699858 342312 699864
rect 336740 699712 336792 699718
rect 336740 699654 336792 699660
rect 339408 699712 339460 699718
rect 339408 699654 339460 699660
rect 327080 565140 327132 565146
rect 327080 565082 327132 565088
rect 328368 565140 328420 565146
rect 328368 565082 328420 565088
rect 329840 565140 329892 565146
rect 329840 565082 329892 565088
rect 331128 565140 331180 565146
rect 331128 565082 331180 565088
rect 332600 565140 332652 565146
rect 332600 565082 332652 565088
rect 333888 565140 333940 565146
rect 333888 565082 333940 565088
rect 325698 560960 325754 560969
rect 325698 560895 325754 560904
rect 325712 560697 325740 560895
rect 325698 560688 325754 560697
rect 325698 560623 325754 560632
rect 325266 559966 325648 559994
rect 327092 559994 327120 565082
rect 328460 563848 328512 563854
rect 328460 563790 328512 563796
rect 328472 560130 328500 563790
rect 329852 560130 329880 565082
rect 328472 560102 328868 560130
rect 329852 560102 330708 560130
rect 328840 559994 328868 560102
rect 330680 559994 330708 560102
rect 332612 559994 332640 565082
rect 333980 563984 334032 563990
rect 333980 563926 334032 563932
rect 333992 560130 334020 563926
rect 333992 560102 334572 560130
rect 334544 559994 334572 560102
rect 336752 559994 336780 699654
rect 339420 560130 339448 699654
rect 340696 563916 340748 563922
rect 340696 563858 340748 563864
rect 339052 560102 339448 560130
rect 339052 559994 339080 560102
rect 327092 559966 327198 559994
rect 328840 559966 329130 559994
rect 330680 559966 331062 559994
rect 332612 559966 332994 559994
rect 334544 559966 334926 559994
rect 336752 559966 336858 559994
rect 338790 559966 339080 559994
rect 340708 559980 340736 563858
rect 342272 559994 342300 699858
rect 343640 699780 343692 699786
rect 343640 699722 343692 699728
rect 343652 560266 343680 699722
rect 345018 560824 345074 560833
rect 345018 560759 345074 560768
rect 344926 560688 344982 560697
rect 344926 560623 344982 560632
rect 344940 560538 344968 560623
rect 345032 560538 345060 560759
rect 344940 560510 345060 560538
rect 343652 560238 344232 560266
rect 344204 559994 344232 560238
rect 346412 559994 346440 699994
rect 347884 559994 347912 700198
rect 348436 563990 348464 700198
rect 348804 699718 348832 703520
rect 351920 700936 351972 700942
rect 351920 700878 351972 700884
rect 349160 700120 349212 700126
rect 349160 700062 349212 700068
rect 348792 699712 348844 699718
rect 348792 699654 348844 699660
rect 348424 563984 348476 563990
rect 348424 563926 348476 563932
rect 349172 560266 349200 700062
rect 349172 560238 349936 560266
rect 349908 559994 349936 560238
rect 351932 559994 351960 700878
rect 356060 700868 356112 700874
rect 356060 700810 356112 700816
rect 353300 700732 353352 700738
rect 353300 700674 353352 700680
rect 353312 560130 353340 700674
rect 353312 560102 353892 560130
rect 353864 559994 353892 560102
rect 356072 559994 356100 700810
rect 357440 700596 357492 700602
rect 357440 700538 357492 700544
rect 357346 560824 357402 560833
rect 357346 560759 357402 560768
rect 357360 560561 357388 560759
rect 357346 560552 357402 560561
rect 357346 560487 357402 560496
rect 357452 560130 357480 700538
rect 361580 700528 361632 700534
rect 361580 700470 361632 700476
rect 358820 700460 358872 700466
rect 358820 700402 358872 700408
rect 358832 560130 358860 700402
rect 357452 560102 357756 560130
rect 358832 560102 359780 560130
rect 357728 559994 357756 560102
rect 359752 559994 359780 560102
rect 361592 559994 361620 700470
rect 362960 700392 363012 700398
rect 362960 700334 363012 700340
rect 362972 560266 363000 700334
rect 364996 700262 365024 703520
rect 365718 700360 365774 700369
rect 365718 700295 365774 700304
rect 367100 700324 367152 700330
rect 364984 700256 365036 700262
rect 364984 700198 365036 700204
rect 362972 560238 363552 560266
rect 363524 559994 363552 560238
rect 365732 559994 365760 700295
rect 367100 700266 367152 700272
rect 367006 560824 367062 560833
rect 367006 560759 367062 560768
rect 367020 560561 367048 560759
rect 367006 560552 367062 560561
rect 367006 560487 367062 560496
rect 367112 560130 367140 700266
rect 397472 699854 397500 703520
rect 413664 699990 413692 703520
rect 413652 699984 413704 699990
rect 413652 699926 413704 699932
rect 397460 699848 397512 699854
rect 397460 699790 397512 699796
rect 429856 688634 429884 703520
rect 462332 700194 462360 703520
rect 478524 701010 478552 703520
rect 494808 703474 494836 703520
rect 494808 703446 494928 703474
rect 478512 701004 478564 701010
rect 478512 700946 478564 700952
rect 462320 700188 462372 700194
rect 462320 700130 462372 700136
rect 429384 688628 429436 688634
rect 429384 688570 429436 688576
rect 429844 688628 429896 688634
rect 429844 688570 429896 688576
rect 429396 685930 429424 688570
rect 494900 686089 494928 703446
rect 527192 700806 527220 703520
rect 527180 700800 527232 700806
rect 527180 700742 527232 700748
rect 543476 700670 543504 703520
rect 543464 700664 543516 700670
rect 543464 700606 543516 700612
rect 559668 688634 559696 703520
rect 580170 698048 580226 698057
rect 580170 697983 580226 697992
rect 580184 696998 580212 697983
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 559104 688628 559156 688634
rect 559104 688570 559156 688576
rect 559656 688628 559708 688634
rect 559656 688570 559708 688576
rect 494886 686080 494942 686089
rect 494886 686015 494942 686024
rect 429304 685902 429424 685930
rect 494242 685944 494298 685953
rect 429304 684486 429332 685902
rect 559116 685930 559144 688570
rect 580170 686352 580226 686361
rect 580170 686287 580226 686296
rect 494242 685879 494298 685888
rect 559024 685902 559144 685930
rect 580184 685914 580212 686287
rect 580172 685908 580224 685914
rect 429292 684480 429344 684486
rect 429292 684422 429344 684428
rect 368480 681760 368532 681766
rect 368480 681702 368532 681708
rect 368492 560266 368520 681702
rect 494256 678994 494284 685879
rect 559024 684486 559052 685902
rect 580172 685850 580224 685856
rect 559012 684480 559064 684486
rect 559012 684422 559064 684428
rect 494072 678966 494284 678994
rect 494072 676190 494100 678966
rect 494060 676184 494112 676190
rect 494060 676126 494112 676132
rect 580170 674656 580226 674665
rect 580170 674591 580226 674600
rect 580184 673538 580212 674591
rect 580172 673532 580224 673538
rect 580172 673474 580224 673480
rect 372620 667956 372672 667962
rect 372620 667898 372672 667904
rect 371240 652792 371292 652798
rect 371240 652734 371292 652740
rect 368492 560238 369256 560266
rect 367112 560102 367416 560130
rect 367388 559994 367416 560102
rect 369228 559994 369256 560238
rect 371252 559994 371280 652734
rect 372250 560144 372306 560153
rect 372632 560130 372660 667898
rect 429660 666596 429712 666602
rect 429660 666538 429712 666544
rect 494152 666596 494204 666602
rect 494152 666538 494204 666544
rect 559380 666596 559432 666602
rect 559380 666538 559432 666544
rect 429672 659682 429700 666538
rect 429488 659654 429700 659682
rect 494164 659682 494192 666538
rect 559392 659682 559420 666538
rect 494164 659654 494284 659682
rect 429488 647290 429516 659654
rect 494256 654158 494284 659654
rect 559208 659654 559420 659682
rect 494060 654152 494112 654158
rect 494060 654094 494112 654100
rect 494244 654152 494296 654158
rect 494244 654094 494296 654100
rect 429384 647284 429436 647290
rect 429384 647226 429436 647232
rect 429476 647284 429528 647290
rect 429476 647226 429528 647232
rect 429396 640422 429424 647226
rect 494072 644450 494100 654094
rect 559208 647290 559236 659654
rect 580170 651128 580226 651137
rect 580170 651063 580226 651072
rect 580184 650078 580212 651063
rect 580172 650072 580224 650078
rect 580172 650014 580224 650020
rect 559104 647284 559156 647290
rect 559104 647226 559156 647232
rect 559196 647284 559248 647290
rect 559196 647226 559248 647232
rect 494072 644422 494284 644450
rect 429384 640416 429436 640422
rect 429384 640358 429436 640364
rect 429476 640416 429528 640422
rect 429476 640358 429528 640364
rect 429488 630698 429516 640358
rect 494256 634846 494284 644422
rect 559116 640422 559144 647226
rect 559104 640416 559156 640422
rect 559104 640358 559156 640364
rect 559196 640416 559248 640422
rect 559196 640358 559248 640364
rect 494060 634840 494112 634846
rect 494060 634782 494112 634788
rect 494244 634840 494296 634846
rect 494244 634782 494296 634788
rect 429292 630692 429344 630698
rect 429292 630634 429344 630640
rect 429476 630692 429528 630698
rect 429476 630634 429528 630640
rect 429304 630578 429332 630634
rect 429304 630550 429424 630578
rect 375380 623824 375432 623830
rect 375380 623766 375432 623772
rect 372632 560102 373212 560130
rect 372250 560079 372306 560088
rect 342272 559966 342654 559994
rect 344204 559966 344586 559994
rect 346412 559966 346518 559994
rect 347884 559966 348450 559994
rect 349908 559966 350382 559994
rect 351932 559966 352314 559994
rect 353864 559966 354246 559994
rect 356072 559966 356178 559994
rect 357728 559966 358110 559994
rect 359752 559966 360042 559994
rect 361592 559966 361974 559994
rect 363524 559966 363906 559994
rect 365732 559966 365838 559994
rect 367388 559966 367770 559994
rect 369228 559966 369702 559994
rect 371252 559966 371634 559994
rect 267648 559914 267700 559920
rect 372264 559910 372292 560079
rect 373184 559994 373212 560102
rect 375392 559994 375420 623766
rect 429396 621058 429424 630550
rect 494072 625138 494100 634782
rect 559208 630698 559236 640358
rect 580170 639432 580226 639441
rect 580170 639367 580226 639376
rect 580184 638994 580212 639367
rect 580172 638988 580224 638994
rect 580172 638930 580224 638936
rect 559012 630692 559064 630698
rect 559012 630634 559064 630640
rect 559196 630692 559248 630698
rect 559196 630634 559248 630640
rect 559024 630578 559052 630634
rect 559024 630550 559144 630578
rect 494072 625110 494284 625138
rect 429396 621030 429516 621058
rect 429488 611386 429516 621030
rect 494256 615534 494284 625110
rect 559116 621058 559144 630550
rect 580170 627736 580226 627745
rect 580170 627671 580226 627680
rect 580184 626618 580212 627671
rect 580172 626612 580224 626618
rect 580172 626554 580224 626560
rect 559116 621030 559236 621058
rect 494060 615528 494112 615534
rect 494060 615470 494112 615476
rect 494244 615528 494296 615534
rect 494244 615470 494296 615476
rect 429292 611380 429344 611386
rect 429292 611322 429344 611328
rect 429476 611380 429528 611386
rect 429476 611322 429528 611328
rect 429304 611266 429332 611322
rect 429304 611238 429424 611266
rect 378140 610020 378192 610026
rect 378140 609962 378192 609968
rect 376760 594856 376812 594862
rect 376760 594798 376812 594804
rect 376772 560130 376800 594798
rect 378152 560130 378180 609962
rect 429396 608598 429424 611238
rect 429384 608592 429436 608598
rect 429384 608534 429436 608540
rect 494072 605826 494100 615470
rect 559208 611386 559236 621030
rect 559012 611380 559064 611386
rect 559012 611322 559064 611328
rect 559196 611380 559248 611386
rect 559196 611322 559248 611328
rect 559024 611266 559052 611322
rect 559024 611238 559144 611266
rect 559116 608598 559144 611238
rect 559104 608592 559156 608598
rect 559104 608534 559156 608540
rect 494072 605798 494284 605826
rect 429568 601724 429620 601730
rect 429568 601666 429620 601672
rect 429580 598942 429608 601666
rect 429568 598936 429620 598942
rect 429568 598878 429620 598884
rect 494256 596222 494284 605798
rect 580170 604208 580226 604217
rect 580170 604143 580226 604152
rect 580184 603158 580212 604143
rect 580172 603152 580224 603158
rect 580172 603094 580224 603100
rect 559288 601724 559340 601730
rect 559288 601666 559340 601672
rect 559300 598942 559328 601666
rect 559288 598936 559340 598942
rect 559288 598878 559340 598884
rect 494060 596216 494112 596222
rect 494244 596216 494296 596222
rect 494112 596164 494192 596170
rect 494060 596158 494192 596164
rect 494244 596158 494296 596164
rect 494072 596142 494192 596158
rect 494164 596034 494192 596142
rect 494164 596006 494284 596034
rect 494256 591954 494284 596006
rect 580170 592512 580226 592521
rect 580170 592447 580226 592456
rect 580184 592074 580212 592447
rect 580172 592068 580224 592074
rect 580172 592010 580224 592016
rect 494164 591926 494284 591954
rect 429660 589348 429712 589354
rect 429660 589290 429712 589296
rect 429672 584474 429700 589290
rect 429488 584446 429700 584474
rect 429488 579714 429516 584446
rect 494164 579714 494192 591926
rect 559380 589348 559432 589354
rect 559380 589290 559432 589296
rect 559392 584474 559420 589290
rect 429488 579686 429608 579714
rect 429580 579630 429608 579686
rect 494072 579686 494192 579714
rect 559208 584446 559420 584474
rect 559208 579714 559236 584446
rect 580170 580816 580226 580825
rect 580170 580751 580226 580760
rect 559208 579686 559328 579714
rect 580184 579698 580212 580751
rect 494072 579630 494100 579686
rect 559300 579630 559328 579686
rect 580172 579692 580224 579698
rect 580172 579634 580224 579640
rect 429568 579624 429620 579630
rect 429568 579566 429620 579572
rect 494060 579624 494112 579630
rect 494060 579566 494112 579572
rect 559288 579624 559340 579630
rect 559288 579566 559340 579572
rect 429476 569968 429528 569974
rect 429476 569910 429528 569916
rect 494244 569968 494296 569974
rect 494244 569910 494296 569916
rect 559380 569968 559432 569974
rect 559380 569910 559432 569916
rect 380900 567248 380952 567254
rect 380900 567190 380952 567196
rect 376772 560102 377076 560130
rect 378152 560102 378916 560130
rect 377048 559994 377076 560102
rect 378888 559994 378916 560102
rect 380912 559994 380940 567190
rect 429488 563854 429516 569910
rect 429476 563848 429528 563854
rect 429476 563790 429528 563796
rect 494256 563786 494284 569910
rect 494244 563780 494296 563786
rect 494244 563722 494296 563728
rect 559392 563718 559420 569910
rect 559380 563712 559432 563718
rect 559380 563654 559432 563660
rect 412088 563032 412140 563038
rect 412088 562974 412140 562980
rect 404358 562864 404414 562873
rect 404358 562799 404414 562808
rect 388904 562420 388956 562426
rect 388904 562362 388956 562368
rect 386972 562352 387024 562358
rect 386972 562294 387024 562300
rect 386234 560960 386290 560969
rect 386234 560895 386290 560904
rect 386248 560561 386276 560895
rect 386234 560552 386290 560561
rect 386234 560487 386290 560496
rect 386418 560552 386474 560561
rect 386418 560487 386474 560496
rect 386432 560402 386460 560487
rect 386510 560416 386566 560425
rect 386432 560374 386510 560402
rect 386510 560351 386566 560360
rect 385130 560008 385186 560017
rect 373184 559966 373566 559994
rect 375392 559966 375498 559994
rect 377048 559966 377430 559994
rect 378888 559966 379270 559994
rect 380912 559966 381202 559994
rect 386984 559980 387012 562294
rect 388916 559980 388944 562362
rect 390836 562284 390888 562290
rect 390836 562226 390888 562232
rect 390652 561060 390704 561066
rect 390652 561002 390704 561008
rect 389086 560144 389142 560153
rect 389086 560079 389142 560088
rect 385130 559943 385186 559952
rect 265808 559904 265860 559910
rect 263534 559842 263640 559858
rect 265466 559852 265808 559858
rect 372252 559904 372304 559910
rect 265466 559846 265860 559852
rect 291566 559872 291622 559881
rect 263534 559836 263652 559842
rect 263534 559830 263600 559836
rect 265466 559830 265848 559846
rect 291566 559807 291622 559816
rect 296626 559872 296682 559881
rect 296626 559807 296682 559816
rect 304262 559872 304318 559881
rect 372252 559846 372304 559852
rect 304262 559807 304318 559816
rect 263600 559778 263652 559784
rect 257738 559706 258120 559722
rect 257738 559700 258132 559706
rect 257738 559694 258080 559700
rect 258080 559642 258132 559648
rect 248788 559632 248840 559638
rect 246146 559570 246528 559586
rect 252192 559632 252244 559638
rect 248788 559574 248840 559580
rect 251942 559580 252192 559586
rect 251942 559574 252244 559580
rect 252650 559600 252706 559609
rect 246146 559564 246540 559570
rect 246146 559558 246488 559564
rect 246488 559506 246540 559512
rect 240140 559496 240192 559502
rect 240138 559464 240140 559473
rect 240600 559496 240652 559502
rect 240192 559464 240194 559473
rect 240350 559444 240600 559450
rect 240350 559438 240652 559444
rect 240350 559422 240640 559438
rect 240138 559399 240194 559408
rect 248800 559337 248828 559574
rect 251942 559558 252232 559574
rect 252650 559535 252706 559544
rect 277306 559600 277362 559609
rect 277306 559535 277362 559544
rect 231030 559328 231086 559337
rect 230782 559286 231030 559314
rect 232870 559328 232926 559337
rect 232622 559286 232870 559314
rect 231030 559263 231086 559272
rect 234618 559328 234674 559337
rect 234554 559286 234618 559314
rect 232870 559263 232926 559272
rect 236734 559328 236790 559337
rect 236486 559286 236734 559314
rect 234618 559263 234674 559272
rect 236734 559263 236790 559272
rect 238206 559328 238262 559337
rect 248786 559328 248842 559337
rect 238262 559286 238418 559314
rect 238206 559263 238262 559272
rect 248786 559263 248842 559272
rect 252558 559328 252614 559337
rect 252664 559314 252692 559535
rect 277320 559337 277348 559535
rect 291580 559337 291608 559807
rect 296640 559609 296668 559807
rect 296626 559600 296682 559609
rect 296626 559535 296682 559544
rect 304276 559473 304304 559807
rect 369858 559600 369914 559609
rect 369858 559535 369914 559544
rect 304262 559464 304318 559473
rect 304262 559399 304318 559408
rect 361316 559422 361528 559450
rect 361316 559337 361344 559422
rect 361500 559337 361528 559422
rect 369872 559366 369900 559535
rect 384868 559434 385066 559450
rect 384856 559428 385066 559434
rect 384908 559422 385066 559428
rect 384856 559370 384908 559376
rect 385144 559366 385172 559943
rect 389100 559910 389128 560079
rect 389088 559904 389140 559910
rect 389088 559846 389140 559852
rect 390560 559768 390612 559774
rect 390664 559722 390692 561002
rect 390848 559980 390876 562226
rect 392768 562216 392820 562222
rect 392768 562158 392820 562164
rect 392780 559980 392808 562158
rect 394700 562148 394752 562154
rect 394700 562090 394752 562096
rect 394712 559980 394740 562090
rect 396632 562080 396684 562086
rect 396632 562022 396684 562028
rect 395802 560416 395858 560425
rect 395986 560416 396042 560425
rect 395858 560374 395986 560402
rect 395802 560351 395858 560360
rect 395986 560351 396042 560360
rect 396644 559980 396672 562022
rect 398564 562012 398616 562018
rect 398564 561954 398616 561960
rect 398576 559980 398604 561954
rect 400496 561944 400548 561950
rect 400496 561886 400548 561892
rect 400218 560824 400274 560833
rect 400218 560759 400220 560768
rect 400272 560759 400274 560768
rect 400220 560730 400272 560736
rect 398930 560552 398986 560561
rect 398760 560510 398930 560538
rect 398760 560425 398788 560510
rect 398930 560487 398986 560496
rect 398746 560416 398802 560425
rect 398746 560351 398802 560360
rect 400218 560416 400274 560425
rect 400218 560351 400220 560360
rect 400272 560351 400274 560360
rect 400220 560322 400272 560328
rect 400218 560280 400274 560289
rect 400218 560215 400220 560224
rect 400272 560215 400274 560224
rect 400220 560186 400272 560192
rect 400218 560144 400274 560153
rect 400218 560079 400220 560088
rect 400272 560079 400274 560088
rect 400220 560050 400272 560056
rect 400218 560008 400274 560017
rect 400508 559980 400536 561886
rect 402428 561876 402480 561882
rect 402428 561818 402480 561824
rect 400586 560824 400642 560833
rect 400586 560759 400588 560768
rect 400640 560759 400642 560768
rect 400588 560730 400640 560736
rect 400586 560416 400642 560425
rect 400586 560351 400588 560360
rect 400640 560351 400642 560360
rect 400588 560322 400640 560328
rect 400586 560280 400642 560289
rect 400586 560215 400588 560224
rect 400640 560215 400642 560224
rect 400588 560186 400640 560192
rect 400586 560144 400642 560153
rect 400586 560079 400588 560088
rect 400640 560079 400642 560088
rect 400588 560050 400640 560056
rect 400586 560008 400642 560017
rect 400218 559943 400220 559952
rect 400272 559943 400274 559952
rect 402440 559980 402468 561818
rect 404372 559980 404400 562799
rect 408224 561808 408276 561814
rect 408224 561750 408276 561756
rect 405738 560552 405794 560561
rect 405738 560487 405794 560496
rect 405752 560402 405780 560487
rect 405830 560416 405886 560425
rect 405752 560374 405830 560402
rect 405830 560351 405886 560360
rect 408236 559980 408264 561750
rect 410156 560584 410208 560590
rect 410156 560526 410208 560532
rect 411352 560584 411404 560590
rect 411352 560526 411404 560532
rect 410168 559980 410196 560526
rect 411258 560416 411314 560425
rect 411258 560351 411314 560360
rect 411272 560266 411300 560351
rect 411364 560266 411392 560526
rect 411272 560238 411392 560266
rect 412100 559980 412128 562974
rect 450452 562964 450504 562970
rect 450452 562906 450504 562912
rect 450360 562896 450412 562902
rect 450360 562838 450412 562844
rect 415950 562728 416006 562737
rect 415950 562663 416006 562672
rect 441066 562728 441122 562737
rect 441066 562663 441122 562672
rect 414020 561740 414072 561746
rect 414020 561682 414072 561688
rect 414032 559980 414060 561682
rect 415964 559980 415992 562663
rect 419814 562320 419870 562329
rect 419814 562255 419870 562264
rect 417884 562148 417936 562154
rect 417884 562090 417936 562096
rect 417896 559980 417924 562090
rect 419828 559980 419856 562255
rect 423678 562184 423734 562193
rect 423678 562119 423734 562128
rect 421748 560516 421800 560522
rect 421748 560458 421800 560464
rect 421760 559980 421788 560458
rect 423692 559980 423720 562119
rect 425610 562048 425666 562057
rect 425610 561983 425666 561992
rect 424322 560824 424378 560833
rect 424322 560759 424378 560768
rect 424336 560590 424364 560759
rect 424324 560584 424376 560590
rect 424324 560526 424376 560532
rect 425624 559980 425652 561983
rect 429474 561912 429530 561921
rect 429474 561847 429530 561856
rect 427544 560448 427596 560454
rect 427544 560390 427596 560396
rect 427556 559980 427584 560390
rect 429488 559980 429516 561847
rect 437202 561776 437258 561785
rect 437202 561711 437258 561720
rect 431866 560824 431922 560833
rect 431866 560759 431922 560768
rect 431880 560561 431908 560759
rect 431866 560552 431922 560561
rect 431866 560487 431922 560496
rect 433340 560380 433392 560386
rect 433340 560322 433392 560328
rect 433352 559980 433380 560322
rect 437216 559980 437244 561711
rect 439136 560312 439188 560318
rect 439136 560254 439188 560260
rect 439148 559980 439176 560254
rect 441080 559980 441108 562663
rect 450268 560856 450320 560862
rect 450268 560798 450320 560804
rect 449624 560788 449676 560794
rect 449624 560730 449676 560736
rect 400586 559943 400588 559952
rect 400220 559914 400272 559920
rect 400640 559943 400642 559952
rect 400588 559914 400640 559920
rect 400312 559904 400364 559910
rect 400310 559872 400312 559881
rect 400680 559904 400732 559910
rect 400364 559872 400366 559881
rect 400310 559807 400366 559816
rect 400678 559872 400680 559881
rect 409880 559904 409932 559910
rect 400732 559872 400734 559881
rect 400678 559807 400734 559816
rect 409878 559872 409880 559881
rect 419356 559904 419408 559910
rect 409932 559872 409934 559881
rect 409878 559807 409934 559816
rect 419354 559872 419356 559881
rect 419408 559872 419410 559881
rect 419354 559807 419410 559816
rect 390612 559716 390692 559722
rect 390560 559710 390692 559716
rect 390572 559694 390692 559710
rect 394054 559600 394110 559609
rect 394054 559535 394110 559544
rect 405922 559600 405978 559609
rect 405978 559558 406318 559586
rect 405922 559535 405978 559544
rect 369860 559360 369912 559366
rect 252614 559286 252692 559314
rect 277306 559328 277362 559337
rect 252558 559263 252614 559272
rect 277306 559263 277362 559272
rect 291566 559328 291622 559337
rect 291566 559263 291622 559272
rect 361302 559328 361358 559337
rect 361302 559263 361358 559272
rect 361486 559328 361542 559337
rect 385132 559360 385184 559366
rect 383198 559328 383254 559337
rect 369860 559302 369912 559308
rect 383134 559286 383198 559314
rect 361486 559263 361542 559272
rect 394068 559337 394096 559535
rect 434626 559464 434682 559473
rect 396092 559434 396396 559450
rect 396092 559428 396408 559434
rect 396092 559422 396356 559428
rect 396092 559366 396120 559422
rect 442814 559464 442870 559473
rect 435008 559434 435298 559450
rect 434626 559399 434682 559408
rect 434996 559428 435298 559434
rect 396356 559370 396408 559376
rect 396080 559360 396132 559366
rect 385132 559302 385184 559308
rect 394054 559328 394110 559337
rect 383198 559263 383254 559272
rect 396080 559302 396132 559308
rect 431132 559360 431184 559366
rect 434640 559337 434668 559399
rect 435048 559422 435298 559428
rect 442870 559422 443026 559450
rect 442814 559399 442870 559408
rect 434996 559370 435048 559376
rect 434626 559328 434682 559337
rect 431184 559308 431434 559314
rect 431132 559302 431434 559308
rect 431144 559286 431434 559302
rect 394054 559263 394110 559272
rect 434626 559263 434682 559272
rect 444562 559328 444618 559337
rect 446586 559328 446642 559337
rect 444618 559286 444958 559314
rect 444562 559263 444618 559272
rect 448518 559328 448574 559337
rect 446642 559286 446890 559314
rect 446586 559263 446642 559272
rect 448574 559286 448822 559314
rect 448518 559263 448574 559272
rect 6644 495576 6696 495582
rect 6644 495518 6696 495524
rect 6552 481160 6604 481166
rect 6552 481102 6604 481108
rect 6460 438728 6512 438734
rect 6460 438670 6512 438676
rect 449636 394618 449664 560730
rect 450280 557326 450308 560798
rect 450268 557320 450320 557326
rect 450268 557262 450320 557268
rect 450372 557190 450400 562838
rect 450360 557184 450412 557190
rect 450360 557126 450412 557132
rect 450464 546446 450492 562906
rect 451096 562828 451148 562834
rect 451096 562770 451148 562776
rect 450728 562760 450780 562766
rect 450728 562702 450780 562708
rect 450636 562556 450688 562562
rect 450636 562498 450688 562504
rect 450544 560720 450596 560726
rect 450544 560662 450596 560668
rect 450452 546440 450504 546446
rect 450452 546382 450504 546388
rect 449636 394590 449756 394618
rect 449728 393310 449756 394590
rect 449716 393304 449768 393310
rect 449716 393246 449768 393252
rect 6368 380656 6420 380662
rect 6368 380598 6420 380604
rect 450556 346390 450584 560662
rect 450648 369850 450676 562498
rect 450740 405686 450768 562702
rect 451004 562692 451056 562698
rect 451004 562634 451056 562640
rect 450820 560992 450872 560998
rect 450820 560934 450872 560940
rect 450832 557530 450860 560934
rect 450820 557524 450872 557530
rect 450820 557466 450872 557472
rect 451016 557410 451044 562634
rect 450832 557382 451044 557410
rect 450832 416770 450860 557382
rect 450912 557320 450964 557326
rect 451108 557274 451136 562770
rect 462964 562624 463016 562630
rect 462964 562566 463016 562572
rect 580538 562592 580594 562601
rect 451188 560924 451240 560930
rect 451188 560866 451240 560872
rect 450912 557262 450964 557268
rect 450924 440230 450952 557262
rect 451016 557246 451136 557274
rect 451016 463690 451044 557246
rect 451096 557184 451148 557190
rect 451096 557126 451148 557132
rect 451108 499526 451136 557126
rect 451200 510610 451228 560866
rect 451188 510604 451240 510610
rect 451188 510546 451240 510552
rect 451096 499520 451148 499526
rect 451096 499462 451148 499468
rect 451004 463684 451056 463690
rect 451004 463626 451056 463632
rect 462976 452606 463004 562566
rect 580538 562527 580594 562536
rect 580354 562456 580410 562465
rect 580354 562391 580410 562400
rect 548524 560652 548576 560658
rect 548524 560594 548576 560600
rect 548536 534070 548564 560594
rect 579804 560244 579856 560250
rect 579804 560186 579856 560192
rect 577596 559972 577648 559978
rect 577596 559914 577648 559920
rect 577504 559904 577556 559910
rect 577504 559846 577556 559852
rect 548524 534064 548576 534070
rect 548524 534006 548576 534012
rect 462964 452600 463016 452606
rect 462964 452542 463016 452548
rect 450912 440224 450964 440230
rect 450912 440166 450964 440172
rect 450820 416764 450872 416770
rect 450820 416706 450872 416712
rect 450728 405680 450780 405686
rect 450728 405622 450780 405628
rect 450636 369844 450688 369850
rect 450636 369786 450688 369792
rect 450544 346384 450596 346390
rect 450544 346326 450596 346332
rect 327460 340190 327842 340218
rect 337396 340190 337778 340218
rect 363892 340190 364182 340218
rect 384422 340190 384804 340218
rect 388470 340190 388852 340218
rect 420302 340190 420684 340218
rect 447718 340190 448100 340218
rect 229112 340054 230046 340082
rect 230124 340054 230414 340082
rect 230492 340054 230874 340082
rect 231044 340054 231334 340082
rect 79324 338088 79376 338094
rect 79324 338030 79376 338036
rect 71044 338020 71096 338026
rect 71044 337962 71096 337968
rect 66904 337952 66956 337958
rect 66904 337894 66956 337900
rect 61384 337884 61436 337890
rect 61384 337826 61436 337832
rect 57244 337816 57296 337822
rect 57244 337758 57296 337764
rect 42064 337748 42116 337754
rect 42064 337690 42116 337696
rect 39304 337680 39356 337686
rect 39304 337622 39356 337628
rect 35164 337612 35216 337618
rect 35164 337554 35216 337560
rect 28264 337544 28316 337550
rect 28264 337486 28316 337492
rect 19984 337476 20036 337482
rect 19984 337418 20036 337424
rect 13084 337408 13136 337414
rect 10322 337376 10378 337385
rect 13084 337350 13136 337356
rect 10322 337311 10378 337320
rect 6276 280152 6328 280158
rect 6276 280094 6328 280100
rect 6184 79484 6236 79490
rect 6184 79426 6236 79432
rect 4122 50102 4200 50130
rect 4066 50079 4122 50088
rect 4066 8256 4122 8265
rect 4066 8191 4122 8200
rect 3974 7576 4030 7585
rect 3974 7511 4030 7520
rect 2872 4956 2924 4962
rect 2872 4898 2924 4904
rect 572 4820 624 4826
rect 572 4762 624 4768
rect 584 480 612 4762
rect 1676 4752 1728 4758
rect 1676 4694 1728 4700
rect 1688 480 1716 4694
rect 2884 480 2912 4898
rect 3988 626 4016 7511
rect 4080 7177 4108 8191
rect 8852 7608 8904 7614
rect 8852 7550 8904 7556
rect 4066 7168 4122 7177
rect 4066 7103 4122 7112
rect 7656 5024 7708 5030
rect 7656 4966 7708 4972
rect 5264 4140 5316 4146
rect 5264 4082 5316 4088
rect 3988 598 4108 626
rect 4080 480 4108 598
rect 5276 480 5304 4082
rect 6458 3360 6514 3369
rect 6458 3295 6514 3304
rect 6472 480 6500 3295
rect 7668 480 7696 4966
rect 8864 480 8892 7550
rect 10336 4146 10364 337311
rect 12440 5092 12492 5098
rect 12440 5034 12492 5040
rect 10324 4140 10376 4146
rect 10324 4082 10376 4088
rect 11244 3596 11296 3602
rect 11244 3538 11296 3544
rect 10048 3324 10100 3330
rect 10048 3266 10100 3272
rect 10060 480 10088 3266
rect 11256 480 11284 3538
rect 12452 480 12480 5034
rect 13096 3330 13124 337350
rect 18328 11756 18380 11762
rect 18328 11698 18380 11704
rect 13636 8968 13688 8974
rect 13636 8910 13688 8916
rect 13084 3324 13136 3330
rect 13084 3266 13136 3272
rect 13648 480 13676 8910
rect 17224 7676 17276 7682
rect 17224 7618 17276 7624
rect 16028 3528 16080 3534
rect 16028 3470 16080 3476
rect 14832 3460 14884 3466
rect 14832 3402 14884 3408
rect 14844 480 14872 3402
rect 16040 480 16068 3470
rect 17236 480 17264 7618
rect 18340 480 18368 11698
rect 19996 3602 20024 337418
rect 23388 13116 23440 13122
rect 23388 13058 23440 13064
rect 21916 7744 21968 7750
rect 21916 7686 21968 7692
rect 20720 3936 20772 3942
rect 20720 3878 20772 3884
rect 19984 3596 20036 3602
rect 19984 3538 20036 3544
rect 19524 3392 19576 3398
rect 19524 3334 19576 3340
rect 19536 480 19564 3334
rect 20732 480 20760 3878
rect 21928 480 21956 7686
rect 23400 610 23428 13058
rect 27896 9036 27948 9042
rect 27896 8978 27948 8984
rect 26700 7812 26752 7818
rect 26700 7754 26752 7760
rect 25504 3664 25556 3670
rect 25504 3606 25556 3612
rect 24308 3596 24360 3602
rect 24308 3538 24360 3544
rect 23112 604 23164 610
rect 23112 546 23164 552
rect 23388 604 23440 610
rect 23388 546 23440 552
rect 23124 480 23152 546
rect 24320 480 24348 3538
rect 25516 480 25544 3606
rect 26712 480 26740 7754
rect 27908 480 27936 8978
rect 28276 3398 28304 337486
rect 31668 14476 31720 14482
rect 31668 14418 31720 14424
rect 30288 7880 30340 7886
rect 30288 7822 30340 7828
rect 28264 3392 28316 3398
rect 28264 3334 28316 3340
rect 29092 3324 29144 3330
rect 29092 3266 29144 3272
rect 29104 480 29132 3266
rect 30300 480 30328 7822
rect 31680 626 31708 14418
rect 33876 7948 33928 7954
rect 33876 7890 33928 7896
rect 32680 3732 32732 3738
rect 32680 3674 32732 3680
rect 31496 598 31708 626
rect 31496 480 31524 598
rect 32692 480 32720 3674
rect 33888 480 33916 7890
rect 34980 3392 35032 3398
rect 34980 3334 35032 3340
rect 34992 480 35020 3334
rect 35176 3330 35204 337554
rect 37372 8016 37424 8022
rect 37372 7958 37424 7964
rect 36176 4140 36228 4146
rect 36176 4082 36228 4088
rect 35164 3324 35216 3330
rect 35164 3266 35216 3272
rect 36188 480 36216 4082
rect 37384 480 37412 7958
rect 39316 4146 39344 337622
rect 40960 9104 41012 9110
rect 40960 9046 41012 9052
rect 39304 4140 39356 4146
rect 39304 4082 39356 4088
rect 39764 3868 39816 3874
rect 39764 3810 39816 3816
rect 38568 3800 38620 3806
rect 38568 3742 38620 3748
rect 38580 480 38608 3742
rect 39776 480 39804 3810
rect 40972 480 41000 9046
rect 42076 3942 42104 337690
rect 56416 10464 56468 10470
rect 56416 10406 56468 10412
rect 52828 10396 52880 10402
rect 52828 10338 52880 10344
rect 49332 10328 49384 10334
rect 49332 10270 49384 10276
rect 44548 9172 44600 9178
rect 44548 9114 44600 9120
rect 42064 3936 42116 3942
rect 42064 3878 42116 3884
rect 42156 3324 42208 3330
rect 42156 3266 42208 3272
rect 42168 480 42196 3266
rect 43352 3256 43404 3262
rect 43352 3198 43404 3204
rect 43364 480 43392 3198
rect 44560 480 44588 9114
rect 48136 5160 48188 5166
rect 48136 5102 48188 5108
rect 46940 4004 46992 4010
rect 46940 3946 46992 3952
rect 45744 3936 45796 3942
rect 45744 3878 45796 3884
rect 45756 480 45784 3878
rect 46952 480 46980 3946
rect 48148 480 48176 5102
rect 49344 480 49372 10270
rect 51632 5228 51684 5234
rect 51632 5170 51684 5176
rect 50528 4072 50580 4078
rect 50528 4014 50580 4020
rect 50540 480 50568 4014
rect 51644 480 51672 5170
rect 52840 480 52868 10338
rect 55218 6216 55274 6225
rect 55218 6151 55274 6160
rect 54024 3188 54076 3194
rect 54024 3130 54076 3136
rect 54036 480 54064 3130
rect 55232 480 55260 6151
rect 56428 480 56456 10406
rect 57256 3398 57284 337758
rect 60004 10532 60056 10538
rect 60004 10474 60056 10480
rect 58808 6180 58860 6186
rect 58808 6122 58860 6128
rect 57612 4140 57664 4146
rect 57612 4082 57664 4088
rect 57244 3392 57296 3398
rect 57244 3334 57296 3340
rect 57624 480 57652 4082
rect 58820 480 58848 6122
rect 60016 480 60044 10474
rect 61396 3262 61424 337826
rect 63592 10600 63644 10606
rect 63592 10542 63644 10548
rect 62396 6248 62448 6254
rect 62396 6190 62448 6196
rect 61384 3256 61436 3262
rect 61384 3198 61436 3204
rect 61200 3120 61252 3126
rect 61200 3062 61252 3068
rect 61212 480 61240 3062
rect 62408 480 62436 6190
rect 63604 480 63632 10542
rect 65984 6316 66036 6322
rect 65984 6258 66036 6264
rect 64696 3392 64748 3398
rect 64696 3334 64748 3340
rect 64708 1714 64736 3334
rect 64708 1686 64828 1714
rect 64800 480 64828 1686
rect 65996 480 66024 6258
rect 66916 3330 66944 337894
rect 69480 6384 69532 6390
rect 69480 6326 69532 6332
rect 67180 5296 67232 5302
rect 67180 5238 67232 5244
rect 66904 3324 66956 3330
rect 66904 3266 66956 3272
rect 67192 480 67220 5238
rect 68284 3052 68336 3058
rect 68284 2994 68336 3000
rect 68296 480 68324 2994
rect 69492 480 69520 6326
rect 70676 3324 70728 3330
rect 70676 3266 70728 3272
rect 70688 480 70716 3266
rect 71056 3194 71084 337962
rect 77944 337272 77996 337278
rect 77944 337214 77996 337220
rect 74448 14544 74500 14550
rect 74448 14486 74500 14492
rect 71688 13184 71740 13190
rect 71688 13126 71740 13132
rect 71700 3330 71728 13126
rect 73068 6452 73120 6458
rect 73068 6394 73120 6400
rect 71688 3324 71740 3330
rect 71688 3266 71740 3272
rect 71872 3324 71924 3330
rect 71872 3266 71924 3272
rect 71044 3188 71096 3194
rect 71044 3130 71096 3136
rect 71884 480 71912 3266
rect 73080 480 73108 6394
rect 74460 3380 74488 14486
rect 76656 6520 76708 6526
rect 76656 6462 76708 6468
rect 74276 3352 74488 3380
rect 74276 480 74304 3352
rect 75460 3188 75512 3194
rect 75460 3130 75512 3136
rect 75472 480 75500 3130
rect 76668 480 76696 6462
rect 77852 3256 77904 3262
rect 77852 3198 77904 3204
rect 77864 480 77892 3198
rect 77956 3126 77984 337214
rect 78588 14612 78640 14618
rect 78588 14554 78640 14560
rect 78600 3262 78628 14554
rect 78588 3256 78640 3262
rect 78588 3198 78640 3204
rect 79336 3194 79364 338030
rect 138020 337340 138072 337346
rect 138020 337282 138072 337288
rect 147588 337340 147640 337346
rect 147588 337282 147640 337288
rect 157340 337340 157392 337346
rect 157340 337282 157392 337288
rect 166908 337340 166960 337346
rect 166908 337282 166960 337288
rect 176660 337340 176712 337346
rect 176660 337282 176712 337288
rect 186228 337340 186280 337346
rect 186228 337282 186280 337288
rect 195980 337340 196032 337346
rect 195980 337282 196032 337288
rect 205548 337340 205600 337346
rect 205548 337282 205600 337288
rect 215300 337340 215352 337346
rect 215300 337282 215352 337288
rect 224868 337340 224920 337346
rect 224868 337282 224920 337288
rect 138032 337249 138060 337282
rect 147600 337249 147628 337282
rect 157352 337249 157380 337282
rect 166920 337249 166948 337282
rect 176672 337249 176700 337282
rect 186240 337249 186268 337282
rect 195992 337249 196020 337282
rect 205560 337249 205588 337282
rect 215312 337249 215340 337282
rect 224880 337249 224908 337282
rect 138018 337240 138074 337249
rect 97264 337204 97316 337210
rect 138018 337175 138074 337184
rect 147586 337240 147642 337249
rect 147586 337175 147642 337184
rect 157338 337240 157394 337249
rect 157338 337175 157394 337184
rect 166906 337240 166962 337249
rect 166906 337175 166962 337184
rect 176658 337240 176714 337249
rect 176658 337175 176714 337184
rect 186226 337240 186282 337249
rect 186226 337175 186282 337184
rect 195978 337240 196034 337249
rect 195978 337175 196034 337184
rect 205546 337240 205602 337249
rect 205546 337175 205602 337184
rect 215298 337240 215354 337249
rect 215298 337175 215354 337184
rect 224866 337240 224922 337249
rect 224866 337175 224922 337184
rect 97264 337146 97316 337152
rect 84844 337136 84896 337142
rect 84844 337078 84896 337084
rect 82728 14680 82780 14686
rect 82728 14622 82780 14628
rect 80244 8084 80296 8090
rect 80244 8026 80296 8032
rect 79324 3188 79376 3194
rect 79324 3130 79376 3136
rect 77944 3120 77996 3126
rect 77944 3062 77996 3068
rect 79048 2984 79100 2990
rect 79048 2926 79100 2932
rect 79060 480 79088 2926
rect 80256 480 80284 8026
rect 82740 3262 82768 14622
rect 83832 8152 83884 8158
rect 83832 8094 83884 8100
rect 81440 3256 81492 3262
rect 81440 3198 81492 3204
rect 82728 3256 82780 3262
rect 82728 3198 82780 3204
rect 81452 480 81480 3198
rect 82636 3188 82688 3194
rect 82636 3130 82688 3136
rect 82648 480 82676 3130
rect 83844 480 83872 8094
rect 84856 3262 84884 337078
rect 96528 14952 96580 14958
rect 96528 14894 96580 14900
rect 92388 14884 92440 14890
rect 92388 14826 92440 14832
rect 89628 14816 89680 14822
rect 89628 14758 89680 14764
rect 85488 14748 85540 14754
rect 85488 14690 85540 14696
rect 85500 3262 85528 14690
rect 87328 8220 87380 8226
rect 87328 8162 87380 8168
rect 84844 3256 84896 3262
rect 84844 3198 84896 3204
rect 84936 3256 84988 3262
rect 84936 3198 84988 3204
rect 85488 3256 85540 3262
rect 85488 3198 85540 3204
rect 84948 480 84976 3198
rect 86132 2984 86184 2990
rect 86132 2926 86184 2932
rect 86144 480 86172 2926
rect 87340 480 87368 8162
rect 89640 3262 89668 14758
rect 91008 10668 91060 10674
rect 91008 10610 91060 10616
rect 91020 3482 91048 10610
rect 92400 3482 92428 14826
rect 95148 10736 95200 10742
rect 95148 10678 95200 10684
rect 90928 3454 91048 3482
rect 92124 3454 92428 3482
rect 88524 3256 88576 3262
rect 88524 3198 88576 3204
rect 89628 3256 89680 3262
rect 89628 3198 89680 3204
rect 88536 480 88564 3198
rect 89720 3120 89772 3126
rect 89720 3062 89772 3068
rect 89732 480 89760 3062
rect 90928 480 90956 3454
rect 92124 480 92152 3454
rect 95160 3126 95188 10678
rect 96540 3126 96568 14894
rect 94504 3120 94556 3126
rect 94504 3062 94556 3068
rect 95148 3120 95200 3126
rect 95148 3062 95200 3068
rect 95700 3120 95752 3126
rect 95700 3062 95752 3068
rect 96528 3120 96580 3126
rect 96528 3062 96580 3068
rect 93308 2916 93360 2922
rect 93308 2858 93360 2864
rect 93320 480 93348 2858
rect 94516 480 94544 3062
rect 95712 480 95740 3062
rect 97276 2922 97304 337146
rect 100668 337136 100720 337142
rect 100668 337078 100720 337084
rect 99288 15020 99340 15026
rect 99288 14962 99340 14968
rect 99196 10804 99248 10810
rect 99196 10746 99248 10752
rect 99208 3126 99236 10746
rect 98092 3120 98144 3126
rect 98092 3062 98144 3068
rect 99196 3120 99248 3126
rect 99196 3062 99248 3068
rect 97264 2916 97316 2922
rect 97264 2858 97316 2864
rect 96896 2848 96948 2854
rect 96896 2790 96948 2796
rect 96908 480 96936 2790
rect 98104 480 98132 3062
rect 99300 480 99328 14962
rect 100680 3346 100708 337078
rect 107568 337068 107620 337074
rect 107568 337010 107620 337016
rect 105544 337000 105596 337006
rect 105544 336942 105596 336948
rect 102784 336864 102836 336870
rect 102784 336806 102836 336812
rect 102048 10872 102100 10878
rect 102048 10814 102100 10820
rect 100496 3318 100708 3346
rect 100496 480 100524 3318
rect 102060 3126 102088 10814
rect 102796 3210 102824 336806
rect 103428 15088 103480 15094
rect 103428 15030 103480 15036
rect 102612 3182 102824 3210
rect 101588 3120 101640 3126
rect 101588 3062 101640 3068
rect 102048 3120 102100 3126
rect 102048 3062 102100 3068
rect 101600 480 101628 3062
rect 102612 3058 102640 3182
rect 103440 3126 103468 15030
rect 102784 3120 102836 3126
rect 102784 3062 102836 3068
rect 103428 3120 103480 3126
rect 103428 3062 103480 3068
rect 105176 3120 105228 3126
rect 105176 3062 105228 3068
rect 102600 3052 102652 3058
rect 102600 2994 102652 3000
rect 102796 480 102824 3062
rect 103980 2916 104032 2922
rect 103980 2858 104032 2864
rect 103992 480 104020 2858
rect 105188 480 105216 3062
rect 105556 2854 105584 336942
rect 107476 15156 107528 15162
rect 107476 15098 107528 15104
rect 106188 10940 106240 10946
rect 106188 10882 106240 10888
rect 106200 3126 106228 10882
rect 107488 3126 107516 15098
rect 106188 3120 106240 3126
rect 106188 3062 106240 3068
rect 106372 3120 106424 3126
rect 106372 3062 106424 3068
rect 107476 3120 107528 3126
rect 107476 3062 107528 3068
rect 105544 2848 105596 2854
rect 105544 2790 105596 2796
rect 106384 480 106412 3062
rect 107580 480 107608 337010
rect 118608 336932 118660 336938
rect 118608 336874 118660 336880
rect 110328 14408 110380 14414
rect 110328 14350 110380 14356
rect 108948 11008 109000 11014
rect 108948 10950 109000 10956
rect 108960 3346 108988 10950
rect 110340 3346 110368 14350
rect 114468 14340 114520 14346
rect 114468 14282 114520 14288
rect 113088 10260 113140 10266
rect 113088 10202 113140 10208
rect 108776 3318 108988 3346
rect 109972 3318 110368 3346
rect 108776 480 108804 3318
rect 109972 480 110000 3318
rect 113100 2990 113128 10202
rect 114480 2990 114508 14282
rect 117228 14272 117280 14278
rect 117228 14214 117280 14220
rect 117136 10192 117188 10198
rect 117136 10134 117188 10140
rect 117148 3618 117176 10134
rect 116964 3590 117176 3618
rect 116964 2990 116992 3590
rect 117240 3482 117268 14214
rect 117148 3454 117268 3482
rect 112352 2984 112404 2990
rect 112352 2926 112404 2932
rect 113088 2984 113140 2990
rect 113088 2926 113140 2932
rect 113548 2984 113600 2990
rect 113548 2926 113600 2932
rect 114468 2984 114520 2990
rect 114468 2926 114520 2932
rect 115940 2984 115992 2990
rect 115940 2926 115992 2932
rect 116952 2984 117004 2990
rect 116952 2926 117004 2932
rect 111156 2916 111208 2922
rect 111156 2858 111208 2864
rect 111168 480 111196 2858
rect 112364 480 112392 2926
rect 113560 480 113588 2926
rect 114744 2848 114796 2854
rect 114744 2790 114796 2796
rect 114756 480 114784 2790
rect 115952 480 115980 2926
rect 117148 480 117176 3454
rect 118620 3346 118648 336874
rect 125508 336796 125560 336802
rect 125508 336738 125560 336744
rect 121368 14204 121420 14210
rect 121368 14146 121420 14152
rect 119988 10124 120040 10130
rect 119988 10066 120040 10072
rect 118252 3318 118648 3346
rect 118252 480 118280 3318
rect 120000 2990 120028 10066
rect 121380 2990 121408 14146
rect 125416 14136 125468 14142
rect 125416 14078 125468 14084
rect 124128 10056 124180 10062
rect 124128 9998 124180 10004
rect 124140 3482 124168 9998
rect 125428 4214 125456 14078
rect 124220 4208 124272 4214
rect 124220 4150 124272 4156
rect 125416 4208 125468 4214
rect 125416 4150 125468 4156
rect 123036 3454 124168 3482
rect 119436 2984 119488 2990
rect 119436 2926 119488 2932
rect 119988 2984 120040 2990
rect 119988 2926 120040 2932
rect 120632 2984 120684 2990
rect 120632 2926 120684 2932
rect 121368 2984 121420 2990
rect 121368 2926 121420 2932
rect 119448 480 119476 2926
rect 120644 480 120672 2926
rect 121828 2848 121880 2854
rect 121828 2790 121880 2796
rect 121840 480 121868 2790
rect 123036 480 123064 3454
rect 124232 480 124260 4150
rect 125520 3482 125548 336738
rect 197268 14068 197320 14074
rect 197268 14010 197320 14016
rect 190368 13796 190420 13802
rect 190368 13738 190420 13744
rect 186228 13728 186280 13734
rect 186228 13670 186280 13676
rect 183468 13660 183520 13666
rect 183468 13602 183520 13608
rect 179328 13592 179380 13598
rect 179328 13534 179380 13540
rect 176568 13524 176620 13530
rect 176568 13466 176620 13472
rect 172428 13456 172480 13462
rect 172428 13398 172480 13404
rect 160008 13388 160060 13394
rect 160008 13330 160060 13336
rect 155868 13320 155920 13326
rect 155868 13262 155920 13268
rect 135168 13252 135220 13258
rect 135168 13194 135220 13200
rect 128268 11892 128320 11898
rect 128268 11834 128320 11840
rect 126888 11824 126940 11830
rect 126888 11766 126940 11772
rect 126900 3482 126928 11766
rect 128280 3482 128308 11834
rect 132590 8936 132646 8945
rect 132590 8871 132646 8880
rect 129004 8288 129056 8294
rect 129004 8230 129056 8236
rect 125428 3454 125548 3482
rect 126624 3454 126928 3482
rect 127820 3454 128308 3482
rect 125428 480 125456 3454
rect 126624 480 126652 3454
rect 127820 480 127848 3454
rect 129016 480 129044 8230
rect 131396 6588 131448 6594
rect 131396 6530 131448 6536
rect 130200 5364 130252 5370
rect 130200 5306 130252 5312
rect 130212 480 130240 5306
rect 131408 480 131436 6530
rect 132604 480 132632 8871
rect 133788 5432 133840 5438
rect 133788 5374 133840 5380
rect 133800 480 133828 5374
rect 135180 626 135208 13194
rect 151728 12164 151780 12170
rect 151728 12106 151780 12112
rect 148968 12096 149020 12102
rect 148968 12038 149020 12044
rect 144828 12028 144880 12034
rect 144828 11970 144880 11976
rect 140872 11960 140924 11966
rect 140872 11902 140924 11908
rect 139676 9308 139728 9314
rect 139676 9250 139728 9256
rect 136088 9240 136140 9246
rect 136088 9182 136140 9188
rect 134904 598 135208 626
rect 134904 480 134932 598
rect 136100 480 136128 9182
rect 138480 7540 138532 7546
rect 138480 7482 138532 7488
rect 137284 5500 137336 5506
rect 137284 5442 137336 5448
rect 137296 480 137324 5442
rect 138492 480 138520 7482
rect 139688 480 139716 9250
rect 140884 480 140912 11902
rect 143264 9376 143316 9382
rect 143264 9318 143316 9324
rect 142068 7472 142120 7478
rect 142068 7414 142120 7420
rect 142080 480 142108 7414
rect 143276 480 143304 9318
rect 144840 626 144868 11970
rect 146852 9444 146904 9450
rect 146852 9386 146904 9392
rect 145656 7404 145708 7410
rect 145656 7346 145708 7352
rect 144472 598 144868 626
rect 144472 480 144500 598
rect 145668 480 145696 7346
rect 146864 480 146892 9386
rect 148980 610 149008 12038
rect 150440 9512 150492 9518
rect 150440 9454 150492 9460
rect 149244 7336 149296 7342
rect 149244 7278 149296 7284
rect 148048 604 148100 610
rect 148048 546 148100 552
rect 148968 604 149020 610
rect 148968 546 149020 552
rect 148060 480 148088 546
rect 149256 480 149284 7278
rect 150452 480 150480 9454
rect 151740 610 151768 12106
rect 154488 9988 154540 9994
rect 154488 9930 154540 9936
rect 152740 7268 152792 7274
rect 152740 7210 152792 7216
rect 151544 604 151596 610
rect 151544 546 151596 552
rect 151728 604 151780 610
rect 151728 546 151780 552
rect 151556 480 151584 546
rect 152752 480 152780 7210
rect 154500 610 154528 9930
rect 155880 610 155908 13262
rect 158628 9920 158680 9926
rect 158628 9862 158680 9868
rect 156328 7200 156380 7206
rect 156328 7142 156380 7148
rect 153936 604 153988 610
rect 153936 546 153988 552
rect 154488 604 154540 610
rect 154488 546 154540 552
rect 155132 604 155184 610
rect 155132 546 155184 552
rect 155868 604 155920 610
rect 155868 546 155920 552
rect 153948 480 153976 546
rect 155144 480 155172 546
rect 156340 480 156368 7142
rect 158640 610 158668 9862
rect 160020 7138 160048 13330
rect 169392 12368 169444 12374
rect 169392 12310 169444 12316
rect 165896 12300 165948 12306
rect 165896 12242 165948 12248
rect 162308 12232 162360 12238
rect 162308 12174 162360 12180
rect 161388 9852 161440 9858
rect 161388 9794 161440 9800
rect 158720 7132 158772 7138
rect 158720 7074 158772 7080
rect 160008 7132 160060 7138
rect 160008 7074 160060 7080
rect 157524 604 157576 610
rect 157524 546 157576 552
rect 158628 604 158680 610
rect 158628 546 158680 552
rect 157536 480 157564 546
rect 158732 480 158760 7074
rect 159916 7064 159968 7070
rect 159916 7006 159968 7012
rect 159928 480 159956 7006
rect 161400 610 161428 9794
rect 161112 604 161164 610
rect 161112 546 161164 552
rect 161388 604 161440 610
rect 161388 546 161440 552
rect 161124 480 161152 546
rect 162320 480 162348 12174
rect 164700 7064 164752 7070
rect 164700 7006 164752 7012
rect 163504 6656 163556 6662
rect 163504 6598 163556 6604
rect 163516 480 163544 6598
rect 164712 480 164740 7006
rect 165908 480 165936 12242
rect 168196 6996 168248 7002
rect 168196 6938 168248 6944
rect 167092 6724 167144 6730
rect 167092 6666 167144 6672
rect 167104 480 167132 6666
rect 168208 480 168236 6938
rect 169404 480 169432 12310
rect 170588 6792 170640 6798
rect 170588 6734 170640 6740
rect 170600 480 170628 6734
rect 172440 610 172468 13398
rect 173808 12436 173860 12442
rect 173808 12378 173860 12384
rect 173820 610 173848 12378
rect 176384 11688 176436 11694
rect 176384 11630 176436 11636
rect 175372 6928 175424 6934
rect 175372 6870 175424 6876
rect 174176 6860 174228 6866
rect 174176 6802 174228 6808
rect 171784 604 171836 610
rect 171784 546 171836 552
rect 172428 604 172480 610
rect 172428 546 172480 552
rect 172980 604 173032 610
rect 172980 546 173032 552
rect 173808 604 173860 610
rect 173808 546 173860 552
rect 171796 480 171824 546
rect 172992 480 173020 546
rect 174188 480 174216 6802
rect 175384 480 175412 6870
rect 176396 2802 176424 11630
rect 176580 6934 176608 13466
rect 176568 6928 176620 6934
rect 176568 6870 176620 6876
rect 177764 6112 177816 6118
rect 177764 6054 177816 6060
rect 176396 2774 176608 2802
rect 176580 480 176608 2774
rect 177776 480 177804 6054
rect 179340 610 179368 13534
rect 180708 11620 180760 11626
rect 180708 11562 180760 11568
rect 180720 610 180748 11562
rect 181352 6044 181404 6050
rect 181352 5986 181404 5992
rect 178960 604 179012 610
rect 178960 546 179012 552
rect 179328 604 179380 610
rect 179328 546 179380 552
rect 180156 604 180208 610
rect 180156 546 180208 552
rect 180708 604 180760 610
rect 180708 546 180760 552
rect 178972 480 179000 546
rect 180168 480 180196 546
rect 181364 480 181392 5986
rect 183480 610 183508 13602
rect 184756 11552 184808 11558
rect 184756 11494 184808 11500
rect 184768 610 184796 11494
rect 184848 5976 184900 5982
rect 184848 5918 184900 5924
rect 182548 604 182600 610
rect 182548 546 182600 552
rect 183468 604 183520 610
rect 183468 546 183520 552
rect 183744 604 183796 610
rect 183744 546 183796 552
rect 184756 604 184808 610
rect 184756 546 184808 552
rect 182560 480 182588 546
rect 183756 480 183784 546
rect 184860 480 184888 5918
rect 186240 626 186268 13670
rect 187608 11484 187660 11490
rect 187608 11426 187660 11432
rect 187620 626 187648 11426
rect 188436 5908 188488 5914
rect 188436 5850 188488 5856
rect 186148 598 186268 626
rect 187344 598 187648 626
rect 186148 592 186176 598
rect 187344 592 187372 598
rect 186056 564 186176 592
rect 187252 564 187372 592
rect 186056 480 186084 564
rect 187252 480 187280 564
rect 188448 480 188476 5850
rect 190380 610 190408 13738
rect 194508 13048 194560 13054
rect 194508 12990 194560 12996
rect 191748 11416 191800 11422
rect 191748 11358 191800 11364
rect 191760 610 191788 11358
rect 194416 11348 194468 11354
rect 194416 11290 194468 11296
rect 193220 6928 193272 6934
rect 193220 6870 193272 6876
rect 192024 5840 192076 5846
rect 192024 5782 192076 5788
rect 189632 604 189684 610
rect 189632 546 189684 552
rect 190368 604 190420 610
rect 190368 546 190420 552
rect 190828 604 190880 610
rect 190828 546 190880 552
rect 191748 604 191800 610
rect 191748 546 191800 552
rect 189644 480 189672 546
rect 190840 480 190868 546
rect 192036 480 192064 5782
rect 193232 480 193260 6870
rect 194428 480 194456 11290
rect 194520 6934 194548 12990
rect 194508 6928 194560 6934
rect 194508 6870 194560 6876
rect 195612 5772 195664 5778
rect 195612 5714 195664 5720
rect 195624 480 195652 5714
rect 197280 610 197308 14010
rect 211068 12980 211120 12986
rect 211068 12922 211120 12928
rect 198648 11280 198700 11286
rect 198648 11222 198700 11228
rect 198660 610 198688 11222
rect 203892 9648 203944 9654
rect 203892 9590 203944 9596
rect 200396 9580 200448 9586
rect 200396 9522 200448 9528
rect 199200 5704 199252 5710
rect 199200 5646 199252 5652
rect 196808 604 196860 610
rect 196808 546 196860 552
rect 197268 604 197320 610
rect 197268 546 197320 552
rect 198004 604 198056 610
rect 198004 546 198056 552
rect 198648 604 198700 610
rect 198648 546 198700 552
rect 196820 480 196848 546
rect 198016 480 198044 546
rect 199212 480 199240 5646
rect 200408 480 200436 9522
rect 202696 5636 202748 5642
rect 202696 5578 202748 5584
rect 201500 4344 201552 4350
rect 201500 4286 201552 4292
rect 201512 480 201540 4286
rect 202708 480 202736 5578
rect 203904 480 203932 9590
rect 207480 8900 207532 8906
rect 207480 8842 207532 8848
rect 206284 5568 206336 5574
rect 206284 5510 206336 5516
rect 205086 4856 205142 4865
rect 205086 4791 205142 4800
rect 205100 480 205128 4791
rect 206296 480 206324 5510
rect 207492 480 207520 8842
rect 210884 8832 210936 8838
rect 210884 8774 210936 8780
rect 209872 6928 209924 6934
rect 209872 6870 209924 6876
rect 208676 4752 208728 4758
rect 208676 4694 208728 4700
rect 208688 480 208716 4694
rect 209884 480 209912 6870
rect 210896 5794 210924 8774
rect 211080 6934 211108 12922
rect 213828 12912 213880 12918
rect 213828 12854 213880 12860
rect 211068 6928 211120 6934
rect 211068 6870 211120 6876
rect 210896 5766 211108 5794
rect 211080 480 211108 5766
rect 212264 4684 212316 4690
rect 212264 4626 212316 4632
rect 212276 480 212304 4626
rect 213840 626 213868 12854
rect 217968 12844 218020 12850
rect 217968 12786 218020 12792
rect 214656 8764 214708 8770
rect 214656 8706 214708 8712
rect 213472 598 213868 626
rect 213472 480 213500 598
rect 214668 480 214696 8706
rect 215852 4616 215904 4622
rect 215852 4558 215904 4564
rect 215864 480 215892 4558
rect 217980 610 218008 12786
rect 220728 12776 220780 12782
rect 220728 12718 220780 12724
rect 218152 8696 218204 8702
rect 218152 8638 218204 8644
rect 217048 604 217100 610
rect 217048 546 217100 552
rect 217968 604 218020 610
rect 217968 546 218020 552
rect 217060 480 217088 546
rect 218164 480 218192 8638
rect 219348 4548 219400 4554
rect 219348 4490 219400 4496
rect 219360 480 219388 4490
rect 220740 610 220768 12718
rect 224868 12708 224920 12714
rect 224868 12650 224920 12656
rect 221740 8628 221792 8634
rect 221740 8570 221792 8576
rect 220544 604 220596 610
rect 220544 546 220596 552
rect 220728 604 220780 610
rect 220728 546 220780 552
rect 220556 480 220584 546
rect 221752 480 221780 8570
rect 222936 4480 222988 4486
rect 222936 4422 222988 4428
rect 222948 480 222976 4422
rect 224880 610 224908 12650
rect 229008 12640 229060 12646
rect 229008 12582 229060 12588
rect 225328 8560 225380 8566
rect 225328 8502 225380 8508
rect 224132 604 224184 610
rect 224132 546 224184 552
rect 224868 604 224920 610
rect 224868 546 224920 552
rect 224144 480 224172 546
rect 225340 480 225368 8502
rect 228916 8492 228968 8498
rect 228916 8434 228968 8440
rect 227720 7608 227772 7614
rect 227720 7550 227772 7556
rect 226524 4412 226576 4418
rect 226524 4354 226576 4360
rect 226536 480 226564 4354
rect 227732 480 227760 7550
rect 228928 480 228956 8434
rect 229020 7614 229048 12582
rect 229008 7608 229060 7614
rect 229008 7550 229060 7556
rect 229112 4282 229140 340054
rect 230124 335594 230152 340054
rect 229296 335566 230152 335594
rect 229296 321570 229324 335566
rect 229284 321564 229336 321570
rect 229284 321506 229336 321512
rect 229468 321564 229520 321570
rect 229468 321506 229520 321512
rect 229480 313954 229508 321506
rect 229468 313948 229520 313954
rect 229468 313890 229520 313896
rect 229652 313948 229704 313954
rect 229652 313890 229704 313896
rect 229664 309126 229692 313890
rect 229468 309120 229520 309126
rect 229468 309062 229520 309068
rect 229652 309120 229704 309126
rect 229652 309062 229704 309068
rect 229480 299606 229508 309062
rect 229468 299600 229520 299606
rect 229468 299542 229520 299548
rect 229284 298172 229336 298178
rect 229284 298114 229336 298120
rect 229296 298058 229324 298114
rect 229374 298072 229430 298081
rect 229296 298030 229374 298058
rect 229374 298007 229430 298016
rect 229558 298072 229614 298081
rect 229558 298007 229614 298016
rect 229572 292466 229600 298007
rect 229376 292460 229428 292466
rect 229376 292402 229428 292408
rect 229560 292460 229612 292466
rect 229560 292402 229612 292408
rect 229388 283014 229416 292402
rect 229376 283008 229428 283014
rect 229376 282950 229428 282956
rect 229376 282804 229428 282810
rect 229376 282746 229428 282752
rect 229388 280158 229416 282746
rect 229376 280152 229428 280158
rect 229376 280094 229428 280100
rect 229376 273148 229428 273154
rect 229376 273090 229428 273096
rect 229388 270502 229416 273090
rect 229376 270496 229428 270502
rect 229376 270438 229428 270444
rect 229376 263492 229428 263498
rect 229376 263434 229428 263440
rect 229388 260846 229416 263434
rect 229376 260840 229428 260846
rect 229376 260782 229428 260788
rect 229376 253836 229428 253842
rect 229376 253778 229428 253784
rect 229388 244390 229416 253778
rect 229376 244384 229428 244390
rect 229376 244326 229428 244332
rect 229284 244248 229336 244254
rect 229284 244190 229336 244196
rect 229296 240145 229324 244190
rect 229282 240136 229338 240145
rect 229282 240071 229338 240080
rect 229558 240136 229614 240145
rect 229558 240071 229614 240080
rect 229572 230518 229600 240071
rect 229376 230512 229428 230518
rect 229376 230454 229428 230460
rect 229560 230512 229612 230518
rect 229560 230454 229612 230460
rect 229388 225078 229416 230454
rect 229376 225072 229428 225078
rect 229376 225014 229428 225020
rect 229284 224936 229336 224942
rect 229284 224878 229336 224884
rect 229296 220794 229324 224878
rect 229284 220788 229336 220794
rect 229284 220730 229336 220736
rect 229284 215280 229336 215286
rect 229284 215222 229336 215228
rect 229296 211154 229324 215222
rect 229296 211126 229416 211154
rect 229388 202910 229416 211126
rect 229284 202904 229336 202910
rect 229282 202872 229284 202881
rect 229376 202904 229428 202910
rect 229336 202872 229338 202881
rect 229376 202846 229428 202852
rect 229558 202872 229614 202881
rect 229282 202807 229338 202816
rect 229558 202807 229614 202816
rect 229572 193254 229600 202807
rect 229376 193248 229428 193254
rect 229376 193190 229428 193196
rect 229560 193248 229612 193254
rect 229560 193190 229612 193196
rect 229388 186266 229416 193190
rect 229296 186238 229416 186266
rect 229296 183569 229324 186238
rect 229282 183560 229338 183569
rect 229282 183495 229338 183504
rect 229558 183560 229614 183569
rect 229558 183495 229614 183504
rect 229572 173942 229600 183495
rect 229376 173936 229428 173942
rect 229376 173878 229428 173884
rect 229560 173936 229612 173942
rect 229560 173878 229612 173884
rect 229388 166954 229416 173878
rect 229296 166926 229416 166954
rect 229296 157418 229324 166926
rect 229284 157412 229336 157418
rect 229284 157354 229336 157360
rect 229376 157344 229428 157350
rect 229376 157286 229428 157292
rect 229388 154562 229416 157286
rect 229376 154556 229428 154562
rect 229376 154498 229428 154504
rect 229560 154556 229612 154562
rect 229560 154498 229612 154504
rect 229572 144945 229600 154498
rect 229282 144936 229338 144945
rect 229282 144871 229338 144880
rect 229558 144936 229614 144945
rect 229558 144871 229614 144880
rect 229296 138038 229324 144871
rect 229284 138032 229336 138038
rect 229284 137974 229336 137980
rect 229376 137964 229428 137970
rect 229376 137906 229428 137912
rect 229388 135250 229416 137906
rect 229376 135244 229428 135250
rect 229376 135186 229428 135192
rect 229560 135244 229612 135250
rect 229560 135186 229612 135192
rect 229572 125633 229600 135186
rect 229282 125624 229338 125633
rect 229282 125559 229338 125568
rect 229558 125624 229614 125633
rect 229558 125559 229614 125568
rect 229296 118726 229324 125559
rect 229284 118720 229336 118726
rect 229284 118662 229336 118668
rect 229376 118652 229428 118658
rect 229376 118594 229428 118600
rect 229388 115938 229416 118594
rect 229376 115932 229428 115938
rect 229376 115874 229428 115880
rect 229284 106344 229336 106350
rect 229284 106286 229336 106292
rect 229296 99414 229324 106286
rect 229284 99408 229336 99414
rect 229284 99350 229336 99356
rect 229376 99340 229428 99346
rect 229376 99282 229428 99288
rect 229388 96626 229416 99282
rect 229376 96620 229428 96626
rect 229376 96562 229428 96568
rect 229284 87032 229336 87038
rect 229284 86974 229336 86980
rect 229296 80102 229324 86974
rect 229284 80096 229336 80102
rect 229284 80038 229336 80044
rect 229376 79960 229428 79966
rect 229376 79902 229428 79908
rect 229388 74526 229416 79902
rect 229376 74520 229428 74526
rect 229376 74462 229428 74468
rect 229284 65000 229336 65006
rect 229284 64942 229336 64948
rect 229296 64870 229324 64942
rect 229284 64864 229336 64870
rect 229284 64806 229336 64812
rect 229468 64864 229520 64870
rect 229468 64806 229520 64812
rect 229480 60602 229508 64806
rect 229388 60574 229508 60602
rect 229388 51134 229416 60574
rect 229376 51128 229428 51134
rect 229376 51070 229428 51076
rect 229284 51060 229336 51066
rect 229284 51002 229336 51008
rect 229296 41478 229324 51002
rect 229284 41472 229336 41478
rect 229284 41414 229336 41420
rect 229376 38752 229428 38758
rect 229296 38700 229376 38706
rect 229296 38694 229428 38700
rect 229296 38678 229416 38694
rect 229296 31822 229324 38678
rect 229284 31816 229336 31822
rect 229284 31758 229336 31764
rect 229376 31680 229428 31686
rect 229376 31622 229428 31628
rect 229388 22273 229416 31622
rect 229374 22264 229430 22273
rect 229374 22199 229430 22208
rect 229374 18048 229430 18057
rect 229374 17983 229430 17992
rect 229388 17950 229416 17983
rect 229376 17944 229428 17950
rect 229376 17886 229428 17892
rect 229192 8356 229244 8362
rect 229192 8298 229244 8304
rect 229204 4894 229232 8298
rect 230492 4894 230520 340054
rect 231044 335730 231072 340054
rect 231780 337385 231808 340068
rect 232148 340054 232254 340082
rect 232424 340054 232714 340082
rect 232792 340054 233174 340082
rect 231766 337376 231822 337385
rect 231766 337311 231822 337320
rect 230584 335702 231072 335730
rect 232044 335708 232096 335714
rect 230584 7585 230612 335702
rect 232044 335650 232096 335656
rect 231952 335640 232004 335646
rect 231952 335582 232004 335588
rect 231308 9716 231360 9722
rect 231308 9658 231360 9664
rect 230570 7576 230626 7585
rect 230570 7511 230626 7520
rect 229192 4888 229244 4894
rect 229192 4830 229244 4836
rect 230480 4888 230532 4894
rect 230480 4830 230532 4836
rect 230112 4820 230164 4826
rect 230112 4762 230164 4768
rect 229100 4276 229152 4282
rect 229100 4218 229152 4224
rect 230124 480 230152 4762
rect 231320 480 231348 9658
rect 231964 5030 231992 335582
rect 232056 6934 232084 335650
rect 232044 6928 232096 6934
rect 232044 6870 232096 6876
rect 231952 5024 232004 5030
rect 231952 4966 232004 4972
rect 232148 3369 232176 340054
rect 232424 335646 232452 340054
rect 232792 335714 232820 340054
rect 233620 337414 233648 340068
rect 233988 337754 234016 340068
rect 234080 340054 234462 340082
rect 233976 337748 234028 337754
rect 233976 337690 234028 337696
rect 233608 337408 233660 337414
rect 233608 337350 233660 337356
rect 232780 335708 232832 335714
rect 232780 335650 232832 335656
rect 232412 335640 232464 335646
rect 232412 335582 232464 335588
rect 234080 334490 234108 340054
rect 234160 337408 234212 337414
rect 234160 337350 234212 337356
rect 234068 334484 234120 334490
rect 234068 334426 234120 334432
rect 234172 334370 234200 337350
rect 234712 335640 234764 335646
rect 234712 335582 234764 335588
rect 233896 334342 234200 334370
rect 233516 328500 233568 328506
rect 233516 328442 233568 328448
rect 233528 302258 233556 328442
rect 233332 302252 233384 302258
rect 233332 302194 233384 302200
rect 233516 302252 233568 302258
rect 233516 302194 233568 302200
rect 233344 302138 233372 302194
rect 233344 302110 233464 302138
rect 233436 292618 233464 302110
rect 233436 292590 233556 292618
rect 233528 282946 233556 292590
rect 233332 282940 233384 282946
rect 233332 282882 233384 282888
rect 233516 282940 233568 282946
rect 233516 282882 233568 282888
rect 233344 282826 233372 282882
rect 233344 282798 233464 282826
rect 233436 273306 233464 282798
rect 233436 273278 233556 273306
rect 233528 263634 233556 273278
rect 233332 263628 233384 263634
rect 233332 263570 233384 263576
rect 233516 263628 233568 263634
rect 233516 263570 233568 263576
rect 233344 263514 233372 263570
rect 233344 263486 233464 263514
rect 233436 253994 233464 263486
rect 233436 253966 233556 253994
rect 233528 244322 233556 253966
rect 233332 244316 233384 244322
rect 233332 244258 233384 244264
rect 233516 244316 233568 244322
rect 233516 244258 233568 244264
rect 233344 244202 233372 244258
rect 233344 244174 233464 244202
rect 233436 234682 233464 244174
rect 233436 234654 233556 234682
rect 233528 225010 233556 234654
rect 233332 225004 233384 225010
rect 233332 224946 233384 224952
rect 233516 225004 233568 225010
rect 233516 224946 233568 224952
rect 233344 224890 233372 224946
rect 233344 224862 233464 224890
rect 233436 215370 233464 224862
rect 233436 215342 233556 215370
rect 233528 205698 233556 215342
rect 233332 205692 233384 205698
rect 233332 205634 233384 205640
rect 233516 205692 233568 205698
rect 233516 205634 233568 205640
rect 233344 205578 233372 205634
rect 233344 205550 233464 205578
rect 233436 196058 233464 205550
rect 233436 196030 233556 196058
rect 233528 186386 233556 196030
rect 233332 186380 233384 186386
rect 233332 186322 233384 186328
rect 233516 186380 233568 186386
rect 233516 186322 233568 186328
rect 233344 186266 233372 186322
rect 233344 186238 233464 186266
rect 233436 183546 233464 186238
rect 233436 183518 233556 183546
rect 233528 167074 233556 183518
rect 233332 167068 233384 167074
rect 233332 167010 233384 167016
rect 233516 167068 233568 167074
rect 233516 167010 233568 167016
rect 233344 166954 233372 167010
rect 233344 166926 233464 166954
rect 233436 159338 233464 166926
rect 233436 159310 233556 159338
rect 233528 147694 233556 159310
rect 233332 147688 233384 147694
rect 233516 147688 233568 147694
rect 233384 147636 233464 147642
rect 233332 147630 233464 147636
rect 233516 147630 233568 147636
rect 233344 147614 233464 147630
rect 233436 132530 233464 147614
rect 233424 132524 233476 132530
rect 233424 132466 233476 132472
rect 233424 131164 233476 131170
rect 233424 131106 233476 131112
rect 233436 125526 233464 131106
rect 233424 125520 233476 125526
rect 233424 125462 233476 125468
rect 233424 121508 233476 121514
rect 233424 121450 233476 121456
rect 233436 118810 233464 121450
rect 233436 118782 233556 118810
rect 233528 104938 233556 118782
rect 233436 104910 233556 104938
rect 233436 100042 233464 104910
rect 233436 100014 233556 100042
rect 233528 89758 233556 100014
rect 233332 89752 233384 89758
rect 233516 89752 233568 89758
rect 233384 89700 233464 89706
rect 233332 89694 233464 89700
rect 233516 89694 233568 89700
rect 233344 89678 233464 89694
rect 233436 77314 233464 89678
rect 233424 77308 233476 77314
rect 233424 77250 233476 77256
rect 233516 77308 233568 77314
rect 233516 77250 233568 77256
rect 233528 64938 233556 77250
rect 233424 64932 233476 64938
rect 233424 64874 233476 64880
rect 233516 64932 233568 64938
rect 233516 64874 233568 64880
rect 233436 60738 233464 64874
rect 233436 60710 233556 60738
rect 233528 51082 233556 60710
rect 233344 51054 233556 51082
rect 233344 50946 233372 51054
rect 233344 50918 233464 50946
rect 233436 31770 233464 50918
rect 233344 31742 233464 31770
rect 233344 12458 233372 31742
rect 233252 12430 233372 12458
rect 232504 8424 232556 8430
rect 232504 8366 232556 8372
rect 232134 3360 232190 3369
rect 232134 3295 232190 3304
rect 232516 480 232544 8366
rect 233252 5098 233280 12430
rect 233896 9042 233924 334342
rect 234618 277400 234674 277409
rect 234618 277335 234674 277344
rect 234632 259486 234660 277335
rect 234620 259480 234672 259486
rect 234620 259422 234672 259428
rect 234724 12510 234752 335582
rect 234908 328522 234936 340068
rect 235000 340054 235382 340082
rect 235460 340054 235842 340082
rect 236196 340054 236302 340082
rect 236472 340054 236762 340082
rect 235000 335646 235028 340054
rect 234988 335640 235040 335646
rect 234988 335582 235040 335588
rect 235460 331974 235488 340054
rect 236092 335640 236144 335646
rect 236092 335582 236144 335588
rect 235448 331968 235500 331974
rect 235448 331910 235500 331916
rect 234816 328494 234936 328522
rect 234816 327078 234844 328494
rect 235080 327140 235132 327146
rect 235080 327082 235132 327088
rect 234804 327072 234856 327078
rect 234804 327014 234856 327020
rect 234896 317484 234948 317490
rect 234896 317426 234948 317432
rect 234908 307766 234936 317426
rect 235092 309126 235120 327082
rect 235080 309120 235132 309126
rect 235080 309062 235132 309068
rect 234896 307760 234948 307766
rect 234896 307702 234948 307708
rect 235080 299532 235132 299538
rect 235080 299474 235132 299480
rect 234896 298172 234948 298178
rect 234896 298114 234948 298120
rect 234908 278746 234936 298114
rect 235092 298110 235120 299474
rect 235080 298104 235132 298110
rect 235080 298046 235132 298052
rect 235080 280220 235132 280226
rect 235080 280162 235132 280168
rect 234816 278718 234936 278746
rect 235092 278730 235120 280162
rect 235080 278724 235132 278730
rect 234816 277409 234844 278718
rect 235080 278666 235132 278672
rect 234802 277400 234858 277409
rect 234802 277335 234858 277344
rect 235080 260908 235132 260914
rect 235080 260850 235132 260856
rect 234896 259480 234948 259486
rect 234896 259422 234948 259428
rect 234908 251258 234936 259422
rect 235092 259418 235120 260850
rect 235080 259412 235132 259418
rect 235080 259354 235132 259360
rect 234896 251252 234948 251258
rect 234896 251194 234948 251200
rect 234988 251116 235040 251122
rect 234988 251058 235040 251064
rect 235000 241534 235028 251058
rect 234896 241528 234948 241534
rect 234896 241470 234948 241476
rect 234988 241528 235040 241534
rect 234988 241470 235040 241476
rect 235080 241528 235132 241534
rect 235080 241470 235132 241476
rect 234908 240106 234936 241470
rect 235092 240145 235120 241470
rect 235078 240136 235134 240145
rect 234896 240100 234948 240106
rect 235078 240071 235134 240080
rect 235262 240136 235318 240145
rect 235262 240071 235318 240080
rect 234896 240042 234948 240048
rect 235276 230518 235304 240071
rect 234896 230512 234948 230518
rect 234896 230454 234948 230460
rect 235080 230512 235132 230518
rect 235080 230454 235132 230460
rect 235264 230512 235316 230518
rect 235264 230454 235316 230460
rect 234908 220833 234936 230454
rect 235092 222358 235120 230454
rect 235080 222352 235132 222358
rect 235080 222294 235132 222300
rect 235080 222216 235132 222222
rect 235080 222158 235132 222164
rect 234894 220824 234950 220833
rect 235092 220794 235120 222158
rect 235170 220824 235226 220833
rect 234894 220759 234950 220768
rect 235080 220788 235132 220794
rect 235170 220759 235226 220768
rect 235080 220730 235132 220736
rect 235080 211200 235132 211206
rect 234894 211168 234950 211177
rect 235184 211177 235212 220759
rect 235080 211142 235132 211148
rect 235170 211168 235226 211177
rect 234894 211103 234950 211112
rect 234908 202910 234936 211103
rect 235092 205850 235120 211142
rect 235170 211103 235226 211112
rect 235000 205822 235120 205850
rect 235000 205578 235028 205822
rect 235000 205550 235120 205578
rect 234804 202904 234856 202910
rect 234804 202846 234856 202852
rect 234896 202904 234948 202910
rect 234896 202846 234948 202852
rect 234816 201482 234844 202846
rect 234804 201476 234856 201482
rect 234804 201418 234856 201424
rect 235092 193254 235120 205550
rect 235080 193248 235132 193254
rect 235080 193190 235132 193196
rect 235264 193180 235316 193186
rect 235264 193122 235316 193128
rect 234804 192296 234856 192302
rect 234804 192238 234856 192244
rect 234816 173942 234844 192238
rect 235276 183598 235304 193122
rect 234988 183592 235040 183598
rect 234988 183534 235040 183540
rect 235264 183592 235316 183598
rect 235264 183534 235316 183540
rect 235000 179382 235028 183534
rect 234988 179376 235040 179382
rect 234988 179318 235040 179324
rect 235172 179376 235224 179382
rect 235172 179318 235224 179324
rect 234804 173936 234856 173942
rect 234804 173878 234856 173884
rect 234896 173936 234948 173942
rect 234948 173884 235028 173890
rect 234896 173878 235028 173884
rect 234908 173862 235028 173878
rect 235000 163146 235028 173862
rect 235000 163118 235120 163146
rect 234988 162988 235040 162994
rect 234988 162930 235040 162936
rect 234894 162888 234950 162897
rect 234894 162823 234950 162832
rect 234908 161362 234936 162823
rect 235000 161430 235028 162930
rect 235092 162897 235120 163118
rect 235184 162994 235212 179318
rect 235172 162988 235224 162994
rect 235172 162930 235224 162936
rect 235078 162888 235134 162897
rect 235078 162823 235134 162832
rect 234988 161424 235040 161430
rect 234988 161366 235040 161372
rect 234896 161356 234948 161362
rect 234896 161298 234948 161304
rect 235080 151836 235132 151842
rect 235080 151778 235132 151784
rect 235092 143721 235120 151778
rect 235078 143712 235134 143721
rect 235078 143647 235134 143656
rect 235170 143576 235226 143585
rect 235170 143511 235226 143520
rect 234804 140888 234856 140894
rect 234804 140830 234856 140836
rect 234816 140758 234844 140830
rect 234804 140752 234856 140758
rect 234804 140694 234856 140700
rect 234988 134632 235040 134638
rect 234988 134574 235040 134580
rect 235000 121530 235028 134574
rect 235184 132546 235212 143511
rect 235092 132518 235212 132546
rect 235092 128382 235120 132518
rect 235080 128376 235132 128382
rect 235080 128318 235132 128324
rect 235080 122868 235132 122874
rect 235080 122810 235132 122816
rect 234908 121502 235028 121530
rect 234908 120086 234936 121502
rect 234896 120080 234948 120086
rect 234896 120022 234948 120028
rect 235092 114510 235120 122810
rect 234988 114504 235040 114510
rect 234988 114446 235040 114452
rect 235080 114504 235132 114510
rect 235080 114446 235132 114452
rect 235000 104854 235028 114446
rect 234988 104848 235040 104854
rect 234988 104790 235040 104796
rect 235080 104848 235132 104854
rect 235080 104790 235132 104796
rect 234804 92064 234856 92070
rect 234804 92006 234856 92012
rect 234816 85785 234844 92006
rect 234802 85776 234858 85785
rect 234802 85711 234858 85720
rect 234802 85640 234858 85649
rect 234802 85575 234858 85584
rect 234816 84182 234844 85575
rect 234804 84176 234856 84182
rect 234804 84118 234856 84124
rect 235092 77314 235120 104790
rect 234988 77308 235040 77314
rect 234988 77250 235040 77256
rect 235080 77308 235132 77314
rect 235080 77250 235132 77256
rect 234804 74588 234856 74594
rect 234804 74530 234856 74536
rect 234816 64870 234844 74530
rect 234804 64864 234856 64870
rect 234804 64806 234856 64812
rect 234804 55276 234856 55282
rect 234804 55218 234856 55224
rect 234816 45558 234844 55218
rect 235000 53122 235028 77250
rect 235000 53094 235212 53122
rect 235184 45558 235212 53094
rect 234804 45552 234856 45558
rect 234804 45494 234856 45500
rect 234988 45552 235040 45558
rect 234988 45494 235040 45500
rect 235172 45552 235224 45558
rect 235172 45494 235224 45500
rect 235000 35986 235028 45494
rect 234804 35964 234856 35970
rect 235000 35958 235120 35986
rect 234804 35906 234856 35912
rect 234816 26246 234844 35906
rect 235092 26246 235120 35958
rect 234804 26240 234856 26246
rect 234804 26182 234856 26188
rect 235080 26240 235132 26246
rect 235080 26182 235132 26188
rect 234896 16652 234948 16658
rect 234896 16594 234948 16600
rect 234712 12504 234764 12510
rect 234712 12446 234764 12452
rect 234712 11212 234764 11218
rect 234712 11154 234764 11160
rect 233884 9036 233936 9042
rect 233884 8978 233936 8984
rect 233240 5092 233292 5098
rect 233240 5034 233292 5040
rect 233700 4888 233752 4894
rect 233700 4830 233752 4836
rect 233712 480 233740 4830
rect 234724 3466 234752 11154
rect 234908 8362 234936 16594
rect 236104 11762 236132 335582
rect 236092 11756 236144 11762
rect 236092 11698 236144 11704
rect 236000 8968 236052 8974
rect 236000 8910 236052 8916
rect 234896 8356 234948 8362
rect 234896 8298 234948 8304
rect 235080 8356 235132 8362
rect 235080 8298 235132 8304
rect 234804 7608 234856 7614
rect 234804 7550 234856 7556
rect 234712 3460 234764 3466
rect 234712 3402 234764 3408
rect 234816 480 234844 7550
rect 235092 3534 235120 8298
rect 235080 3528 235132 3534
rect 235080 3470 235132 3476
rect 236012 480 236040 8910
rect 236196 7682 236224 340054
rect 236472 335646 236500 340054
rect 237208 337482 237236 340068
rect 237576 337550 237604 340068
rect 237668 340054 238050 340082
rect 238128 340054 238510 340082
rect 237564 337544 237616 337550
rect 237564 337486 237616 337492
rect 237196 337476 237248 337482
rect 237196 337418 237248 337424
rect 236460 335640 236512 335646
rect 236460 335582 236512 335588
rect 237472 335640 237524 335646
rect 237472 335582 237524 335588
rect 237484 13122 237512 335582
rect 237472 13116 237524 13122
rect 237472 13058 237524 13064
rect 237668 7750 237696 340054
rect 238128 335646 238156 340054
rect 238116 335640 238168 335646
rect 238116 335582 238168 335588
rect 238668 333328 238720 333334
rect 238668 333270 238720 333276
rect 238680 330834 238708 333270
rect 238956 331242 238984 340068
rect 239048 340054 239430 340082
rect 239048 333334 239076 340054
rect 239876 338162 239904 340068
rect 239128 338156 239180 338162
rect 239128 338098 239180 338104
rect 239864 338156 239916 338162
rect 239864 338098 239916 338104
rect 239140 336734 239168 338098
rect 240336 337414 240364 340068
rect 240796 337618 240824 340068
rect 240888 340054 241178 340082
rect 241638 340054 241744 340082
rect 240784 337612 240836 337618
rect 240784 337554 240836 337560
rect 240324 337408 240376 337414
rect 240324 337350 240376 337356
rect 239128 336728 239180 336734
rect 239128 336670 239180 336676
rect 239036 333328 239088 333334
rect 239036 333270 239088 333276
rect 238772 331214 238984 331242
rect 238772 330970 238800 331214
rect 238772 330942 238892 330970
rect 238680 330806 238800 330834
rect 238772 321570 238800 330806
rect 238760 321564 238812 321570
rect 238760 321506 238812 321512
rect 238864 309806 238892 330942
rect 240888 327146 240916 340054
rect 241520 335640 241572 335646
rect 241520 335582 241572 335588
rect 240416 327140 240468 327146
rect 240416 327082 240468 327088
rect 240876 327140 240928 327146
rect 240876 327082 240928 327088
rect 238944 321564 238996 321570
rect 238944 321506 238996 321512
rect 238852 309800 238904 309806
rect 238852 309742 238904 309748
rect 238852 309664 238904 309670
rect 238852 309606 238904 309612
rect 238760 204604 238812 204610
rect 238760 204546 238812 204552
rect 238772 198370 238800 204546
rect 238864 198490 238892 309606
rect 238956 204610 238984 321506
rect 239128 318844 239180 318850
rect 239128 318786 239180 318792
rect 239140 298110 239168 318786
rect 240428 298110 240456 327082
rect 239036 298104 239088 298110
rect 239036 298046 239088 298052
rect 239128 298104 239180 298110
rect 239128 298046 239180 298052
rect 240416 298104 240468 298110
rect 240416 298046 240468 298052
rect 239048 296721 239076 298046
rect 239034 296712 239090 296721
rect 239034 296647 239090 296656
rect 239310 296712 239366 296721
rect 239310 296647 239366 296656
rect 239324 278798 239352 296647
rect 240416 288448 240468 288454
rect 240416 288390 240468 288396
rect 239128 278792 239180 278798
rect 239128 278734 239180 278740
rect 239312 278792 239364 278798
rect 240428 278769 240456 288390
rect 239312 278734 239364 278740
rect 240230 278760 240286 278769
rect 239140 274106 239168 278734
rect 240230 278695 240286 278704
rect 240414 278760 240470 278769
rect 240414 278695 240470 278704
rect 239128 274100 239180 274106
rect 239128 274042 239180 274048
rect 240244 269142 240272 278695
rect 240232 269136 240284 269142
rect 240232 269078 240284 269084
rect 240416 269136 240468 269142
rect 240416 269078 240468 269084
rect 239312 267776 239364 267782
rect 239312 267718 239364 267724
rect 239140 259486 239168 259517
rect 239324 259486 239352 267718
rect 239128 259480 239180 259486
rect 239312 259480 239364 259486
rect 239180 259428 239260 259434
rect 239128 259422 239260 259428
rect 240428 259457 240456 269078
rect 239312 259422 239364 259428
rect 240230 259448 240286 259457
rect 239140 259406 239260 259422
rect 239232 249898 239260 259406
rect 240230 259383 240286 259392
rect 240414 259448 240470 259457
rect 240414 259383 240470 259392
rect 239220 249892 239272 249898
rect 239220 249834 239272 249840
rect 240244 249830 240272 259383
rect 240232 249824 240284 249830
rect 240232 249766 240284 249772
rect 240416 249824 240468 249830
rect 240416 249766 240468 249772
rect 239128 240168 239180 240174
rect 239126 240136 239128 240145
rect 240428 240145 240456 249766
rect 239180 240136 239182 240145
rect 239126 240071 239182 240080
rect 240230 240136 240286 240145
rect 240230 240071 240286 240080
rect 240414 240136 240470 240145
rect 240414 240071 240470 240080
rect 239218 240000 239274 240009
rect 239218 239935 239274 239944
rect 239232 220862 239260 239935
rect 240244 230518 240272 240071
rect 240232 230512 240284 230518
rect 240232 230454 240284 230460
rect 240416 230512 240468 230518
rect 240416 230454 240468 230460
rect 239128 220856 239180 220862
rect 239126 220824 239128 220833
rect 239220 220856 239272 220862
rect 239180 220824 239182 220833
rect 240428 220833 240456 230454
rect 239220 220798 239272 220804
rect 240230 220824 240286 220833
rect 239126 220759 239182 220768
rect 240230 220759 240286 220768
rect 240414 220824 240470 220833
rect 240414 220759 240470 220768
rect 239034 220688 239090 220697
rect 239034 220623 239090 220632
rect 239048 211274 239076 220623
rect 239036 211268 239088 211274
rect 239036 211210 239088 211216
rect 239128 211268 239180 211274
rect 239128 211210 239180 211216
rect 239140 211138 239168 211210
rect 240244 211177 240272 220759
rect 240230 211168 240286 211177
rect 239128 211132 239180 211138
rect 240230 211103 240286 211112
rect 240414 211168 240470 211177
rect 240414 211103 240470 211112
rect 239128 211074 239180 211080
rect 238944 204604 238996 204610
rect 238944 204546 238996 204552
rect 239128 202836 239180 202842
rect 239128 202778 239180 202784
rect 238852 198484 238904 198490
rect 238852 198426 238904 198432
rect 238772 198342 238984 198370
rect 238852 198076 238904 198082
rect 238852 198018 238904 198024
rect 238760 186380 238812 186386
rect 238760 186322 238812 186328
rect 238772 176662 238800 186322
rect 238760 176656 238812 176662
rect 238760 176598 238812 176604
rect 238760 167068 238812 167074
rect 238760 167010 238812 167016
rect 238772 159610 238800 167010
rect 238864 159730 238892 198018
rect 238956 186386 238984 198342
rect 239140 193254 239168 202778
rect 240428 201482 240456 211103
rect 240416 201476 240468 201482
rect 240416 201418 240468 201424
rect 239128 193248 239180 193254
rect 239128 193190 239180 193196
rect 239220 193180 239272 193186
rect 239220 193122 239272 193128
rect 240508 193180 240560 193186
rect 240508 193122 240560 193128
rect 238944 186380 238996 186386
rect 238944 186322 238996 186328
rect 239232 183598 239260 193122
rect 239128 183592 239180 183598
rect 239128 183534 239180 183540
rect 239220 183592 239272 183598
rect 239220 183534 239272 183540
rect 239140 182170 239168 183534
rect 239128 182164 239180 182170
rect 239128 182106 239180 182112
rect 238944 176656 238996 176662
rect 238944 176598 238996 176604
rect 238956 167074 238984 176598
rect 240520 173942 240548 193122
rect 240416 173936 240468 173942
rect 240414 173904 240416 173913
rect 240508 173936 240560 173942
rect 240468 173904 240470 173913
rect 239128 173868 239180 173874
rect 240508 173878 240560 173884
rect 240598 173904 240654 173913
rect 240414 173839 240470 173848
rect 240598 173839 240654 173848
rect 239128 173810 239180 173816
rect 239140 169114 239168 173810
rect 239128 169108 239180 169114
rect 239128 169050 239180 169056
rect 239312 169108 239364 169114
rect 239312 169050 239364 169056
rect 238944 167068 238996 167074
rect 238944 167010 238996 167016
rect 239324 164257 239352 169050
rect 239126 164248 239182 164257
rect 239126 164183 239182 164192
rect 239310 164248 239366 164257
rect 240612 164234 240640 173839
rect 239310 164183 239366 164192
rect 240520 164206 240640 164234
rect 238852 159724 238904 159730
rect 238852 159666 238904 159672
rect 238772 159582 238984 159610
rect 238852 159384 238904 159390
rect 238852 159326 238904 159332
rect 238864 147762 238892 159326
rect 238956 147830 238984 159582
rect 239140 154698 239168 164183
rect 239128 154692 239180 154698
rect 239128 154634 239180 154640
rect 240520 154630 240548 164206
rect 240508 154624 240560 154630
rect 240508 154566 240560 154572
rect 240416 153332 240468 153338
rect 240416 153274 240468 153280
rect 240428 153202 240456 153274
rect 240416 153196 240468 153202
rect 240416 153138 240468 153144
rect 239036 151836 239088 151842
rect 239036 151778 239088 151784
rect 238944 147824 238996 147830
rect 238944 147766 238996 147772
rect 238852 147756 238904 147762
rect 238852 147698 238904 147704
rect 238852 147620 238904 147626
rect 238852 147562 238904 147568
rect 238944 147620 238996 147626
rect 238944 147562 238996 147568
rect 238760 143540 238812 143546
rect 238760 143482 238812 143488
rect 238772 128314 238800 143482
rect 238760 128308 238812 128314
rect 238760 128250 238812 128256
rect 238760 109064 238812 109070
rect 238760 109006 238812 109012
rect 238666 32600 238722 32609
rect 238666 32535 238722 32544
rect 238680 29209 238708 32535
rect 238666 29200 238722 29209
rect 238666 29135 238722 29144
rect 237656 7744 237708 7750
rect 237656 7686 237708 7692
rect 236184 7676 236236 7682
rect 236184 7618 236236 7624
rect 238392 7676 238444 7682
rect 238392 7618 238444 7624
rect 237196 4956 237248 4962
rect 237196 4898 237248 4904
rect 237208 480 237236 4898
rect 238404 480 238432 7618
rect 238772 3670 238800 109006
rect 238760 3664 238812 3670
rect 238760 3606 238812 3612
rect 238864 3602 238892 147562
rect 238956 143546 238984 147562
rect 239048 143546 239076 151778
rect 240324 143608 240376 143614
rect 240324 143550 240376 143556
rect 238944 143540 238996 143546
rect 238944 143482 238996 143488
rect 239036 143540 239088 143546
rect 239036 143482 239088 143488
rect 239128 143540 239180 143546
rect 239128 143482 239180 143488
rect 239140 142118 239168 143482
rect 240336 142118 240364 143550
rect 239128 142112 239180 142118
rect 239128 142054 239180 142060
rect 240324 142112 240376 142118
rect 240324 142054 240376 142060
rect 239128 132524 239180 132530
rect 239128 132466 239180 132472
rect 240416 132524 240468 132530
rect 240416 132466 240468 132472
rect 238944 128308 238996 128314
rect 238944 128250 238996 128256
rect 238956 109070 238984 128250
rect 239140 109138 239168 132466
rect 240428 122806 240456 132466
rect 240416 122800 240468 122806
rect 240416 122742 240468 122748
rect 239128 109132 239180 109138
rect 239128 109074 239180 109080
rect 238944 109064 238996 109070
rect 238944 109006 238996 109012
rect 238944 108928 238996 108934
rect 238944 108870 238996 108876
rect 238956 100094 238984 108870
rect 240324 104916 240376 104922
rect 240324 104858 240376 104864
rect 240336 104802 240364 104858
rect 240336 104774 240548 104802
rect 238944 100088 238996 100094
rect 238944 100030 238996 100036
rect 239128 100088 239180 100094
rect 239128 100030 239180 100036
rect 239140 57934 239168 100030
rect 240520 99226 240548 104774
rect 240428 99198 240548 99226
rect 240428 95198 240456 99198
rect 240416 95192 240468 95198
rect 240416 95134 240468 95140
rect 240508 95192 240560 95198
rect 240508 95134 240560 95140
rect 240520 93838 240548 95134
rect 240508 93832 240560 93838
rect 240508 93774 240560 93780
rect 240046 91216 240102 91225
rect 240046 91151 240102 91160
rect 240060 87145 240088 91151
rect 240046 87136 240102 87145
rect 240046 87071 240102 87080
rect 240416 84244 240468 84250
rect 240416 84186 240468 84192
rect 240428 75886 240456 84186
rect 240416 75880 240468 75886
rect 240416 75822 240468 75828
rect 240416 66360 240468 66366
rect 240416 66302 240468 66308
rect 240428 64870 240456 66302
rect 240416 64864 240468 64870
rect 240416 64806 240468 64812
rect 239128 57928 239180 57934
rect 239128 57870 239180 57876
rect 240324 55276 240376 55282
rect 240324 55218 240376 55224
rect 239036 51060 239088 51066
rect 239036 51002 239088 51008
rect 239048 48278 239076 51002
rect 240336 48346 240364 55218
rect 240324 48340 240376 48346
rect 240324 48282 240376 48288
rect 240416 48340 240468 48346
rect 240416 48282 240468 48288
rect 239036 48272 239088 48278
rect 239036 48214 239088 48220
rect 239128 48272 239180 48278
rect 239128 48214 239180 48220
rect 239140 26246 239168 48214
rect 239128 26240 239180 26246
rect 239128 26182 239180 26188
rect 240428 18193 240456 48282
rect 240414 18184 240470 18193
rect 240414 18119 240470 18128
rect 240322 18048 240378 18057
rect 240322 17983 240378 17992
rect 240336 17950 240364 17983
rect 240324 17944 240376 17950
rect 240324 17886 240376 17892
rect 239588 9036 239640 9042
rect 239588 8978 239640 8984
rect 239036 8356 239088 8362
rect 239036 8298 239088 8304
rect 239048 7818 239076 8298
rect 239036 7812 239088 7818
rect 239036 7754 239088 7760
rect 238852 3596 238904 3602
rect 238852 3538 238904 3544
rect 239600 480 239628 8978
rect 240232 8356 240284 8362
rect 240232 8298 240284 8304
rect 240244 7886 240272 8298
rect 240232 7880 240284 7886
rect 240232 7822 240284 7828
rect 240784 5024 240836 5030
rect 240784 4966 240836 4972
rect 240796 480 240824 4966
rect 241532 3738 241560 335582
rect 241612 111104 241664 111110
rect 241612 111046 241664 111052
rect 241624 106321 241652 111046
rect 241610 106312 241666 106321
rect 241610 106247 241666 106256
rect 241610 18048 241666 18057
rect 241610 17983 241666 17992
rect 241624 17950 241652 17983
rect 241612 17944 241664 17950
rect 241612 17886 241664 17892
rect 241716 14482 241744 340054
rect 241808 340054 242098 340082
rect 242176 340054 242558 340082
rect 241808 335646 241836 340054
rect 241796 335640 241848 335646
rect 241796 335582 241848 335588
rect 242176 327146 242204 340054
rect 243004 337822 243032 340068
rect 242992 337816 243044 337822
rect 242992 337758 243044 337764
rect 243464 337686 243492 340068
rect 243556 340054 243938 340082
rect 243452 337680 243504 337686
rect 243452 337622 243504 337628
rect 243556 335696 243584 340054
rect 243096 335668 243584 335696
rect 241888 327140 241940 327146
rect 241888 327082 241940 327088
rect 242164 327140 242216 327146
rect 242164 327082 242216 327088
rect 241900 298110 241928 327082
rect 241888 298104 241940 298110
rect 241888 298046 241940 298052
rect 241888 288448 241940 288454
rect 241888 288390 241940 288396
rect 241900 278769 241928 288390
rect 241886 278760 241942 278769
rect 241886 278695 241942 278704
rect 242070 278760 242126 278769
rect 242070 278695 242126 278704
rect 242084 269142 242112 278695
rect 241888 269136 241940 269142
rect 241888 269078 241940 269084
rect 242072 269136 242124 269142
rect 242072 269078 242124 269084
rect 241900 259457 241928 269078
rect 241886 259448 241942 259457
rect 241886 259383 241942 259392
rect 242070 259448 242126 259457
rect 242070 259383 242126 259392
rect 242084 249830 242112 259383
rect 241888 249824 241940 249830
rect 241888 249766 241940 249772
rect 242072 249824 242124 249830
rect 242072 249766 242124 249772
rect 241900 240145 241928 249766
rect 241886 240136 241942 240145
rect 241886 240071 241942 240080
rect 242070 240136 242126 240145
rect 242070 240071 242126 240080
rect 242084 230518 242112 240071
rect 241888 230512 241940 230518
rect 241888 230454 241940 230460
rect 242072 230512 242124 230518
rect 242072 230454 242124 230460
rect 241900 220833 241928 230454
rect 241886 220824 241942 220833
rect 241886 220759 241942 220768
rect 242070 220824 242126 220833
rect 242070 220759 242126 220768
rect 242084 211177 242112 220759
rect 241886 211168 241942 211177
rect 241886 211103 241942 211112
rect 242070 211168 242126 211177
rect 242070 211103 242126 211112
rect 241900 183666 241928 211103
rect 241888 183660 241940 183666
rect 241888 183602 241940 183608
rect 241796 183592 241848 183598
rect 241796 183534 241848 183540
rect 241808 178838 241836 183534
rect 241796 178832 241848 178838
rect 241796 178774 241848 178780
rect 241796 173936 241848 173942
rect 241796 173878 241848 173884
rect 241808 164234 241836 173878
rect 241808 164206 241928 164234
rect 241900 162858 241928 164206
rect 241888 162852 241940 162858
rect 241888 162794 241940 162800
rect 241888 153264 241940 153270
rect 241888 153206 241940 153212
rect 241900 147642 241928 153206
rect 241808 147614 241928 147642
rect 241808 144906 241836 147614
rect 241796 144900 241848 144906
rect 241796 144842 241848 144848
rect 241980 144900 242032 144906
rect 241980 144842 242032 144848
rect 241992 135266 242020 144842
rect 241900 135250 242020 135266
rect 241888 135244 242020 135250
rect 241940 135238 242020 135244
rect 241888 135186 241940 135192
rect 241900 135155 241928 135186
rect 241888 125656 241940 125662
rect 241888 125598 241940 125604
rect 241900 124166 241928 125598
rect 241888 124160 241940 124166
rect 241888 124102 241940 124108
rect 241888 114572 241940 114578
rect 241888 114514 241940 114520
rect 241900 111110 241928 114514
rect 241888 111104 241940 111110
rect 241888 111046 241940 111052
rect 241794 106312 241850 106321
rect 241794 106247 241850 106256
rect 241808 104854 241836 106247
rect 241796 104848 241848 104854
rect 241796 104790 241848 104796
rect 241888 95260 241940 95266
rect 241888 95202 241940 95208
rect 241900 57882 241928 95202
rect 241808 57854 241928 57882
rect 241808 50402 241836 57854
rect 241808 50374 241928 50402
rect 241900 45642 241928 50374
rect 241808 45614 241928 45642
rect 241808 44130 241836 45614
rect 241796 44124 241848 44130
rect 241796 44066 241848 44072
rect 241796 29028 241848 29034
rect 241796 28970 241848 28976
rect 241808 18193 241836 28970
rect 241794 18184 241850 18193
rect 241794 18119 241850 18128
rect 241704 14476 241756 14482
rect 241704 14418 241756 14424
rect 241704 8356 241756 8362
rect 241704 8298 241756 8304
rect 241716 7954 241744 8298
rect 243096 8022 243124 335668
rect 244384 331294 244412 340068
rect 244476 340054 244858 340082
rect 244936 340054 245226 340082
rect 244476 331362 244504 340054
rect 244936 331786 244964 340054
rect 245672 337958 245700 340068
rect 245660 337952 245712 337958
rect 245660 337894 245712 337900
rect 246132 337890 246160 340068
rect 246224 340054 246606 340082
rect 246120 337884 246172 337890
rect 246120 337826 246172 337832
rect 244568 331758 244964 331786
rect 244464 331356 244516 331362
rect 244464 331298 244516 331304
rect 244372 331288 244424 331294
rect 244372 331230 244424 331236
rect 244280 331220 244332 331226
rect 244280 331162 244332 331168
rect 244292 309074 244320 331162
rect 244372 331152 244424 331158
rect 244372 331094 244424 331100
rect 244200 309046 244320 309074
rect 244200 299606 244228 309046
rect 244188 299600 244240 299606
rect 244188 299542 244240 299548
rect 244280 299532 244332 299538
rect 244280 299474 244332 299480
rect 244292 270502 244320 299474
rect 244280 270496 244332 270502
rect 244280 270438 244332 270444
rect 244280 260908 244332 260914
rect 244280 260850 244332 260856
rect 244292 251190 244320 260850
rect 244280 251184 244332 251190
rect 244280 251126 244332 251132
rect 244280 241528 244332 241534
rect 244280 241470 244332 241476
rect 244292 231826 244320 241470
rect 244200 231798 244320 231826
rect 244200 222222 244228 231798
rect 244188 222216 244240 222222
rect 244188 222158 244240 222164
rect 244280 222216 244332 222222
rect 244280 222158 244332 222164
rect 244292 202881 244320 222158
rect 244094 202872 244150 202881
rect 244094 202807 244150 202816
rect 244278 202872 244334 202881
rect 244278 202807 244334 202816
rect 244108 193254 244136 202807
rect 244096 193248 244148 193254
rect 244096 193190 244148 193196
rect 244280 193248 244332 193254
rect 244280 193190 244332 193196
rect 244292 189446 244320 193190
rect 244280 189440 244332 189446
rect 244280 189382 244332 189388
rect 244280 173936 244332 173942
rect 244280 173878 244332 173884
rect 244292 144906 244320 173878
rect 244096 144900 244148 144906
rect 244096 144842 244148 144848
rect 244280 144900 244332 144906
rect 244280 144842 244332 144848
rect 244108 135289 244136 144842
rect 244094 135280 244150 135289
rect 244094 135215 244150 135224
rect 244278 135280 244334 135289
rect 244278 135215 244334 135224
rect 244292 67590 244320 135215
rect 244280 67584 244332 67590
rect 244280 67526 244332 67532
rect 244280 57996 244332 58002
rect 244280 57938 244332 57944
rect 243176 8356 243228 8362
rect 243176 8298 243228 8304
rect 243084 8016 243136 8022
rect 243084 7958 243136 7964
rect 241704 7948 241756 7954
rect 241704 7890 241756 7896
rect 241980 7744 242032 7750
rect 241980 7686 242032 7692
rect 241520 3732 241572 3738
rect 241520 3674 241572 3680
rect 241992 480 242020 7686
rect 243188 480 243216 8298
rect 244292 3874 244320 57938
rect 244384 5250 244412 331094
rect 244568 316690 244596 331758
rect 246224 327146 246252 340054
rect 247052 337278 247080 340068
rect 247236 340054 247526 340082
rect 247696 340054 247986 340082
rect 248446 340054 248552 340082
rect 246304 337272 246356 337278
rect 246304 337214 246356 337220
rect 247040 337272 247092 337278
rect 247040 337214 247092 337220
rect 245936 327140 245988 327146
rect 245936 327082 245988 327088
rect 246212 327140 246264 327146
rect 246212 327082 246264 327088
rect 244476 316662 244596 316690
rect 244476 307034 244504 316662
rect 244476 307006 244596 307034
rect 244568 297378 244596 307006
rect 244476 297350 244596 297378
rect 244476 287722 244504 297350
rect 244476 287694 244596 287722
rect 244568 277794 244596 287694
rect 244476 277766 244596 277794
rect 244476 270586 244504 277766
rect 244476 270558 244596 270586
rect 244568 258482 244596 270558
rect 245948 270502 245976 327082
rect 245936 270496 245988 270502
rect 245936 270438 245988 270444
rect 245936 260908 245988 260914
rect 245936 260850 245988 260856
rect 244476 258454 244596 258482
rect 244476 251274 244504 258454
rect 244476 251246 244596 251274
rect 244568 239442 244596 251246
rect 245948 251190 245976 260850
rect 245936 251184 245988 251190
rect 245936 251126 245988 251132
rect 245936 241528 245988 241534
rect 245936 241470 245988 241476
rect 244476 239414 244596 239442
rect 244476 231810 244504 239414
rect 245948 231849 245976 241470
rect 245750 231840 245806 231849
rect 244464 231804 244516 231810
rect 244464 231746 244516 231752
rect 244556 231804 244608 231810
rect 245750 231775 245806 231784
rect 245934 231840 245990 231849
rect 245934 231775 245990 231784
rect 244556 231746 244608 231752
rect 244568 217954 244596 231746
rect 245764 222222 245792 231775
rect 245752 222216 245804 222222
rect 245752 222158 245804 222164
rect 245936 222216 245988 222222
rect 245936 222158 245988 222164
rect 244476 217926 244596 217954
rect 244476 210746 244504 217926
rect 244476 210718 244596 210746
rect 244568 198642 244596 210718
rect 244476 198614 244596 198642
rect 244476 191434 244504 198614
rect 244476 191406 244596 191434
rect 244464 189440 244516 189446
rect 244464 189382 244516 189388
rect 244476 173942 244504 189382
rect 244464 173936 244516 173942
rect 244464 173878 244516 173884
rect 244568 162194 244596 191406
rect 244476 162166 244596 162194
rect 244476 152538 244504 162166
rect 245948 154562 245976 222158
rect 245752 154556 245804 154562
rect 245752 154498 245804 154504
rect 245936 154556 245988 154562
rect 245936 154498 245988 154504
rect 244476 152510 244596 152538
rect 244568 123570 244596 152510
rect 245764 144945 245792 154498
rect 245750 144936 245806 144945
rect 245750 144871 245806 144880
rect 245934 144936 245990 144945
rect 245934 144871 245990 144880
rect 245948 135250 245976 144871
rect 245752 135244 245804 135250
rect 245752 135186 245804 135192
rect 245936 135244 245988 135250
rect 245936 135186 245988 135192
rect 245764 125633 245792 135186
rect 245750 125624 245806 125633
rect 245750 125559 245806 125568
rect 245934 125624 245990 125633
rect 245934 125559 245990 125568
rect 244476 123542 244596 123570
rect 244476 113914 244504 123542
rect 245948 115938 245976 125559
rect 245936 115932 245988 115938
rect 245936 115874 245988 115880
rect 244476 113886 244596 113914
rect 244568 104258 244596 113886
rect 245936 106344 245988 106350
rect 245936 106286 245988 106292
rect 244476 104230 244596 104258
rect 244476 94654 244504 104230
rect 244464 94648 244516 94654
rect 244464 94590 244516 94596
rect 244464 85604 244516 85610
rect 244464 85546 244516 85552
rect 244476 77314 244504 85546
rect 244464 77308 244516 77314
rect 244464 77250 244516 77256
rect 244556 77308 244608 77314
rect 244556 77250 244608 77256
rect 244568 75886 244596 77250
rect 244464 75880 244516 75886
rect 244464 75822 244516 75828
rect 244556 75880 244608 75886
rect 244556 75822 244608 75828
rect 244476 55842 244504 75822
rect 245948 57934 245976 106286
rect 245936 57928 245988 57934
rect 245936 57870 245988 57876
rect 244476 55814 244596 55842
rect 244568 19446 244596 55814
rect 245936 48340 245988 48346
rect 245936 48282 245988 48288
rect 245948 38622 245976 48282
rect 245936 38616 245988 38622
rect 245936 38558 245988 38564
rect 245936 29028 245988 29034
rect 245936 28970 245988 28976
rect 245948 22166 245976 28970
rect 245936 22160 245988 22166
rect 245936 22102 245988 22108
rect 245752 22092 245804 22098
rect 245752 22034 245804 22040
rect 244556 19440 244608 19446
rect 244556 19382 244608 19388
rect 244464 19372 244516 19378
rect 244464 19314 244516 19320
rect 244476 9110 244504 19314
rect 245764 9178 245792 22034
rect 245752 9172 245804 9178
rect 245752 9114 245804 9120
rect 244464 9104 244516 9110
rect 244464 9046 244516 9052
rect 245568 7812 245620 7818
rect 245568 7754 245620 7760
rect 244384 5222 244504 5250
rect 244372 5092 244424 5098
rect 244372 5034 244424 5040
rect 244280 3868 244332 3874
rect 244280 3810 244332 3816
rect 244384 480 244412 5034
rect 244476 3806 244504 5222
rect 244464 3800 244516 3806
rect 244464 3742 244516 3748
rect 245580 480 245608 7754
rect 246316 3942 246344 337214
rect 247132 335640 247184 335646
rect 247132 335582 247184 335588
rect 246764 9104 246816 9110
rect 246764 9046 246816 9052
rect 246304 3936 246356 3942
rect 246304 3878 246356 3884
rect 246776 480 246804 9046
rect 247144 5166 247172 335582
rect 247132 5160 247184 5166
rect 247132 5102 247184 5108
rect 247236 4010 247264 340054
rect 247696 335646 247724 340054
rect 247776 337272 247828 337278
rect 247776 337214 247828 337220
rect 247684 335640 247736 335646
rect 247684 335582 247736 335588
rect 247788 335458 247816 337214
rect 247696 335430 247816 335458
rect 247696 4078 247724 335430
rect 248524 10334 248552 340054
rect 248800 337278 248828 340068
rect 248892 340054 249274 340082
rect 249352 340054 249734 340082
rect 248788 337272 248840 337278
rect 248788 337214 248840 337220
rect 248604 332444 248656 332450
rect 248604 332386 248656 332392
rect 248616 10402 248644 332386
rect 248892 325718 248920 340054
rect 249064 337272 249116 337278
rect 249064 337214 249116 337220
rect 248880 325712 248932 325718
rect 248880 325654 248932 325660
rect 248788 322244 248840 322250
rect 248788 322186 248840 322192
rect 248800 317506 248828 322186
rect 248800 317478 248920 317506
rect 248892 311982 248920 317478
rect 248880 311976 248932 311982
rect 248880 311918 248932 311924
rect 248788 299532 248840 299538
rect 248788 299474 248840 299480
rect 248800 297378 248828 299474
rect 248708 297350 248828 297378
rect 248708 287722 248736 297350
rect 248708 287694 248828 287722
rect 248800 277794 248828 287694
rect 248708 277766 248828 277794
rect 248708 270586 248736 277766
rect 248708 270558 248828 270586
rect 248800 258482 248828 270558
rect 248708 258454 248828 258482
rect 248708 251274 248736 258454
rect 248708 251246 248828 251274
rect 248800 239442 248828 251246
rect 248708 239414 248828 239442
rect 248708 229786 248736 239414
rect 248708 229758 248828 229786
rect 248800 217954 248828 229758
rect 248708 217926 248828 217954
rect 248708 210746 248736 217926
rect 248708 210718 248828 210746
rect 248800 198642 248828 210718
rect 248708 198614 248828 198642
rect 248708 191434 248736 198614
rect 248708 191406 248828 191434
rect 248800 176798 248828 191406
rect 248788 176792 248840 176798
rect 248788 176734 248840 176740
rect 248696 176656 248748 176662
rect 248696 176598 248748 176604
rect 248708 171850 248736 176598
rect 248708 171822 248828 171850
rect 248800 162194 248828 171822
rect 248708 162166 248828 162194
rect 248708 152538 248736 162166
rect 248708 152510 248828 152538
rect 248800 123570 248828 152510
rect 248708 123542 248828 123570
rect 248708 113914 248736 123542
rect 248708 113886 248828 113914
rect 248800 104258 248828 113886
rect 248708 104230 248828 104258
rect 248708 94654 248736 104230
rect 248696 94648 248748 94654
rect 248696 94590 248748 94596
rect 248788 85604 248840 85610
rect 248788 85546 248840 85552
rect 248800 75886 248828 85546
rect 248788 75880 248840 75886
rect 248788 75822 248840 75828
rect 248788 66292 248840 66298
rect 248788 66234 248840 66240
rect 248800 62778 248828 66234
rect 248708 62750 248828 62778
rect 248708 55842 248736 62750
rect 248708 55814 248828 55842
rect 248800 19446 248828 55814
rect 248788 19440 248840 19446
rect 248788 19382 248840 19388
rect 248696 19372 248748 19378
rect 248696 19314 248748 19320
rect 248604 10396 248656 10402
rect 248604 10338 248656 10344
rect 248512 10328 248564 10334
rect 248512 10270 248564 10276
rect 248708 5234 248736 19314
rect 248696 5228 248748 5234
rect 248696 5170 248748 5176
rect 247960 5160 248012 5166
rect 247960 5102 248012 5108
rect 247684 4072 247736 4078
rect 247684 4014 247736 4020
rect 247224 4004 247276 4010
rect 247224 3946 247276 3952
rect 247972 480 248000 5102
rect 249076 4146 249104 337214
rect 249352 332450 249380 340054
rect 250180 338026 250208 340068
rect 250272 340054 250654 340082
rect 250824 340054 251114 340082
rect 250168 338020 250220 338026
rect 250168 337962 250220 337968
rect 249892 335640 249944 335646
rect 250272 335594 250300 340054
rect 250444 337884 250496 337890
rect 250444 337826 250496 337832
rect 249892 335582 249944 335588
rect 249340 332444 249392 332450
rect 249340 332386 249392 332392
rect 249248 325712 249300 325718
rect 249248 325654 249300 325660
rect 249260 322250 249288 325654
rect 249248 322244 249300 322250
rect 249248 322186 249300 322192
rect 249706 29336 249762 29345
rect 249706 29271 249762 29280
rect 249720 28937 249748 29271
rect 249706 28928 249762 28937
rect 249706 28863 249762 28872
rect 249904 10470 249932 335582
rect 250180 335566 250300 335594
rect 250180 335345 250208 335566
rect 250166 335336 250222 335345
rect 250166 335271 250222 335280
rect 250258 335200 250314 335209
rect 250258 335135 250314 335144
rect 250272 325689 250300 335135
rect 249982 325680 250038 325689
rect 249982 325615 250038 325624
rect 250258 325680 250314 325689
rect 250258 325615 250314 325624
rect 249996 316130 250024 325615
rect 249984 316124 250036 316130
rect 249984 316066 250036 316072
rect 250168 316124 250220 316130
rect 250168 316066 250220 316072
rect 250180 315994 250208 316066
rect 250168 315988 250220 315994
rect 250168 315930 250220 315936
rect 250076 299532 250128 299538
rect 250076 299474 250128 299480
rect 250088 297378 250116 299474
rect 249996 297350 250116 297378
rect 249996 287722 250024 297350
rect 249996 287694 250116 287722
rect 250088 277794 250116 287694
rect 249996 277766 250116 277794
rect 249996 270586 250024 277766
rect 249996 270558 250116 270586
rect 250088 258482 250116 270558
rect 249996 258454 250116 258482
rect 249996 251274 250024 258454
rect 249996 251246 250116 251274
rect 250088 239442 250116 251246
rect 249996 239414 250116 239442
rect 249996 229786 250024 239414
rect 249996 229758 250116 229786
rect 250088 217954 250116 229758
rect 249996 217926 250116 217954
rect 249996 210746 250024 217926
rect 249996 210718 250116 210746
rect 250088 198642 250116 210718
rect 249996 198614 250116 198642
rect 249996 191434 250024 198614
rect 249996 191406 250116 191434
rect 250088 178786 250116 191406
rect 249996 178758 250116 178786
rect 249996 171850 250024 178758
rect 249996 171822 250116 171850
rect 250088 162194 250116 171822
rect 249996 162166 250116 162194
rect 249996 152538 250024 162166
rect 249996 152510 250116 152538
rect 250088 123570 250116 152510
rect 249996 123542 250116 123570
rect 249996 113914 250024 123542
rect 249996 113886 250116 113914
rect 250088 104258 250116 113886
rect 249996 104230 250116 104258
rect 249996 94602 250024 104230
rect 249996 94574 250116 94602
rect 250088 56642 250116 94574
rect 249984 56636 250036 56642
rect 249984 56578 250036 56584
rect 250076 56636 250128 56642
rect 250076 56578 250128 56584
rect 249996 55842 250024 56578
rect 249996 55814 250116 55842
rect 250088 19378 250116 55814
rect 249984 19372 250036 19378
rect 249984 19314 250036 19320
rect 250076 19372 250128 19378
rect 250076 19314 250128 19320
rect 249892 10464 249944 10470
rect 249892 10406 249944 10412
rect 249156 7880 249208 7886
rect 249156 7822 249208 7828
rect 249064 4140 249116 4146
rect 249064 4082 249116 4088
rect 249168 480 249196 7822
rect 249996 6225 250024 19314
rect 250352 9172 250404 9178
rect 250352 9114 250404 9120
rect 249982 6216 250038 6225
rect 249982 6151 250038 6160
rect 250364 480 250392 9114
rect 250456 3398 250484 337826
rect 250824 335646 250852 340054
rect 251560 337278 251588 340068
rect 251652 340054 252034 340082
rect 252112 340054 252402 340082
rect 251548 337272 251600 337278
rect 251548 337214 251600 337220
rect 250812 335640 250864 335646
rect 250812 335582 250864 335588
rect 251272 335640 251324 335646
rect 251652 335594 251680 340054
rect 251824 337952 251876 337958
rect 251824 337894 251876 337900
rect 251272 335582 251324 335588
rect 251178 288416 251234 288425
rect 251178 288351 251234 288360
rect 251192 278798 251220 288351
rect 251180 278792 251232 278798
rect 251180 278734 251232 278740
rect 251180 224256 251232 224262
rect 251180 224198 251232 224204
rect 251192 219473 251220 224198
rect 251178 219464 251234 219473
rect 251178 219399 251234 219408
rect 251180 151836 251232 151842
rect 251180 151778 251232 151784
rect 251192 143585 251220 151778
rect 251178 143576 251234 143585
rect 251178 143511 251234 143520
rect 251180 133952 251232 133958
rect 251178 133920 251180 133929
rect 251232 133920 251234 133929
rect 251178 133855 251234 133864
rect 251180 95192 251232 95198
rect 251180 95134 251232 95140
rect 251192 85649 251220 95134
rect 251178 85640 251234 85649
rect 251178 85575 251234 85584
rect 251284 10538 251312 335582
rect 251468 335566 251680 335594
rect 251468 328438 251496 335566
rect 251456 328432 251508 328438
rect 251456 328374 251508 328380
rect 251640 328432 251692 328438
rect 251640 328374 251692 328380
rect 251652 318918 251680 328374
rect 251640 318912 251692 318918
rect 251640 318854 251692 318860
rect 251456 318776 251508 318782
rect 251456 318718 251508 318724
rect 251362 288416 251418 288425
rect 251468 288402 251496 318718
rect 251418 288374 251496 288402
rect 251362 288351 251418 288360
rect 251456 278792 251508 278798
rect 251456 278734 251508 278740
rect 251468 273902 251496 278734
rect 251456 273896 251508 273902
rect 251456 273838 251508 273844
rect 251456 260908 251508 260914
rect 251456 260850 251508 260856
rect 251468 259418 251496 260850
rect 251456 259412 251508 259418
rect 251456 259354 251508 259360
rect 251548 251116 251600 251122
rect 251548 251058 251600 251064
rect 251560 249778 251588 251058
rect 251468 249750 251588 249778
rect 251468 241534 251496 249750
rect 251456 241528 251508 241534
rect 251456 241470 251508 241476
rect 251456 240168 251508 240174
rect 251456 240110 251508 240116
rect 251468 240038 251496 240110
rect 251456 240032 251508 240038
rect 251456 239974 251508 239980
rect 251456 230512 251508 230518
rect 251456 230454 251508 230460
rect 251468 224262 251496 230454
rect 251456 224256 251508 224262
rect 251456 224198 251508 224204
rect 251362 219464 251418 219473
rect 251362 219399 251418 219408
rect 251376 209778 251404 219399
rect 251364 209772 251416 209778
rect 251364 209714 251416 209720
rect 251732 209772 251784 209778
rect 251732 209714 251784 209720
rect 251744 200161 251772 209714
rect 251546 200152 251602 200161
rect 251546 200087 251602 200096
rect 251730 200152 251786 200161
rect 251730 200087 251786 200096
rect 251560 191894 251588 200087
rect 251456 191888 251508 191894
rect 251456 191830 251508 191836
rect 251548 191888 251600 191894
rect 251548 191830 251600 191836
rect 251468 182345 251496 191830
rect 251454 182336 251510 182345
rect 251454 182271 251510 182280
rect 251638 182064 251694 182073
rect 251638 181999 251694 182008
rect 251652 172553 251680 181999
rect 251454 172544 251510 172553
rect 251364 172508 251416 172514
rect 251454 172479 251456 172488
rect 251364 172450 251416 172456
rect 251508 172479 251510 172488
rect 251638 172544 251694 172553
rect 251638 172479 251694 172488
rect 251456 172450 251508 172456
rect 251376 171086 251404 172450
rect 251364 171080 251416 171086
rect 251364 171022 251416 171028
rect 251456 161492 251508 161498
rect 251456 161434 251508 161440
rect 251468 161378 251496 161434
rect 251376 161350 251496 161378
rect 251376 151842 251404 161350
rect 251364 151836 251416 151842
rect 251364 151778 251416 151784
rect 251362 143576 251418 143585
rect 251362 143511 251364 143520
rect 251416 143511 251418 143520
rect 251364 143482 251416 143488
rect 251548 135244 251600 135250
rect 251548 135186 251600 135192
rect 251560 133890 251588 135186
rect 251548 133884 251600 133890
rect 251548 133826 251600 133832
rect 251456 124228 251508 124234
rect 251456 124170 251508 124176
rect 251468 114458 251496 124170
rect 251376 114430 251496 114458
rect 251376 105097 251404 114430
rect 251362 105088 251418 105097
rect 251362 105023 251418 105032
rect 251454 104952 251510 104961
rect 251454 104887 251510 104896
rect 251468 104854 251496 104887
rect 251456 104848 251508 104854
rect 251456 104790 251508 104796
rect 251456 95328 251508 95334
rect 251456 95270 251508 95276
rect 251468 95198 251496 95270
rect 251456 95192 251508 95198
rect 251456 95134 251508 95140
rect 251362 85640 251418 85649
rect 251362 85575 251418 85584
rect 251376 79370 251404 85575
rect 251376 79342 251496 79370
rect 251468 56817 251496 79342
rect 251454 56808 251510 56817
rect 251454 56743 251510 56752
rect 251454 56536 251510 56545
rect 251454 56471 251510 56480
rect 251468 46918 251496 56471
rect 251364 46912 251416 46918
rect 251364 46854 251416 46860
rect 251456 46912 251508 46918
rect 251456 46854 251508 46860
rect 251376 37346 251404 46854
rect 251376 37318 251496 37346
rect 251468 27606 251496 37318
rect 251456 27600 251508 27606
rect 251456 27542 251508 27548
rect 251548 17944 251600 17950
rect 251548 17886 251600 17892
rect 251272 10532 251324 10538
rect 251272 10474 251324 10480
rect 251560 8401 251588 17886
rect 251362 8392 251418 8401
rect 251362 8327 251418 8336
rect 251546 8392 251602 8401
rect 251546 8327 251602 8336
rect 251376 8242 251404 8327
rect 251284 8214 251404 8242
rect 251284 6186 251312 8214
rect 251272 6180 251324 6186
rect 251272 6122 251324 6128
rect 251456 5228 251508 5234
rect 251456 5170 251508 5176
rect 250444 3392 250496 3398
rect 250444 3334 250496 3340
rect 251468 480 251496 5170
rect 251836 3330 251864 337894
rect 252112 335646 252140 340054
rect 252848 337414 252876 340068
rect 252940 340054 253322 340082
rect 253400 340054 253782 340082
rect 252836 337408 252888 337414
rect 252836 337350 252888 337356
rect 252100 335640 252152 335646
rect 252100 335582 252152 335588
rect 252652 335640 252704 335646
rect 252652 335582 252704 335588
rect 252664 10606 252692 335582
rect 252940 311794 252968 340054
rect 253204 337272 253256 337278
rect 253204 337214 253256 337220
rect 252848 311766 252968 311794
rect 252848 297378 252876 311766
rect 252756 297350 252876 297378
rect 252756 287722 252784 297350
rect 252756 287694 252876 287722
rect 252848 277794 252876 287694
rect 252756 277766 252876 277794
rect 252756 270586 252784 277766
rect 252756 270558 252876 270586
rect 252848 258482 252876 270558
rect 252756 258454 252876 258482
rect 252756 251274 252784 258454
rect 252756 251246 252876 251274
rect 252848 239442 252876 251246
rect 252756 239414 252876 239442
rect 252756 229786 252784 239414
rect 252756 229758 252876 229786
rect 252848 217954 252876 229758
rect 252756 217926 252876 217954
rect 252756 210746 252784 217926
rect 252756 210718 252876 210746
rect 252848 198642 252876 210718
rect 252756 198614 252876 198642
rect 252756 191434 252784 198614
rect 252756 191406 252876 191434
rect 252848 172530 252876 191406
rect 252756 172502 252876 172530
rect 252756 171850 252784 172502
rect 252756 171822 252876 171850
rect 252848 162194 252876 171822
rect 252756 162166 252876 162194
rect 252756 152538 252784 162166
rect 252756 152510 252876 152538
rect 252848 123622 252876 152510
rect 252836 123616 252888 123622
rect 252836 123558 252888 123564
rect 252744 123548 252796 123554
rect 252744 123490 252796 123496
rect 252756 113914 252784 123490
rect 252756 113886 252876 113914
rect 252848 104258 252876 113886
rect 252756 104230 252876 104258
rect 252756 94602 252784 104230
rect 252756 94574 252876 94602
rect 252848 67590 252876 94574
rect 252744 67584 252796 67590
rect 252744 67526 252796 67532
rect 252836 67584 252888 67590
rect 252836 67526 252888 67532
rect 252756 53174 252784 67526
rect 252744 53168 252796 53174
rect 252744 53110 252796 53116
rect 252836 53100 252888 53106
rect 252836 53042 252888 53048
rect 252848 22778 252876 53042
rect 252836 22772 252888 22778
rect 252836 22714 252888 22720
rect 252652 10600 252704 10606
rect 252652 10542 252704 10548
rect 252744 9716 252796 9722
rect 252744 9658 252796 9664
rect 252652 7948 252704 7954
rect 252652 7890 252704 7896
rect 251824 3324 251876 3330
rect 251824 3266 251876 3272
rect 252664 480 252692 7890
rect 252756 6254 252784 9658
rect 252744 6248 252796 6254
rect 252744 6190 252796 6196
rect 253216 3262 253244 337214
rect 253400 335646 253428 340054
rect 254228 337890 254256 340068
rect 254320 340054 254702 340082
rect 254780 340054 255162 340082
rect 254216 337884 254268 337890
rect 254216 337826 254268 337832
rect 253388 335640 253440 335646
rect 254320 335628 254348 340054
rect 254780 338042 254808 340054
rect 253388 335582 253440 335588
rect 254044 335600 254348 335628
rect 254412 338014 254808 338042
rect 253938 306368 253994 306377
rect 253938 306303 253994 306312
rect 253952 296750 253980 306303
rect 253940 296744 253992 296750
rect 253940 296686 253992 296692
rect 253754 87136 253810 87145
rect 253938 87136 253994 87145
rect 253810 87094 253938 87122
rect 253754 87071 253810 87080
rect 253938 87071 253994 87080
rect 253940 32428 253992 32434
rect 253940 32370 253992 32376
rect 253952 22778 253980 32370
rect 253940 22772 253992 22778
rect 253940 22714 253992 22720
rect 254044 6322 254072 335600
rect 254412 335458 254440 338014
rect 254584 337816 254636 337822
rect 254584 337758 254636 337764
rect 254228 335430 254440 335458
rect 254228 328438 254256 335430
rect 254216 328432 254268 328438
rect 254216 328374 254268 328380
rect 254308 328432 254360 328438
rect 254308 328374 254360 328380
rect 254320 322266 254348 328374
rect 254136 322238 254348 322266
rect 254136 316010 254164 322238
rect 254136 315982 254348 316010
rect 254320 306474 254348 315982
rect 254124 306468 254176 306474
rect 254124 306410 254176 306416
rect 254308 306468 254360 306474
rect 254308 306410 254360 306416
rect 254136 306377 254164 306410
rect 254122 306368 254178 306377
rect 254122 306303 254178 306312
rect 254216 296744 254268 296750
rect 254216 296686 254268 296692
rect 254228 292670 254256 296686
rect 254216 292664 254268 292670
rect 254216 292606 254268 292612
rect 254216 292528 254268 292534
rect 254216 292470 254268 292476
rect 254228 280158 254256 292470
rect 254216 280152 254268 280158
rect 254216 280094 254268 280100
rect 254216 270564 254268 270570
rect 254216 270506 254268 270512
rect 254228 260846 254256 270506
rect 254216 260840 254268 260846
rect 254216 260782 254268 260788
rect 254216 251252 254268 251258
rect 254216 251194 254268 251200
rect 254228 241505 254256 251194
rect 254214 241496 254270 241505
rect 254214 241431 254270 241440
rect 254398 241496 254454 241505
rect 254398 241431 254454 241440
rect 254412 231878 254440 241431
rect 254216 231872 254268 231878
rect 254216 231814 254268 231820
rect 254400 231872 254452 231878
rect 254400 231814 254452 231820
rect 254228 222193 254256 231814
rect 254214 222184 254270 222193
rect 254214 222119 254270 222128
rect 254398 222184 254454 222193
rect 254398 222119 254454 222128
rect 254412 212566 254440 222119
rect 254216 212560 254268 212566
rect 254216 212502 254268 212508
rect 254400 212560 254452 212566
rect 254400 212502 254452 212508
rect 254228 196654 254256 212502
rect 254216 196648 254268 196654
rect 254216 196590 254268 196596
rect 254400 196648 254452 196654
rect 254400 196590 254452 196596
rect 254412 191865 254440 196590
rect 254214 191856 254270 191865
rect 254214 191791 254270 191800
rect 254398 191856 254454 191865
rect 254398 191791 254454 191800
rect 254228 164218 254256 191791
rect 254216 164212 254268 164218
rect 254216 164154 254268 164160
rect 254400 164212 254452 164218
rect 254400 164154 254452 164160
rect 254412 154601 254440 164154
rect 254214 154592 254270 154601
rect 254214 154527 254270 154536
rect 254398 154592 254454 154601
rect 254398 154527 254454 154536
rect 254228 144906 254256 154527
rect 254216 144900 254268 144906
rect 254216 144842 254268 144848
rect 254400 144900 254452 144906
rect 254400 144842 254452 144848
rect 254412 135289 254440 144842
rect 254214 135280 254270 135289
rect 254214 135215 254270 135224
rect 254398 135280 254454 135289
rect 254398 135215 254454 135224
rect 254228 125594 254256 135215
rect 254216 125588 254268 125594
rect 254216 125530 254268 125536
rect 254216 116000 254268 116006
rect 254216 115942 254268 115948
rect 254228 99498 254256 115942
rect 254136 99470 254256 99498
rect 254136 99362 254164 99470
rect 254136 99334 254256 99362
rect 254228 80102 254256 99334
rect 254216 80096 254268 80102
rect 254216 80038 254268 80044
rect 254216 79960 254268 79966
rect 254216 79902 254268 79908
rect 254228 56658 254256 79902
rect 254136 56630 254256 56658
rect 254136 56574 254164 56630
rect 254124 56568 254176 56574
rect 254124 56510 254176 56516
rect 254124 46980 254176 46986
rect 254124 46922 254176 46928
rect 254136 37330 254164 46922
rect 254124 37324 254176 37330
rect 254124 37266 254176 37272
rect 254216 37324 254268 37330
rect 254216 37266 254268 37272
rect 254228 32434 254256 37266
rect 254216 32428 254268 32434
rect 254216 32370 254268 32376
rect 254124 9716 254176 9722
rect 254124 9658 254176 9664
rect 254032 6316 254084 6322
rect 254032 6258 254084 6264
rect 253848 6180 253900 6186
rect 253848 6122 253900 6128
rect 253204 3256 253256 3262
rect 253204 3198 253256 3204
rect 253860 480 253888 6122
rect 254136 5302 254164 9658
rect 254124 5296 254176 5302
rect 254124 5238 254176 5244
rect 254596 3194 254624 337758
rect 254860 337680 254912 337686
rect 254860 337622 254912 337628
rect 254872 334506 254900 337622
rect 255608 336870 255636 340068
rect 255884 340054 256082 340082
rect 256160 340054 256450 340082
rect 255596 336864 255648 336870
rect 255596 336806 255648 336812
rect 255412 335640 255464 335646
rect 255412 335582 255464 335588
rect 254688 334478 254900 334506
rect 254584 3188 254636 3194
rect 254584 3130 254636 3136
rect 254688 3126 254716 334478
rect 255320 153196 255372 153202
rect 255320 153138 255372 153144
rect 255332 143585 255360 153138
rect 255318 143576 255374 143585
rect 255318 143511 255374 143520
rect 255320 22772 255372 22778
rect 255320 22714 255372 22720
rect 255332 12322 255360 22714
rect 255424 13190 255452 335582
rect 255884 331242 255912 340054
rect 255964 337340 256016 337346
rect 255964 337282 256016 337288
rect 255608 331214 255912 331242
rect 255608 331106 255636 331214
rect 255608 331078 255728 331106
rect 255700 321638 255728 331078
rect 255688 321632 255740 321638
rect 255688 321574 255740 321580
rect 255688 321428 255740 321434
rect 255688 321370 255740 321376
rect 255700 292618 255728 321370
rect 255608 292590 255728 292618
rect 255608 288402 255636 292590
rect 255516 288374 255636 288402
rect 255516 278798 255544 288374
rect 255504 278792 255556 278798
rect 255504 278734 255556 278740
rect 255872 278792 255924 278798
rect 255872 278734 255924 278740
rect 255884 270570 255912 278734
rect 255596 270564 255648 270570
rect 255596 270506 255648 270512
rect 255872 270564 255924 270570
rect 255872 270506 255924 270512
rect 255608 270434 255636 270506
rect 255596 270428 255648 270434
rect 255596 270370 255648 270376
rect 255688 260908 255740 260914
rect 255688 260850 255740 260856
rect 255700 260778 255728 260850
rect 255688 260772 255740 260778
rect 255688 260714 255740 260720
rect 255596 251252 255648 251258
rect 255596 251194 255648 251200
rect 255608 251161 255636 251194
rect 255594 251152 255650 251161
rect 255594 251087 255650 251096
rect 255778 251152 255834 251161
rect 255778 251087 255834 251096
rect 255792 241534 255820 251087
rect 255780 241528 255832 241534
rect 255780 241470 255832 241476
rect 255872 241528 255924 241534
rect 255872 241470 255924 241476
rect 255884 230518 255912 241470
rect 255780 230512 255832 230518
rect 255780 230454 255832 230460
rect 255872 230512 255924 230518
rect 255872 230454 255924 230460
rect 255792 220810 255820 230454
rect 255608 220782 255820 220810
rect 255608 202978 255636 220782
rect 255596 202972 255648 202978
rect 255596 202914 255648 202920
rect 255688 202972 255740 202978
rect 255688 202914 255740 202920
rect 255700 192001 255728 202914
rect 255686 191992 255742 192001
rect 255686 191927 255742 191936
rect 255594 191856 255650 191865
rect 255594 191791 255596 191800
rect 255648 191791 255650 191800
rect 255596 191762 255648 191768
rect 255596 186312 255648 186318
rect 255596 186254 255648 186260
rect 255608 182186 255636 186254
rect 255608 182170 255728 182186
rect 255608 182164 255740 182170
rect 255608 182158 255688 182164
rect 255688 182106 255740 182112
rect 255596 172576 255648 172582
rect 255596 172518 255648 172524
rect 255608 164286 255636 172518
rect 255596 164280 255648 164286
rect 255596 164222 255648 164228
rect 255688 164144 255740 164150
rect 255688 164086 255740 164092
rect 255700 154698 255728 164086
rect 255596 154692 255648 154698
rect 255596 154634 255648 154640
rect 255688 154692 255740 154698
rect 255688 154634 255740 154640
rect 255608 153202 255636 154634
rect 255596 153196 255648 153202
rect 255596 153138 255648 153144
rect 255502 143576 255558 143585
rect 255502 143511 255558 143520
rect 255516 130490 255544 143511
rect 255504 130484 255556 130490
rect 255504 130426 255556 130432
rect 255780 130484 255832 130490
rect 255780 130426 255832 130432
rect 255792 116090 255820 130426
rect 255700 116062 255820 116090
rect 255700 115954 255728 116062
rect 255608 115926 255728 115954
rect 255608 114510 255636 115926
rect 255596 114504 255648 114510
rect 255596 114446 255648 114452
rect 255596 104916 255648 104922
rect 255596 104858 255648 104864
rect 255608 98734 255636 104858
rect 255596 98728 255648 98734
rect 255596 98670 255648 98676
rect 255688 93900 255740 93906
rect 255688 93842 255740 93848
rect 255700 93770 255728 93842
rect 255688 93764 255740 93770
rect 255688 93706 255740 93712
rect 255780 84244 255832 84250
rect 255780 84186 255832 84192
rect 255792 77586 255820 84186
rect 255596 77580 255648 77586
rect 255596 77522 255648 77528
rect 255780 77580 255832 77586
rect 255780 77522 255832 77528
rect 255608 66230 255636 77522
rect 255596 66224 255648 66230
rect 255596 66166 255648 66172
rect 255780 64728 255832 64734
rect 255780 64670 255832 64676
rect 255792 55214 255820 64670
rect 255780 55208 255832 55214
rect 255780 55150 255832 55156
rect 255596 45688 255648 45694
rect 255596 45630 255648 45636
rect 255608 45558 255636 45630
rect 255596 45552 255648 45558
rect 255596 45494 255648 45500
rect 255688 45552 255740 45558
rect 255688 45494 255740 45500
rect 255700 22778 255728 45494
rect 255688 22772 255740 22778
rect 255688 22714 255740 22720
rect 255412 13184 255464 13190
rect 255412 13126 255464 13132
rect 255332 12294 255452 12322
rect 255424 6390 255452 12294
rect 255412 6384 255464 6390
rect 255412 6326 255464 6332
rect 255044 3460 255096 3466
rect 255044 3402 255096 3408
rect 254676 3120 254728 3126
rect 254676 3062 254728 3068
rect 255056 480 255084 3402
rect 255976 3058 256004 337282
rect 256160 335646 256188 340054
rect 256896 337958 256924 340068
rect 256988 340054 257370 340082
rect 257448 340054 257830 340082
rect 256884 337952 256936 337958
rect 256884 337894 256936 337900
rect 256148 335640 256200 335646
rect 256148 335582 256200 335588
rect 256792 334076 256844 334082
rect 256792 334018 256844 334024
rect 256804 14550 256832 334018
rect 256792 14544 256844 14550
rect 256792 14486 256844 14492
rect 256240 8016 256292 8022
rect 256240 7958 256292 7964
rect 255964 3052 256016 3058
rect 255964 2994 256016 3000
rect 256252 480 256280 7958
rect 256988 6458 257016 340054
rect 257344 337476 257396 337482
rect 257344 337418 257396 337424
rect 256976 6452 257028 6458
rect 256976 6394 257028 6400
rect 257356 2990 257384 337418
rect 257448 334082 257476 340054
rect 258276 338094 258304 340068
rect 258368 340054 258750 340082
rect 258920 340054 259210 340082
rect 258264 338088 258316 338094
rect 258264 338030 258316 338036
rect 258172 335640 258224 335646
rect 258172 335582 258224 335588
rect 257436 334076 257488 334082
rect 257436 334018 257488 334024
rect 258184 14618 258212 335582
rect 258172 14612 258224 14618
rect 258172 14554 258224 14560
rect 258368 6526 258396 340054
rect 258816 337612 258868 337618
rect 258816 337554 258868 337560
rect 258724 337544 258776 337550
rect 258724 337486 258776 337492
rect 258356 6520 258408 6526
rect 258356 6462 258408 6468
rect 257436 6248 257488 6254
rect 257436 6190 257488 6196
rect 257344 2984 257396 2990
rect 257344 2926 257396 2932
rect 257448 480 257476 6190
rect 258632 3596 258684 3602
rect 258632 3538 258684 3544
rect 258644 480 258672 3538
rect 258736 2922 258764 337486
rect 258724 2916 258776 2922
rect 258724 2858 258776 2864
rect 258828 2854 258856 337554
rect 258920 335646 258948 340054
rect 259552 337952 259604 337958
rect 259552 337894 259604 337900
rect 259460 337680 259512 337686
rect 259564 337668 259592 337894
rect 259512 337640 259592 337668
rect 259460 337622 259512 337628
rect 259656 337278 259684 340068
rect 259748 340054 260038 340082
rect 260208 340054 260498 340082
rect 259644 337272 259696 337278
rect 259644 337214 259696 337220
rect 258908 335640 258960 335646
rect 258908 335582 258960 335588
rect 259552 335640 259604 335646
rect 259552 335582 259604 335588
rect 259564 14686 259592 335582
rect 259552 14680 259604 14686
rect 259552 14622 259604 14628
rect 259748 8090 259776 340054
rect 260208 335646 260236 340054
rect 260944 337822 260972 340068
rect 261036 340054 261418 340082
rect 261588 340054 261878 340082
rect 260932 337816 260984 337822
rect 260932 337758 260984 337764
rect 260196 335640 260248 335646
rect 260196 335582 260248 335588
rect 260746 134192 260802 134201
rect 260746 134127 260802 134136
rect 260760 133958 260788 134127
rect 260748 133952 260800 133958
rect 260748 133894 260800 133900
rect 261036 8158 261064 340054
rect 261588 331242 261616 340054
rect 262324 337006 262352 340068
rect 262416 340054 262798 340082
rect 263060 340054 263258 340082
rect 262312 337000 262364 337006
rect 262312 336942 262364 336948
rect 261220 331214 261616 331242
rect 261220 321638 261248 331214
rect 261208 321632 261260 321638
rect 261208 321574 261260 321580
rect 261300 321428 261352 321434
rect 261300 321370 261352 321376
rect 261312 289882 261340 321370
rect 261208 289876 261260 289882
rect 261208 289818 261260 289824
rect 261300 289876 261352 289882
rect 261300 289818 261352 289824
rect 261220 273222 261248 289818
rect 262416 278934 262444 340054
rect 263060 328506 263088 340054
rect 263612 338026 263640 340068
rect 263796 340054 264086 340082
rect 264256 340054 264546 340082
rect 263600 338020 263652 338026
rect 263600 337962 263652 337968
rect 263692 335640 263744 335646
rect 263692 335582 263744 335588
rect 262680 328500 262732 328506
rect 262680 328442 262732 328448
rect 263048 328500 263100 328506
rect 263048 328442 263100 328448
rect 262692 318782 262720 328442
rect 262680 318776 262732 318782
rect 262680 318718 262732 318724
rect 262680 312180 262732 312186
rect 262680 312122 262732 312128
rect 262692 299470 262720 312122
rect 262680 299464 262732 299470
rect 262680 299406 262732 299412
rect 262588 289944 262640 289950
rect 262588 289886 262640 289892
rect 262600 288386 262628 289886
rect 262588 288380 262640 288386
rect 262588 288322 262640 288328
rect 262404 278928 262456 278934
rect 262404 278870 262456 278876
rect 262496 278860 262548 278866
rect 262496 278802 262548 278808
rect 262404 278792 262456 278798
rect 262404 278734 262456 278740
rect 261208 273216 261260 273222
rect 261208 273158 261260 273164
rect 261208 273080 261260 273086
rect 261208 273022 261260 273028
rect 261220 253910 261248 273022
rect 261208 253904 261260 253910
rect 261208 253846 261260 253852
rect 261208 253768 261260 253774
rect 261208 253710 261260 253716
rect 261220 234598 261248 253710
rect 261208 234592 261260 234598
rect 261208 234534 261260 234540
rect 261208 234456 261260 234462
rect 261208 234398 261260 234404
rect 261220 216034 261248 234398
rect 261208 216028 261260 216034
rect 261208 215970 261260 215976
rect 261392 216028 261444 216034
rect 261392 215970 261444 215976
rect 261404 211177 261432 215970
rect 261206 211168 261262 211177
rect 261206 211103 261262 211112
rect 261390 211168 261446 211177
rect 261390 211103 261446 211112
rect 261220 186454 261248 211103
rect 261208 186448 261260 186454
rect 261208 186390 261260 186396
rect 261208 186312 261260 186318
rect 261208 186254 261260 186260
rect 261220 173942 261248 186254
rect 261208 173936 261260 173942
rect 261208 173878 261260 173884
rect 261300 173936 261352 173942
rect 261300 173878 261352 173884
rect 261312 171034 261340 173878
rect 261312 171006 261432 171034
rect 261404 162858 261432 171006
rect 261392 162852 261444 162858
rect 261392 162794 261444 162800
rect 261300 153264 261352 153270
rect 261300 153206 261352 153212
rect 261312 133906 261340 153206
rect 261312 133878 261432 133906
rect 261404 125769 261432 133878
rect 261390 125760 261446 125769
rect 261390 125695 261446 125704
rect 261298 125624 261354 125633
rect 261298 125559 261354 125568
rect 261312 124166 261340 125559
rect 261300 124160 261352 124166
rect 261300 124102 261352 124108
rect 261208 118652 261260 118658
rect 261208 118594 261260 118600
rect 261220 99498 261248 118594
rect 261128 99470 261248 99498
rect 261128 99362 261156 99470
rect 261128 99334 261248 99362
rect 261220 82226 261248 99334
rect 261128 82198 261248 82226
rect 261128 77246 261156 82198
rect 261116 77240 261168 77246
rect 261116 77182 261168 77188
rect 261300 77172 261352 77178
rect 261300 77114 261352 77120
rect 261312 60858 261340 77114
rect 261300 60852 261352 60858
rect 261300 60794 261352 60800
rect 261208 60716 261260 60722
rect 261208 60658 261260 60664
rect 261220 53174 261248 60658
rect 261208 53168 261260 53174
rect 261208 53110 261260 53116
rect 261300 48340 261352 48346
rect 261300 48282 261352 48288
rect 261312 37346 261340 48282
rect 261220 37318 261340 37346
rect 261220 31822 261248 37318
rect 261208 31816 261260 31822
rect 261208 31758 261260 31764
rect 261208 27668 261260 27674
rect 261208 27610 261260 27616
rect 261220 19378 261248 27610
rect 261116 19372 261168 19378
rect 261116 19314 261168 19320
rect 261208 19372 261260 19378
rect 261208 19314 261260 19320
rect 261128 14754 261156 19314
rect 261116 14748 261168 14754
rect 261116 14690 261168 14696
rect 262416 8226 262444 278734
rect 262508 278730 262536 278802
rect 262496 278724 262548 278730
rect 262496 278666 262548 278672
rect 262680 263492 262732 263498
rect 262680 263434 262732 263440
rect 262692 260846 262720 263434
rect 262680 260840 262732 260846
rect 262680 260782 262732 260788
rect 262588 251252 262640 251258
rect 262588 251194 262640 251200
rect 262600 246378 262628 251194
rect 262600 246350 262812 246378
rect 262784 241534 262812 246350
rect 262772 241528 262824 241534
rect 262772 241470 262824 241476
rect 262864 241528 262916 241534
rect 262864 241470 262916 241476
rect 262876 231878 262904 241470
rect 262588 231872 262640 231878
rect 262588 231814 262640 231820
rect 262864 231872 262916 231878
rect 262864 231814 262916 231820
rect 262600 227066 262628 231814
rect 262508 227038 262628 227066
rect 262508 222222 262536 227038
rect 262496 222216 262548 222222
rect 262496 222158 262548 222164
rect 262864 222216 262916 222222
rect 262864 222158 262916 222164
rect 262876 212566 262904 222158
rect 262588 212560 262640 212566
rect 262588 212502 262640 212508
rect 262864 212560 262916 212566
rect 262864 212502 262916 212508
rect 262600 193390 262628 212502
rect 262588 193384 262640 193390
rect 262588 193326 262640 193332
rect 262588 193248 262640 193254
rect 262588 193190 262640 193196
rect 262600 191826 262628 193190
rect 262588 191820 262640 191826
rect 262588 191762 262640 191768
rect 262588 183524 262640 183530
rect 262588 183466 262640 183472
rect 262600 182186 262628 183466
rect 262600 182158 262720 182186
rect 262692 173942 262720 182158
rect 262680 173936 262732 173942
rect 262680 173878 262732 173884
rect 262772 173800 262824 173806
rect 262772 173742 262824 173748
rect 262784 164286 262812 173742
rect 262680 164280 262732 164286
rect 262680 164222 262732 164228
rect 262772 164280 262824 164286
rect 262772 164222 262824 164228
rect 262692 162858 262720 164222
rect 262680 162852 262732 162858
rect 262680 162794 262732 162800
rect 262496 153264 262548 153270
rect 262496 153206 262548 153212
rect 262508 144945 262536 153206
rect 262494 144936 262550 144945
rect 262494 144871 262550 144880
rect 262678 144936 262734 144945
rect 262678 144871 262734 144880
rect 262692 139398 262720 144871
rect 262680 139392 262732 139398
rect 262680 139334 262732 139340
rect 262864 129804 262916 129810
rect 262864 129746 262916 129752
rect 262876 120086 262904 129746
rect 262864 120080 262916 120086
rect 262864 120022 262916 120028
rect 262680 102196 262732 102202
rect 262680 102138 262732 102144
rect 262692 99482 262720 102138
rect 262680 99476 262732 99482
rect 262680 99418 262732 99424
rect 262496 86964 262548 86970
rect 262496 86906 262548 86912
rect 262508 77246 262536 86906
rect 262496 77240 262548 77246
rect 262496 77182 262548 77188
rect 262864 77240 262916 77246
rect 262864 77182 262916 77188
rect 262876 75886 262904 77182
rect 262864 75880 262916 75886
rect 262864 75822 262916 75828
rect 262772 66292 262824 66298
rect 262772 66234 262824 66240
rect 262784 66178 262812 66234
rect 262784 66150 262904 66178
rect 262876 56642 262904 66150
rect 262680 56636 262732 56642
rect 262680 56578 262732 56584
rect 262864 56636 262916 56642
rect 262864 56578 262916 56584
rect 262692 56506 262720 56578
rect 262680 56500 262732 56506
rect 262680 56442 262732 56448
rect 262864 56500 262916 56506
rect 262864 56442 262916 56448
rect 262876 46918 262904 56442
rect 262864 46912 262916 46918
rect 262864 46854 262916 46860
rect 262680 37324 262732 37330
rect 262680 37266 262732 37272
rect 262692 24206 262720 37266
rect 262680 24200 262732 24206
rect 262680 24142 262732 24148
rect 262588 19372 262640 19378
rect 262588 19314 262640 19320
rect 262600 14822 262628 19314
rect 263704 14890 263732 335582
rect 263692 14884 263744 14890
rect 263692 14826 263744 14832
rect 262588 14816 262640 14822
rect 262588 14758 262640 14764
rect 263796 10674 263824 340054
rect 264256 335646 264284 340054
rect 264992 337210 265020 340068
rect 265176 340054 265466 340082
rect 265544 340054 265926 340082
rect 264980 337204 265032 337210
rect 264980 337146 265032 337152
rect 264244 335640 264296 335646
rect 264244 335582 264296 335588
rect 265072 334348 265124 334354
rect 265072 334290 265124 334296
rect 265084 14958 265112 334290
rect 265072 14952 265124 14958
rect 265072 14894 265124 14900
rect 265176 10742 265204 340054
rect 265544 334354 265572 340054
rect 266372 337958 266400 340068
rect 266556 340054 266846 340082
rect 267016 340054 267306 340082
rect 266360 337952 266412 337958
rect 266360 337894 266412 337900
rect 266452 335640 266504 335646
rect 266452 335582 266504 335588
rect 265532 334348 265584 334354
rect 265532 334290 265584 334296
rect 266464 15026 266492 335582
rect 266452 15020 266504 15026
rect 266452 14962 266504 14968
rect 266556 10810 266584 340054
rect 267016 335646 267044 340054
rect 267660 337142 267688 340068
rect 267936 340054 268134 340082
rect 268304 340054 268594 340082
rect 268672 340054 269054 340082
rect 269316 340054 269514 340082
rect 269592 340054 269974 340082
rect 267648 337136 267700 337142
rect 267648 337078 267700 337084
rect 267004 335640 267056 335646
rect 267004 335582 267056 335588
rect 267832 335640 267884 335646
rect 267832 335582 267884 335588
rect 267004 328500 267056 328506
rect 267004 328442 267056 328448
rect 267016 328386 267044 328442
rect 267016 328358 267136 328386
rect 267108 321638 267136 328358
rect 267096 321632 267148 321638
rect 267096 321574 267148 321580
rect 267004 321428 267056 321434
rect 267004 321370 267056 321376
rect 267016 311930 267044 321370
rect 266924 311902 267044 311930
rect 266924 309194 266952 311902
rect 266912 309188 266964 309194
rect 266912 309130 266964 309136
rect 267004 309188 267056 309194
rect 267004 309130 267056 309136
rect 267016 309058 267044 309130
rect 267004 309052 267056 309058
rect 267004 308994 267056 309000
rect 267280 299532 267332 299538
rect 267280 299474 267332 299480
rect 267292 292602 267320 299474
rect 267004 292596 267056 292602
rect 267004 292538 267056 292544
rect 267280 292596 267332 292602
rect 267280 292538 267332 292544
rect 267016 289814 267044 292538
rect 267004 289808 267056 289814
rect 267004 289750 267056 289756
rect 267280 289808 267332 289814
rect 267280 289750 267332 289756
rect 267292 270745 267320 289750
rect 267278 270736 267334 270745
rect 267278 270671 267334 270680
rect 267002 270600 267058 270609
rect 267002 270535 267058 270544
rect 267016 269113 267044 270535
rect 267002 269104 267058 269113
rect 267002 269039 267058 269048
rect 267186 269104 267242 269113
rect 267186 269039 267242 269048
rect 267200 259486 267228 269039
rect 267188 259480 267240 259486
rect 267188 259422 267240 259428
rect 267280 259480 267332 259486
rect 267280 259422 267332 259428
rect 267292 249830 267320 259422
rect 267004 249824 267056 249830
rect 267004 249766 267056 249772
rect 267280 249824 267332 249830
rect 267280 249766 267332 249772
rect 267016 241534 267044 249766
rect 267004 241528 267056 241534
rect 267004 241470 267056 241476
rect 267004 241392 267056 241398
rect 267004 241334 267056 241340
rect 267016 230518 267044 241334
rect 266820 230512 266872 230518
rect 267004 230512 267056 230518
rect 266872 230460 266952 230466
rect 266820 230454 266952 230460
rect 267004 230454 267056 230460
rect 266832 230438 266952 230454
rect 266924 220862 266952 230438
rect 266912 220856 266964 220862
rect 266912 220798 266964 220804
rect 267004 220856 267056 220862
rect 267004 220798 267056 220804
rect 267016 215354 267044 220798
rect 267004 215348 267056 215354
rect 267004 215290 267056 215296
rect 267004 212560 267056 212566
rect 267004 212502 267056 212508
rect 267016 211138 267044 212502
rect 267004 211132 267056 211138
rect 267004 211074 267056 211080
rect 267096 202836 267148 202842
rect 267096 202778 267148 202784
rect 267108 200122 267136 202778
rect 267096 200116 267148 200122
rect 267096 200058 267148 200064
rect 267004 190528 267056 190534
rect 267004 190470 267056 190476
rect 267016 186946 267044 190470
rect 267016 186918 267136 186946
rect 267108 174010 267136 186918
rect 267096 174004 267148 174010
rect 267096 173946 267148 173952
rect 267004 173936 267056 173942
rect 267004 173878 267056 173884
rect 267016 164257 267044 173878
rect 267002 164248 267058 164257
rect 267002 164183 267058 164192
rect 267278 164112 267334 164121
rect 267278 164047 267334 164056
rect 267292 154601 267320 164047
rect 267002 154592 267058 154601
rect 267002 154527 267058 154536
rect 267278 154592 267334 154601
rect 267278 154527 267334 154536
rect 267016 147642 267044 154527
rect 267016 147614 267228 147642
rect 267200 138106 267228 147614
rect 267188 138100 267240 138106
rect 267188 138042 267240 138048
rect 267096 137964 267148 137970
rect 267096 137906 267148 137912
rect 267108 135250 267136 137906
rect 267096 135244 267148 135250
rect 267096 135186 267148 135192
rect 267096 128308 267148 128314
rect 267096 128250 267148 128256
rect 267108 125610 267136 128250
rect 267108 125582 267228 125610
rect 267200 118726 267228 125582
rect 267004 118720 267056 118726
rect 267004 118662 267056 118668
rect 267188 118720 267240 118726
rect 267188 118662 267240 118668
rect 267016 115938 267044 118662
rect 267004 115932 267056 115938
rect 267004 115874 267056 115880
rect 267188 115932 267240 115938
rect 267188 115874 267240 115880
rect 267200 108746 267228 115874
rect 267108 108718 267228 108746
rect 267108 102134 267136 108718
rect 267096 102128 267148 102134
rect 267096 102070 267148 102076
rect 267096 82884 267148 82890
rect 267096 82826 267148 82832
rect 267108 77994 267136 82826
rect 267096 77988 267148 77994
rect 267096 77930 267148 77936
rect 267096 67652 267148 67658
rect 267096 67594 267148 67600
rect 267108 61130 267136 67594
rect 267096 61124 267148 61130
rect 267096 61066 267148 61072
rect 267004 56636 267056 56642
rect 267004 56578 267056 56584
rect 267016 56114 267044 56578
rect 267016 56086 267228 56114
rect 267200 48278 267228 56086
rect 267188 48272 267240 48278
rect 267188 48214 267240 48220
rect 267096 38684 267148 38690
rect 267096 38626 267148 38632
rect 267108 37262 267136 38626
rect 267096 37256 267148 37262
rect 267096 37198 267148 37204
rect 267004 27668 267056 27674
rect 267004 27610 267056 27616
rect 267016 19281 267044 27610
rect 267002 19272 267058 19281
rect 267002 19207 267058 19216
rect 267278 19136 267334 19145
rect 267278 19071 267334 19080
rect 266544 10804 266596 10810
rect 266544 10746 266596 10752
rect 265164 10736 265216 10742
rect 265164 10678 265216 10684
rect 263784 10668 263836 10674
rect 263784 10610 263836 10616
rect 262404 8220 262456 8226
rect 262404 8162 262456 8168
rect 267004 8220 267056 8226
rect 267004 8162 267056 8168
rect 261024 8152 261076 8158
rect 261024 8094 261076 8100
rect 263416 8152 263468 8158
rect 263416 8094 263468 8100
rect 259736 8084 259788 8090
rect 259736 8026 259788 8032
rect 259828 8084 259880 8090
rect 259828 8026 259880 8032
rect 258816 2848 258868 2854
rect 258816 2790 258868 2796
rect 259840 480 259868 8026
rect 261024 6316 261076 6322
rect 261024 6258 261076 6264
rect 261036 480 261064 6258
rect 262220 3800 262272 3806
rect 262220 3742 262272 3748
rect 262232 480 262260 3742
rect 263428 480 263456 8094
rect 265808 4004 265860 4010
rect 265808 3946 265860 3952
rect 264612 3732 264664 3738
rect 264612 3674 264664 3680
rect 264624 480 264652 3674
rect 265820 480 265848 3946
rect 267016 480 267044 8162
rect 267292 4350 267320 19071
rect 267844 15094 267872 335582
rect 267832 15088 267884 15094
rect 267832 15030 267884 15036
rect 267936 10878 267964 340054
rect 268304 335646 268332 340054
rect 268672 337414 268700 340054
rect 268660 337408 268712 337414
rect 268660 337350 268712 337356
rect 269028 337408 269080 337414
rect 269028 337350 269080 337356
rect 268292 335640 268344 335646
rect 268292 335582 268344 335588
rect 267924 10872 267976 10878
rect 267924 10814 267976 10820
rect 267280 4344 267332 4350
rect 267280 4286 267332 4292
rect 269040 4146 269068 337350
rect 269212 335640 269264 335646
rect 269212 335582 269264 335588
rect 269118 134192 269174 134201
rect 269118 134127 269120 134136
rect 269172 134127 269174 134136
rect 269120 134098 269172 134104
rect 269224 15162 269252 335582
rect 269212 15156 269264 15162
rect 269212 15098 269264 15104
rect 269316 10946 269344 340054
rect 269592 335646 269620 340054
rect 270420 337074 270448 340068
rect 270696 340054 270894 340082
rect 270592 338428 270644 338434
rect 270592 338370 270644 338376
rect 270408 337068 270460 337074
rect 270408 337010 270460 337016
rect 269580 335640 269632 335646
rect 269580 335582 269632 335588
rect 270500 180872 270552 180878
rect 270498 180840 270500 180849
rect 270552 180840 270554 180849
rect 270498 180775 270554 180784
rect 270500 40384 270552 40390
rect 270498 40352 270500 40361
rect 270552 40352 270554 40361
rect 270498 40287 270554 40296
rect 270500 29232 270552 29238
rect 270498 29200 270500 29209
rect 270552 29200 270554 29209
rect 270498 29135 270554 29144
rect 270604 14414 270632 338370
rect 270592 14408 270644 14414
rect 270592 14350 270644 14356
rect 270696 11014 270724 340054
rect 271248 338434 271276 340068
rect 271236 338428 271288 338434
rect 271236 338370 271288 338376
rect 271708 337482 271736 340068
rect 272076 340054 272182 340082
rect 272352 340054 272642 340082
rect 271696 337476 271748 337482
rect 271696 337418 271748 337424
rect 271788 337476 271840 337482
rect 271788 337418 271840 337424
rect 270684 11008 270736 11014
rect 270684 10950 270736 10956
rect 269304 10940 269356 10946
rect 269304 10882 269356 10888
rect 268108 4140 268160 4146
rect 268108 4082 268160 4088
rect 269028 4140 269080 4146
rect 269028 4082 269080 4088
rect 268120 480 268148 4082
rect 269304 4072 269356 4078
rect 269304 4014 269356 4020
rect 269316 480 269344 4014
rect 271800 3874 271828 337418
rect 271972 335640 272024 335646
rect 271972 335582 272024 335588
rect 271984 14346 272012 335582
rect 271972 14340 272024 14346
rect 271972 14282 272024 14288
rect 272076 10266 272104 340054
rect 272352 335646 272380 340054
rect 273088 337550 273116 340068
rect 273076 337544 273128 337550
rect 273076 337486 273128 337492
rect 272340 335640 272392 335646
rect 272340 335582 272392 335588
rect 273548 335442 273576 340068
rect 273640 340054 274022 340082
rect 273536 335436 273588 335442
rect 273536 335378 273588 335384
rect 273444 335232 273496 335238
rect 273444 335174 273496 335180
rect 273352 333328 273404 333334
rect 273352 333270 273404 333276
rect 273364 215286 273392 333270
rect 273352 215280 273404 215286
rect 273352 215222 273404 215228
rect 273352 196036 273404 196042
rect 273352 195978 273404 195984
rect 272982 63880 273038 63889
rect 273166 63880 273222 63889
rect 273038 63838 273166 63866
rect 272982 63815 273038 63824
rect 273166 63815 273222 63824
rect 273364 60722 273392 195978
rect 273352 60716 273404 60722
rect 273352 60658 273404 60664
rect 273260 38684 273312 38690
rect 273260 38626 273312 38632
rect 273272 31634 273300 38626
rect 273272 31606 273392 31634
rect 273364 14278 273392 31606
rect 273352 14272 273404 14278
rect 273352 14214 273404 14220
rect 272064 10260 272116 10266
rect 272064 10202 272116 10208
rect 273456 10198 273484 335174
rect 273640 333334 273668 340054
rect 273902 337376 273958 337385
rect 273902 337311 273958 337320
rect 273628 333328 273680 333334
rect 273628 333270 273680 333276
rect 273536 215280 273588 215286
rect 273536 215222 273588 215228
rect 273548 196042 273576 215222
rect 273536 196036 273588 196042
rect 273536 195978 273588 195984
rect 273536 60648 273588 60654
rect 273536 60590 273588 60596
rect 273548 38690 273576 60590
rect 273536 38684 273588 38690
rect 273536 38626 273588 38632
rect 273444 10192 273496 10198
rect 273444 10134 273496 10140
rect 272892 4004 272944 4010
rect 272892 3946 272944 3952
rect 270500 3868 270552 3874
rect 270500 3810 270552 3816
rect 271788 3868 271840 3874
rect 271788 3810 271840 3816
rect 270512 480 270540 3810
rect 271696 2984 271748 2990
rect 271696 2926 271748 2932
rect 271708 480 271736 2926
rect 272904 480 272932 3946
rect 273916 2990 273944 337311
rect 274468 336938 274496 340068
rect 274548 337544 274600 337550
rect 274548 337486 274600 337492
rect 274456 336932 274508 336938
rect 274456 336874 274508 336880
rect 273994 29336 274050 29345
rect 273994 29271 274050 29280
rect 274008 29238 274036 29271
rect 273996 29232 274048 29238
rect 273996 29174 274048 29180
rect 274560 4146 274588 337486
rect 274732 335640 274784 335646
rect 274732 335582 274784 335588
rect 274744 14210 274772 335582
rect 274732 14204 274784 14210
rect 274732 14146 274784 14152
rect 274836 10130 274864 340068
rect 274928 340054 275310 340082
rect 274928 335646 274956 340054
rect 275756 337618 275784 340068
rect 275744 337612 275796 337618
rect 275744 337554 275796 337560
rect 274916 335640 274968 335646
rect 274916 335582 274968 335588
rect 276112 186380 276164 186386
rect 276112 186322 276164 186328
rect 275374 181112 275430 181121
rect 275374 181047 275430 181056
rect 275388 180878 275416 181047
rect 275376 180872 275428 180878
rect 275376 180814 275428 180820
rect 276124 176662 276152 186322
rect 276112 176656 276164 176662
rect 276112 176598 276164 176604
rect 275376 134156 275428 134162
rect 275376 134098 275428 134104
rect 275388 134065 275416 134098
rect 275374 134056 275430 134065
rect 275374 133991 275430 134000
rect 276112 70440 276164 70446
rect 276112 70382 276164 70388
rect 276124 14142 276152 70382
rect 276112 14136 276164 14142
rect 276112 14078 276164 14084
rect 274824 10124 274876 10130
rect 274824 10066 274876 10072
rect 276216 10062 276244 340068
rect 276308 340054 276690 340082
rect 276308 186454 276336 340054
rect 276756 337748 276808 337754
rect 276756 337690 276808 337696
rect 276664 337612 276716 337618
rect 276664 337554 276716 337560
rect 276296 186448 276348 186454
rect 276296 186390 276348 186396
rect 276296 176588 276348 176594
rect 276296 176530 276348 176536
rect 276308 70514 276336 176530
rect 276296 70508 276348 70514
rect 276296 70450 276348 70456
rect 276204 10056 276256 10062
rect 276204 9998 276256 10004
rect 276676 4146 276704 337554
rect 274088 4140 274140 4146
rect 274088 4082 274140 4088
rect 274548 4140 274600 4146
rect 274548 4082 274600 4088
rect 275284 4140 275336 4146
rect 275284 4082 275336 4088
rect 276664 4140 276716 4146
rect 276664 4082 276716 4088
rect 273904 2984 273956 2990
rect 273904 2926 273956 2932
rect 274100 480 274128 4082
rect 275296 480 275324 4082
rect 276768 3890 276796 337690
rect 277136 336802 277164 340068
rect 277124 336796 277176 336802
rect 277124 336738 277176 336744
rect 277400 335708 277452 335714
rect 277400 335650 277452 335656
rect 277412 8294 277440 335650
rect 277492 335640 277544 335646
rect 277492 335582 277544 335588
rect 277504 11898 277532 335582
rect 277492 11892 277544 11898
rect 277492 11834 277544 11840
rect 277596 11830 277624 340068
rect 277688 340054 278070 340082
rect 278148 340054 278438 340082
rect 278792 340054 278898 340082
rect 279068 340054 279358 340082
rect 279528 340054 279818 340082
rect 280172 340054 280278 340082
rect 280356 340054 280738 340082
rect 280908 340054 281198 340082
rect 281552 340054 281658 340082
rect 281828 340054 282118 340082
rect 282196 340054 282486 340082
rect 282946 340054 283144 340082
rect 277688 335646 277716 340054
rect 278148 335714 278176 340054
rect 278136 335708 278188 335714
rect 278136 335650 278188 335656
rect 277676 335640 277728 335646
rect 277676 335582 277728 335588
rect 277584 11824 277636 11830
rect 277584 11766 277636 11772
rect 277400 8288 277452 8294
rect 277400 8230 277452 8236
rect 278792 5370 278820 340054
rect 278964 335640 279016 335646
rect 278964 335582 279016 335588
rect 278976 8945 279004 335582
rect 278962 8936 279018 8945
rect 278962 8871 279018 8880
rect 279068 6594 279096 340054
rect 279528 335646 279556 340054
rect 279976 337340 280028 337346
rect 279976 337282 280028 337288
rect 279516 335640 279568 335646
rect 279516 335582 279568 335588
rect 279056 6588 279108 6594
rect 279056 6530 279108 6536
rect 278780 5364 278832 5370
rect 278780 5306 278832 5312
rect 279988 4146 280016 337282
rect 280172 5438 280200 340054
rect 280252 63504 280304 63510
rect 280252 63446 280304 63452
rect 280264 44538 280292 63446
rect 280252 44532 280304 44538
rect 280252 44474 280304 44480
rect 280356 13258 280384 340054
rect 280908 331242 280936 340054
rect 280632 331214 280936 331242
rect 280632 318850 280660 331214
rect 280528 318844 280580 318850
rect 280528 318786 280580 318792
rect 280620 318844 280672 318850
rect 280620 318786 280672 318792
rect 280540 311930 280568 318786
rect 280540 311902 280660 311930
rect 280632 302258 280660 311902
rect 280436 302252 280488 302258
rect 280436 302194 280488 302200
rect 280620 302252 280672 302258
rect 280620 302194 280672 302200
rect 280448 302138 280476 302194
rect 280448 302110 280568 302138
rect 280540 292618 280568 302110
rect 280540 292590 280660 292618
rect 280632 282946 280660 292590
rect 280436 282940 280488 282946
rect 280436 282882 280488 282888
rect 280620 282940 280672 282946
rect 280620 282882 280672 282888
rect 280448 282826 280476 282882
rect 280448 282798 280568 282826
rect 280540 273306 280568 282798
rect 280540 273278 280660 273306
rect 280632 263634 280660 273278
rect 280436 263628 280488 263634
rect 280436 263570 280488 263576
rect 280620 263628 280672 263634
rect 280620 263570 280672 263576
rect 280448 263514 280476 263570
rect 280448 263486 280568 263514
rect 280540 253994 280568 263486
rect 280540 253966 280660 253994
rect 280632 234734 280660 253966
rect 280620 234728 280672 234734
rect 280620 234670 280672 234676
rect 280528 234592 280580 234598
rect 280528 234534 280580 234540
rect 280540 225026 280568 234534
rect 280448 224998 280568 225026
rect 280448 224890 280476 224998
rect 280448 224862 280568 224890
rect 280540 205714 280568 224862
rect 280448 205686 280568 205714
rect 280448 205578 280476 205686
rect 280448 205550 280568 205578
rect 280540 186402 280568 205550
rect 280448 186374 280568 186402
rect 280448 186318 280476 186374
rect 280436 186312 280488 186318
rect 280436 186254 280488 186260
rect 280620 186312 280672 186318
rect 280620 186254 280672 186260
rect 280632 176746 280660 186254
rect 280632 176718 280752 176746
rect 280724 176610 280752 176718
rect 280540 176582 280752 176610
rect 280540 167090 280568 176582
rect 280448 167062 280568 167090
rect 280448 166954 280476 167062
rect 280448 166926 280568 166954
rect 280540 157418 280568 166926
rect 280528 157412 280580 157418
rect 280528 157354 280580 157360
rect 280620 157276 280672 157282
rect 280620 157218 280672 157224
rect 280632 147694 280660 157218
rect 280436 147688 280488 147694
rect 280620 147688 280672 147694
rect 280488 147636 280568 147642
rect 280436 147630 280568 147636
rect 280620 147630 280672 147636
rect 280448 147614 280568 147630
rect 280540 128466 280568 147614
rect 280448 128438 280568 128466
rect 280448 128330 280476 128438
rect 280448 128302 280568 128330
rect 280540 118726 280568 128302
rect 280528 118720 280580 118726
rect 280528 118662 280580 118668
rect 280620 118652 280672 118658
rect 280620 118594 280672 118600
rect 280632 109070 280660 118594
rect 280436 109064 280488 109070
rect 280620 109064 280672 109070
rect 280488 109012 280568 109018
rect 280436 109006 280568 109012
rect 280620 109006 280672 109012
rect 280448 108990 280568 109006
rect 280540 104854 280568 108990
rect 280528 104848 280580 104854
rect 280528 104790 280580 104796
rect 280620 95260 280672 95266
rect 280620 95202 280672 95208
rect 280632 89758 280660 95202
rect 280436 89752 280488 89758
rect 280620 89752 280672 89758
rect 280488 89700 280620 89706
rect 280436 89694 280672 89700
rect 280448 89678 280660 89694
rect 280632 73234 280660 89678
rect 280528 73228 280580 73234
rect 280528 73170 280580 73176
rect 280620 73228 280672 73234
rect 280620 73170 280672 73176
rect 280540 63510 280568 73170
rect 280528 63504 280580 63510
rect 280528 63446 280580 63452
rect 280528 40384 280580 40390
rect 280526 40352 280528 40361
rect 280580 40352 280582 40361
rect 280526 40287 280582 40296
rect 280528 28892 280580 28898
rect 280528 28834 280580 28840
rect 280540 18018 280568 28834
rect 280436 18012 280488 18018
rect 280436 17954 280488 17960
rect 280528 18012 280580 18018
rect 280528 17954 280580 17960
rect 280344 13252 280396 13258
rect 280344 13194 280396 13200
rect 280448 9246 280476 17954
rect 280436 9240 280488 9246
rect 280436 9182 280488 9188
rect 281552 5506 281580 340054
rect 281724 335640 281776 335646
rect 281724 335582 281776 335588
rect 281736 9314 281764 335582
rect 281724 9308 281776 9314
rect 281724 9250 281776 9256
rect 281828 7546 281856 340054
rect 282196 335646 282224 340054
rect 282184 335640 282236 335646
rect 282184 335582 282236 335588
rect 283012 335640 283064 335646
rect 283012 335582 283064 335588
rect 282734 134056 282790 134065
rect 282918 134056 282974 134065
rect 282790 134014 282918 134042
rect 282734 133991 282790 134000
rect 282918 133991 282974 134000
rect 282826 87272 282882 87281
rect 282826 87207 282828 87216
rect 282880 87207 282882 87216
rect 282828 87178 282880 87184
rect 283024 9382 283052 335582
rect 283116 11966 283144 340054
rect 283208 340054 283406 340082
rect 283576 340054 283866 340082
rect 284326 340054 284524 340082
rect 283104 11960 283156 11966
rect 283104 11902 283156 11908
rect 283012 9376 283064 9382
rect 283012 9318 283064 9324
rect 281816 7540 281868 7546
rect 281816 7482 281868 7488
rect 283208 7478 283236 340054
rect 283576 335646 283604 340054
rect 283564 335640 283616 335646
rect 283564 335582 283616 335588
rect 284392 333192 284444 333198
rect 284392 333134 284444 333140
rect 284404 9450 284432 333134
rect 284496 12034 284524 340054
rect 284588 340054 284786 340082
rect 284864 340054 285246 340082
rect 285706 340054 285996 340082
rect 284484 12028 284536 12034
rect 284484 11970 284536 11976
rect 284392 9444 284444 9450
rect 284392 9386 284444 9392
rect 283196 7472 283248 7478
rect 283196 7414 283248 7420
rect 284588 7410 284616 340054
rect 284864 333198 284892 340054
rect 285588 337816 285640 337822
rect 285588 337758 285640 337764
rect 284852 333192 284904 333198
rect 284852 333134 284904 333140
rect 284942 29336 284998 29345
rect 284942 29271 284998 29280
rect 284956 29073 284984 29271
rect 284942 29064 284998 29073
rect 284942 28999 284998 29008
rect 284576 7404 284628 7410
rect 284576 7346 284628 7352
rect 284208 6384 284260 6390
rect 284208 6326 284260 6332
rect 281540 5500 281592 5506
rect 281540 5442 281592 5448
rect 280160 5432 280212 5438
rect 280160 5374 280212 5380
rect 283656 5364 283708 5370
rect 283656 5306 283708 5312
rect 280068 5296 280120 5302
rect 280068 5238 280120 5244
rect 278872 4140 278924 4146
rect 278872 4082 278924 4088
rect 279976 4140 280028 4146
rect 279976 4082 280028 4088
rect 276400 3862 276796 3890
rect 276400 3738 276428 3862
rect 276388 3732 276440 3738
rect 276388 3674 276440 3680
rect 276480 3732 276532 3738
rect 276480 3674 276532 3680
rect 276492 480 276520 3674
rect 277676 3664 277728 3670
rect 277676 3606 277728 3612
rect 277688 480 277716 3606
rect 278884 480 278912 4082
rect 280080 480 280108 5238
rect 281264 4140 281316 4146
rect 281264 4082 281316 4088
rect 281276 480 281304 4082
rect 282460 3188 282512 3194
rect 282460 3130 282512 3136
rect 282472 480 282500 3130
rect 283668 480 283696 5306
rect 284220 3738 284248 6326
rect 285600 4146 285628 337758
rect 285864 335708 285916 335714
rect 285864 335650 285916 335656
rect 285772 335640 285824 335646
rect 285772 335582 285824 335588
rect 285784 9518 285812 335582
rect 285876 12170 285904 335650
rect 285864 12164 285916 12170
rect 285864 12106 285916 12112
rect 285968 12102 285996 340054
rect 285956 12096 286008 12102
rect 285956 12038 286008 12044
rect 285772 9512 285824 9518
rect 285772 9454 285824 9460
rect 286060 7342 286088 340068
rect 286152 340054 286534 340082
rect 286704 340054 286994 340082
rect 287072 340054 287454 340082
rect 287532 340054 287914 340082
rect 287992 340054 288374 340082
rect 288452 340054 288834 340082
rect 288912 340054 289294 340082
rect 289556 340054 289662 340082
rect 289832 340054 290122 340082
rect 290200 340054 290582 340082
rect 290660 340054 291042 340082
rect 291212 340054 291502 340082
rect 291580 340054 291962 340082
rect 292132 340054 292422 340082
rect 292592 340054 292882 340082
rect 292960 340054 293342 340082
rect 293604 340054 293710 340082
rect 293972 340054 294170 340082
rect 294248 340054 294630 340082
rect 294800 340054 295090 340082
rect 295352 340054 295550 340082
rect 295628 340054 296010 340082
rect 296088 340054 296470 340082
rect 296732 340054 296930 340082
rect 297008 340054 297298 340082
rect 297376 340054 297758 340082
rect 298112 340054 298218 340082
rect 298296 340054 298678 340082
rect 298940 340054 299138 340082
rect 299492 340054 299598 340082
rect 299676 340054 300058 340082
rect 300228 340054 300518 340082
rect 286152 335646 286180 340054
rect 286704 335714 286732 340054
rect 286692 335708 286744 335714
rect 286692 335650 286744 335656
rect 286140 335640 286192 335646
rect 286140 335582 286192 335588
rect 286048 7336 286100 7342
rect 286048 7278 286100 7284
rect 287072 7274 287100 340054
rect 287532 335594 287560 340054
rect 287164 335566 287560 335594
rect 287164 9994 287192 335566
rect 287992 334354 288020 340054
rect 288072 337340 288124 337346
rect 288072 337282 288124 337288
rect 287980 334348 288032 334354
rect 287980 334290 288032 334296
rect 288084 334234 288112 337282
rect 287716 334206 288112 334234
rect 287428 327140 287480 327146
rect 287428 327082 287480 327088
rect 287440 318866 287468 327082
rect 287348 318838 287468 318866
rect 287348 317422 287376 318838
rect 287336 317416 287388 317422
rect 287336 317358 287388 317364
rect 287336 311840 287388 311846
rect 287336 311782 287388 311788
rect 287348 299470 287376 311782
rect 287336 299464 287388 299470
rect 287336 299406 287388 299412
rect 287336 289876 287388 289882
rect 287336 289818 287388 289824
rect 287348 280158 287376 289818
rect 287336 280152 287388 280158
rect 287336 280094 287388 280100
rect 287336 270564 287388 270570
rect 287336 270506 287388 270512
rect 287348 260846 287376 270506
rect 287336 260840 287388 260846
rect 287336 260782 287388 260788
rect 287336 251252 287388 251258
rect 287336 251194 287388 251200
rect 287348 234598 287376 251194
rect 287336 234592 287388 234598
rect 287336 234534 287388 234540
rect 287336 234456 287388 234462
rect 287336 234398 287388 234404
rect 287348 222193 287376 234398
rect 287334 222184 287390 222193
rect 287334 222119 287390 222128
rect 287518 222184 287574 222193
rect 287518 222119 287574 222128
rect 287532 212566 287560 222119
rect 287336 212560 287388 212566
rect 287336 212502 287388 212508
rect 287520 212560 287572 212566
rect 287520 212502 287572 212508
rect 287348 202881 287376 212502
rect 287334 202872 287390 202881
rect 287334 202807 287390 202816
rect 287518 202872 287574 202881
rect 287518 202807 287574 202816
rect 287532 193254 287560 202807
rect 287336 193248 287388 193254
rect 287336 193190 287388 193196
rect 287520 193248 287572 193254
rect 287520 193190 287572 193196
rect 287348 183546 287376 193190
rect 287256 183518 287376 183546
rect 287256 176730 287284 183518
rect 287244 176724 287296 176730
rect 287244 176666 287296 176672
rect 287336 176656 287388 176662
rect 287336 176598 287388 176604
rect 287348 164218 287376 176598
rect 287336 164212 287388 164218
rect 287336 164154 287388 164160
rect 287336 154624 287388 154630
rect 287336 154566 287388 154572
rect 287348 145042 287376 154566
rect 287244 145036 287296 145042
rect 287244 144978 287296 144984
rect 287336 145036 287388 145042
rect 287336 144978 287388 144984
rect 287256 143546 287284 144978
rect 287244 143540 287296 143546
rect 287244 143482 287296 143488
rect 287428 137828 287480 137834
rect 287428 137770 287480 137776
rect 287440 133906 287468 137770
rect 287348 133890 287468 133906
rect 287336 133884 287468 133890
rect 287388 133878 287468 133884
rect 287520 133884 287572 133890
rect 287336 133826 287388 133832
rect 287520 133826 287572 133832
rect 287348 133795 287376 133826
rect 287532 124273 287560 133826
rect 287242 124264 287298 124273
rect 287242 124199 287298 124208
rect 287518 124264 287574 124273
rect 287518 124199 287574 124208
rect 287256 124166 287284 124199
rect 287244 124160 287296 124166
rect 287244 124102 287296 124108
rect 287428 124092 287480 124098
rect 287428 124034 287480 124040
rect 287440 115818 287468 124034
rect 287348 115790 287468 115818
rect 287348 114510 287376 115790
rect 287336 114504 287388 114510
rect 287336 114446 287388 114452
rect 287336 104916 287388 104922
rect 287336 104858 287388 104864
rect 287348 99498 287376 104858
rect 287348 99470 287468 99498
rect 287440 85610 287468 99470
rect 287336 85604 287388 85610
rect 287336 85546 287388 85552
rect 287428 85604 287480 85610
rect 287428 85546 287480 85552
rect 287348 80170 287376 85546
rect 287336 80164 287388 80170
rect 287336 80106 287388 80112
rect 287336 80028 287388 80034
rect 287336 79970 287388 79976
rect 287348 70514 287376 79970
rect 287336 70508 287388 70514
rect 287336 70450 287388 70456
rect 287336 70372 287388 70378
rect 287336 70314 287388 70320
rect 287348 67697 287376 70314
rect 287334 67688 287390 67697
rect 287334 67623 287390 67632
rect 287426 67552 287482 67561
rect 287426 67487 287482 67496
rect 287440 58002 287468 67487
rect 287336 57996 287388 58002
rect 287336 57938 287388 57944
rect 287428 57996 287480 58002
rect 287428 57938 287480 57944
rect 287348 51270 287376 57938
rect 287336 51264 287388 51270
rect 287336 51206 287388 51212
rect 287244 51060 287296 51066
rect 287244 51002 287296 51008
rect 287256 38758 287284 51002
rect 287244 38752 287296 38758
rect 287244 38694 287296 38700
rect 287244 38616 287296 38622
rect 287244 38558 287296 38564
rect 287256 28937 287284 38558
rect 287242 28928 287298 28937
rect 287242 28863 287298 28872
rect 287334 28792 287390 28801
rect 287334 28727 287390 28736
rect 287348 13326 287376 28727
rect 287336 13320 287388 13326
rect 287336 13262 287388 13268
rect 287152 9988 287204 9994
rect 287152 9930 287204 9936
rect 287060 7268 287112 7274
rect 287060 7210 287112 7216
rect 287152 5432 287204 5438
rect 287152 5374 287204 5380
rect 284760 4140 284812 4146
rect 284760 4082 284812 4088
rect 285588 4140 285640 4146
rect 285588 4082 285640 4088
rect 284208 3732 284260 3738
rect 284208 3674 284260 3680
rect 284772 480 284800 4082
rect 285956 3732 286008 3738
rect 285956 3674 286008 3680
rect 285968 480 285996 3674
rect 287164 480 287192 5374
rect 287716 3670 287744 334206
rect 288452 7206 288480 340054
rect 288912 335594 288940 340054
rect 288544 335566 288940 335594
rect 288544 9926 288572 335566
rect 289556 328506 289584 340054
rect 288808 328500 288860 328506
rect 288808 328442 288860 328448
rect 289544 328500 289596 328506
rect 289544 328442 289596 328448
rect 288820 311930 288848 328442
rect 288728 311902 288848 311930
rect 288728 302326 288756 311902
rect 288716 302320 288768 302326
rect 288716 302262 288768 302268
rect 288716 302184 288768 302190
rect 288716 302126 288768 302132
rect 288728 299520 288756 302126
rect 288728 299492 288848 299520
rect 288820 299441 288848 299492
rect 288806 299432 288862 299441
rect 288806 299367 288862 299376
rect 288990 299432 289046 299441
rect 288990 299367 289046 299376
rect 289004 289882 289032 299367
rect 288716 289876 288768 289882
rect 288716 289818 288768 289824
rect 288992 289876 289044 289882
rect 288992 289818 289044 289824
rect 288728 289746 288756 289818
rect 288716 289740 288768 289746
rect 288716 289682 288768 289688
rect 288716 282872 288768 282878
rect 288716 282814 288768 282820
rect 288728 280242 288756 282814
rect 288728 280214 288848 280242
rect 288820 280140 288848 280214
rect 288728 280112 288848 280140
rect 288728 273306 288756 280112
rect 288636 273278 288756 273306
rect 288636 270570 288664 273278
rect 288624 270564 288676 270570
rect 288624 270506 288676 270512
rect 288716 270564 288768 270570
rect 288716 270506 288768 270512
rect 288728 270434 288756 270506
rect 288716 270428 288768 270434
rect 288716 270370 288768 270376
rect 288716 263560 288768 263566
rect 288716 263502 288768 263508
rect 288728 260930 288756 263502
rect 288728 260902 288848 260930
rect 288820 260828 288848 260902
rect 288728 260800 288848 260828
rect 288728 253994 288756 260800
rect 288636 253966 288756 253994
rect 288636 251258 288664 253966
rect 288624 251252 288676 251258
rect 288624 251194 288676 251200
rect 288716 251252 288768 251258
rect 288716 251194 288768 251200
rect 288728 244322 288756 251194
rect 288716 244316 288768 244322
rect 288716 244258 288768 244264
rect 288808 244180 288860 244186
rect 288808 244122 288860 244128
rect 288820 241482 288848 244122
rect 288728 241454 288848 241482
rect 288728 240106 288756 241454
rect 288716 240100 288768 240106
rect 288716 240042 288768 240048
rect 288808 231872 288860 231878
rect 288808 231814 288860 231820
rect 288820 225010 288848 231814
rect 288808 225004 288860 225010
rect 288808 224946 288860 224952
rect 288808 224868 288860 224874
rect 288808 224810 288860 224816
rect 288820 222170 288848 224810
rect 288728 222142 288848 222170
rect 288728 215354 288756 222142
rect 288716 215348 288768 215354
rect 288716 215290 288768 215296
rect 288808 212560 288860 212566
rect 288808 212502 288860 212508
rect 288820 205698 288848 212502
rect 288808 205692 288860 205698
rect 288808 205634 288860 205640
rect 288820 202910 288848 202941
rect 288808 202904 288860 202910
rect 288728 202852 288808 202858
rect 288728 202846 288860 202852
rect 288728 202830 288848 202846
rect 288728 196042 288756 202830
rect 288716 196036 288768 196042
rect 288716 195978 288768 195984
rect 288808 193248 288860 193254
rect 288808 193190 288860 193196
rect 288820 186386 288848 193190
rect 288808 186380 288860 186386
rect 288808 186322 288860 186328
rect 288808 183592 288860 183598
rect 288808 183534 288860 183540
rect 288820 176798 288848 183534
rect 288808 176792 288860 176798
rect 288808 176734 288860 176740
rect 288808 176656 288860 176662
rect 288808 176598 288860 176604
rect 288820 162858 288848 176598
rect 288716 162852 288768 162858
rect 288716 162794 288768 162800
rect 288808 162852 288860 162858
rect 288808 162794 288860 162800
rect 288728 161430 288756 162794
rect 288716 161424 288768 161430
rect 288716 161366 288768 161372
rect 288808 153876 288860 153882
rect 288808 153818 288860 153824
rect 288820 149054 288848 153818
rect 288808 149048 288860 149054
rect 288808 148990 288860 148996
rect 288808 139528 288860 139534
rect 288808 139470 288860 139476
rect 288820 139398 288848 139470
rect 288808 139392 288860 139398
rect 288808 139334 288860 139340
rect 288900 139392 288952 139398
rect 288900 139334 288952 139340
rect 288912 128194 288940 139334
rect 288820 128166 288940 128194
rect 288820 114594 288848 128166
rect 288728 114566 288848 114594
rect 288728 114510 288756 114566
rect 288716 114504 288768 114510
rect 288716 114446 288768 114452
rect 288808 104916 288860 104922
rect 288808 104858 288860 104864
rect 288820 99482 288848 104858
rect 288808 99476 288860 99482
rect 288808 99418 288860 99424
rect 288624 86148 288676 86154
rect 288624 86090 288676 86096
rect 288636 73846 288664 86090
rect 288624 73840 288676 73846
rect 288624 73782 288676 73788
rect 288716 57996 288768 58002
rect 288716 57938 288768 57944
rect 288728 53122 288756 57938
rect 288728 53094 288940 53122
rect 288912 50946 288940 53094
rect 288820 50918 288940 50946
rect 288820 48278 288848 50918
rect 288624 48272 288676 48278
rect 288624 48214 288676 48220
rect 288808 48272 288860 48278
rect 288808 48214 288860 48220
rect 288636 38706 288664 48214
rect 288636 38678 288756 38706
rect 288728 33810 288756 38678
rect 288728 33782 289032 33810
rect 289004 19378 289032 33782
rect 288716 19372 288768 19378
rect 288716 19314 288768 19320
rect 288992 19372 289044 19378
rect 288992 19314 289044 19320
rect 288728 13394 288756 19314
rect 288716 13388 288768 13394
rect 288716 13330 288768 13336
rect 288532 9920 288584 9926
rect 288532 9862 288584 9868
rect 288440 7200 288492 7206
rect 288440 7142 288492 7148
rect 289832 7138 289860 340054
rect 290200 335594 290228 340054
rect 289924 335566 290228 335594
rect 289924 9858 289952 335566
rect 290464 329452 290516 329458
rect 290464 329394 290516 329400
rect 290004 328500 290056 328506
rect 290004 328442 290056 328448
rect 290016 321638 290044 328442
rect 290004 321632 290056 321638
rect 290004 321574 290056 321580
rect 290096 321496 290148 321502
rect 290096 321438 290148 321444
rect 290108 315926 290136 321438
rect 290096 315920 290148 315926
rect 290096 315862 290148 315868
rect 290280 307828 290332 307834
rect 290280 307770 290332 307776
rect 290292 299538 290320 307770
rect 290096 299532 290148 299538
rect 290096 299474 290148 299480
rect 290280 299532 290332 299538
rect 290280 299474 290332 299480
rect 290108 292482 290136 299474
rect 290016 292454 290136 292482
rect 290016 292210 290044 292454
rect 290016 292182 290136 292210
rect 290108 280158 290136 292182
rect 290096 280152 290148 280158
rect 290096 280094 290148 280100
rect 290096 273012 290148 273018
rect 290096 272954 290148 272960
rect 290108 260846 290136 272954
rect 290096 260840 290148 260846
rect 290096 260782 290148 260788
rect 290096 252884 290148 252890
rect 290096 252826 290148 252832
rect 290108 176610 290136 252826
rect 290016 176582 290136 176610
rect 290016 176338 290044 176582
rect 290016 176310 290136 176338
rect 290108 157434 290136 176310
rect 290108 157406 290228 157434
rect 290200 157332 290228 157406
rect 290108 157304 290228 157332
rect 290108 154562 290136 157304
rect 290096 154556 290148 154562
rect 290096 154498 290148 154504
rect 290188 154556 290240 154562
rect 290188 154498 290240 154504
rect 290200 135425 290228 154498
rect 290186 135416 290242 135425
rect 290186 135351 290242 135360
rect 290094 135280 290150 135289
rect 290094 135215 290150 135224
rect 290108 116090 290136 135215
rect 290108 116062 290228 116090
rect 290200 104938 290228 116062
rect 290108 104910 290228 104938
rect 290108 99482 290136 104910
rect 290096 99476 290148 99482
rect 290096 99418 290148 99424
rect 290096 99340 290148 99346
rect 290096 99282 290148 99288
rect 290108 75954 290136 99282
rect 290096 75948 290148 75954
rect 290096 75890 290148 75896
rect 290188 75812 290240 75818
rect 290188 75754 290240 75760
rect 290200 70922 290228 75754
rect 290004 70916 290056 70922
rect 290004 70858 290056 70864
rect 290188 70916 290240 70922
rect 290188 70858 290240 70864
rect 290016 56658 290044 70858
rect 290016 56630 290136 56658
rect 290108 55350 290136 56630
rect 290096 55344 290148 55350
rect 290096 55286 290148 55292
rect 290004 55276 290056 55282
rect 290004 55218 290056 55224
rect 290016 55146 290044 55218
rect 290004 55140 290056 55146
rect 290004 55082 290056 55088
rect 290004 45620 290056 45626
rect 290004 45562 290056 45568
rect 290016 37210 290044 45562
rect 290016 37182 290136 37210
rect 290108 35986 290136 37182
rect 290016 35958 290136 35986
rect 290016 35902 290044 35958
rect 290004 35896 290056 35902
rect 290004 35838 290056 35844
rect 290188 26308 290240 26314
rect 290188 26250 290240 26256
rect 290200 26058 290228 26250
rect 290108 26030 290228 26058
rect 290108 12510 290136 26030
rect 290096 12504 290148 12510
rect 290096 12446 290148 12452
rect 289912 9852 289964 9858
rect 289912 9794 289964 9800
rect 289820 7132 289872 7138
rect 289820 7074 289872 7080
rect 290476 3942 290504 329394
rect 290660 328506 290688 340054
rect 290648 328500 290700 328506
rect 290648 328442 290700 328448
rect 291212 6662 291240 340054
rect 291580 335594 291608 340054
rect 291304 335566 291608 335594
rect 291304 7070 291332 335566
rect 292132 328506 292160 340054
rect 292488 338088 292540 338094
rect 292488 338030 292540 338036
rect 291568 328500 291620 328506
rect 291568 328442 291620 328448
rect 292120 328500 292172 328506
rect 292120 328442 292172 328448
rect 291580 309194 291608 328442
rect 291476 309188 291528 309194
rect 291476 309130 291528 309136
rect 291568 309188 291620 309194
rect 291568 309130 291620 309136
rect 291488 304314 291516 309130
rect 291488 304286 291608 304314
rect 291580 299470 291608 304286
rect 291476 299464 291528 299470
rect 291476 299406 291528 299412
rect 291568 299464 291620 299470
rect 291568 299406 291620 299412
rect 291488 298110 291516 299406
rect 291476 298104 291528 298110
rect 291476 298046 291528 298052
rect 291476 288448 291528 288454
rect 291476 288390 291528 288396
rect 291488 285002 291516 288390
rect 291396 284974 291516 285002
rect 291396 282690 291424 284974
rect 291396 282662 291608 282690
rect 291580 280158 291608 282662
rect 291476 280152 291528 280158
rect 291476 280094 291528 280100
rect 291568 280152 291620 280158
rect 291568 280094 291620 280100
rect 291488 278769 291516 280094
rect 291474 278760 291530 278769
rect 291474 278695 291530 278704
rect 291658 278760 291714 278769
rect 291658 278695 291714 278704
rect 291672 269142 291700 278695
rect 291476 269136 291528 269142
rect 291476 269078 291528 269084
rect 291660 269136 291712 269142
rect 291660 269078 291712 269084
rect 291488 263634 291516 269078
rect 291476 263628 291528 263634
rect 291476 263570 291528 263576
rect 291568 263492 291620 263498
rect 291568 263434 291620 263440
rect 291580 260846 291608 263434
rect 291568 260840 291620 260846
rect 291568 260782 291620 260788
rect 291476 251320 291528 251326
rect 291476 251262 291528 251268
rect 291488 251190 291516 251262
rect 291476 251184 291528 251190
rect 291476 251126 291528 251132
rect 291568 241528 291620 241534
rect 291568 241470 291620 241476
rect 291580 233594 291608 241470
rect 291580 233566 291700 233594
rect 291672 230518 291700 233566
rect 291568 230512 291620 230518
rect 291566 230480 291568 230489
rect 291660 230512 291712 230518
rect 291620 230480 291622 230489
rect 291660 230454 291712 230460
rect 291750 230480 291806 230489
rect 291566 230415 291622 230424
rect 291750 230415 291806 230424
rect 291764 220930 291792 230415
rect 291384 220924 291436 220930
rect 291384 220866 291436 220872
rect 291752 220924 291804 220930
rect 291752 220866 291804 220872
rect 291396 220794 291424 220866
rect 291384 220788 291436 220794
rect 291384 220730 291436 220736
rect 291384 202972 291436 202978
rect 291384 202914 291436 202920
rect 291396 201482 291424 202914
rect 291384 201476 291436 201482
rect 291384 201418 291436 201424
rect 291660 201476 291712 201482
rect 291660 201418 291712 201424
rect 291672 186266 291700 201418
rect 291580 186238 291700 186266
rect 291580 183569 291608 186238
rect 291382 183560 291438 183569
rect 291382 183495 291438 183504
rect 291566 183560 291622 183569
rect 291566 183495 291622 183504
rect 291396 173942 291424 183495
rect 291384 173936 291436 173942
rect 291476 173936 291528 173942
rect 291384 173878 291436 173884
rect 291474 173904 291476 173913
rect 291528 173904 291530 173913
rect 291474 173839 291530 173848
rect 291750 173904 291806 173913
rect 291750 173839 291806 173848
rect 291764 164257 291792 173839
rect 291566 164248 291622 164257
rect 291566 164183 291622 164192
rect 291750 164248 291806 164257
rect 291750 164183 291806 164192
rect 291580 154737 291608 164183
rect 291566 154728 291622 154737
rect 291566 154663 291622 154672
rect 291658 154456 291714 154465
rect 291658 154391 291714 154400
rect 291672 147506 291700 154391
rect 291580 147478 291700 147506
rect 291580 135425 291608 147478
rect 291566 135416 291622 135425
rect 291566 135351 291622 135360
rect 291566 135144 291622 135153
rect 291566 135079 291622 135088
rect 291580 124234 291608 135079
rect 291568 124228 291620 124234
rect 291568 124170 291620 124176
rect 291568 121508 291620 121514
rect 291568 121450 291620 121456
rect 291580 102105 291608 121450
rect 291566 102096 291622 102105
rect 291566 102031 291622 102040
rect 291474 101960 291530 101969
rect 291474 101895 291530 101904
rect 291488 84250 291516 101895
rect 291476 84244 291528 84250
rect 291476 84186 291528 84192
rect 291568 84244 291620 84250
rect 291568 84186 291620 84192
rect 291580 79354 291608 84186
rect 291568 79348 291620 79354
rect 291568 79290 291620 79296
rect 291476 66156 291528 66162
rect 291476 66098 291528 66104
rect 291488 46986 291516 66098
rect 291476 46980 291528 46986
rect 291476 46922 291528 46928
rect 291568 46980 291620 46986
rect 291568 46922 291620 46928
rect 291580 41426 291608 46922
rect 291580 41398 291700 41426
rect 291672 41290 291700 41398
rect 291580 41262 291700 41290
rect 291580 37210 291608 41262
rect 291580 37182 291700 37210
rect 291672 12306 291700 37182
rect 291842 29608 291898 29617
rect 291842 29543 291898 29552
rect 291856 29073 291884 29543
rect 291842 29064 291898 29073
rect 291842 28999 291898 29008
rect 291660 12300 291712 12306
rect 291660 12242 291712 12248
rect 291292 7064 291344 7070
rect 291292 7006 291344 7012
rect 291200 6656 291252 6662
rect 291200 6598 291252 6604
rect 290740 5500 290792 5506
rect 290740 5442 290792 5448
rect 290464 3936 290516 3942
rect 290464 3878 290516 3884
rect 287704 3664 287756 3670
rect 287704 3606 287756 3612
rect 288348 3664 288400 3670
rect 288348 3606 288400 3612
rect 288360 480 288388 3606
rect 289544 3188 289596 3194
rect 289544 3130 289596 3136
rect 289556 480 289584 3130
rect 290752 480 290780 5442
rect 292500 4146 292528 338030
rect 292592 6730 292620 340054
rect 292960 335628 292988 340054
rect 292684 335600 292988 335628
rect 292684 7002 292712 335600
rect 293604 328506 293632 340054
rect 292764 328500 292816 328506
rect 292764 328442 292816 328448
rect 293592 328500 293644 328506
rect 293592 328442 293644 328448
rect 292776 321638 292804 328442
rect 292764 321632 292816 321638
rect 292764 321574 292816 321580
rect 292856 321496 292908 321502
rect 292856 321438 292908 321444
rect 292868 318782 292896 321438
rect 292856 318776 292908 318782
rect 292856 318718 292908 318724
rect 292856 309188 292908 309194
rect 292856 309130 292908 309136
rect 292868 176610 292896 309130
rect 292776 176582 292896 176610
rect 292776 176338 292804 176582
rect 292776 176310 292896 176338
rect 292868 118794 292896 176310
rect 292856 118788 292908 118794
rect 292856 118730 292908 118736
rect 292856 118652 292908 118658
rect 292856 118594 292908 118600
rect 292868 99498 292896 118594
rect 292776 99470 292896 99498
rect 292776 99362 292804 99470
rect 292776 99334 292896 99362
rect 292762 87272 292818 87281
rect 292762 87207 292764 87216
rect 292816 87207 292818 87216
rect 292764 87178 292816 87184
rect 292868 80186 292896 99334
rect 292868 80158 292988 80186
rect 292960 80016 292988 80158
rect 292868 79988 292988 80016
rect 292868 71074 292896 79988
rect 292776 71046 292896 71074
rect 292776 64870 292804 71046
rect 292764 64864 292816 64870
rect 292764 64806 292816 64812
rect 292856 64864 292908 64870
rect 292856 64806 292908 64812
rect 292868 47002 292896 64806
rect 292776 46974 292896 47002
rect 292776 40746 292804 46974
rect 292776 40718 292896 40746
rect 292868 30734 292896 40718
rect 292856 30728 292908 30734
rect 292856 30670 292908 30676
rect 292764 26308 292816 26314
rect 292764 26250 292816 26256
rect 292776 19378 292804 26250
rect 292764 19372 292816 19378
rect 292764 19314 292816 19320
rect 292856 19372 292908 19378
rect 292856 19314 292908 19320
rect 292868 12458 292896 19314
rect 292868 12430 292988 12458
rect 292960 12374 292988 12430
rect 292948 12368 293000 12374
rect 292948 12310 293000 12316
rect 292672 6996 292724 7002
rect 292672 6938 292724 6944
rect 293972 6798 294000 340054
rect 294052 335640 294104 335646
rect 294052 335582 294104 335588
rect 294064 12442 294092 335582
rect 294248 13462 294276 340054
rect 294800 335646 294828 340054
rect 294788 335640 294840 335646
rect 294788 335582 294840 335588
rect 294236 13456 294288 13462
rect 294236 13398 294288 13404
rect 294052 12436 294104 12442
rect 294052 12378 294104 12384
rect 295352 6866 295380 340054
rect 295432 331628 295484 331634
rect 295432 331570 295484 331576
rect 295444 11694 295472 331570
rect 295628 13530 295656 340054
rect 296088 331634 296116 340054
rect 296076 331628 296128 331634
rect 296076 331570 296128 331576
rect 295616 13524 295668 13530
rect 295616 13466 295668 13472
rect 295432 11688 295484 11694
rect 295432 11630 295484 11636
rect 295340 6860 295392 6866
rect 295340 6802 295392 6808
rect 293960 6792 294012 6798
rect 293960 6734 294012 6740
rect 292580 6724 292632 6730
rect 292580 6666 292632 6672
rect 296732 6118 296760 340054
rect 296812 335640 296864 335646
rect 296812 335582 296864 335588
rect 296824 11626 296852 335582
rect 297008 13598 297036 340054
rect 297376 335646 297404 340054
rect 297916 337204 297968 337210
rect 297916 337146 297968 337152
rect 297364 335640 297416 335646
rect 297364 335582 297416 335588
rect 297546 40352 297602 40361
rect 297546 40287 297602 40296
rect 297560 40089 297588 40287
rect 297546 40080 297602 40089
rect 297546 40015 297602 40024
rect 296996 13592 297048 13598
rect 296996 13534 297048 13540
rect 296812 11620 296864 11626
rect 296812 11562 296864 11568
rect 296720 6112 296772 6118
rect 296720 6054 296772 6060
rect 294328 4344 294380 4350
rect 294328 4286 294380 4292
rect 291936 4140 291988 4146
rect 291936 4082 291988 4088
rect 292488 4140 292540 4146
rect 292488 4082 292540 4088
rect 291948 480 291976 4082
rect 293132 3936 293184 3942
rect 293132 3878 293184 3884
rect 293144 480 293172 3878
rect 294340 480 294368 4286
rect 297928 4146 297956 337146
rect 298112 6050 298140 340054
rect 298296 13666 298324 340054
rect 298940 331498 298968 340054
rect 298468 331492 298520 331498
rect 298468 331434 298520 331440
rect 298928 331492 298980 331498
rect 298928 331434 298980 331440
rect 298480 321314 298508 331434
rect 298480 321286 298600 321314
rect 298572 318782 298600 321286
rect 298468 318776 298520 318782
rect 298468 318718 298520 318724
rect 298560 318776 298612 318782
rect 298560 318718 298612 318724
rect 298480 317422 298508 318718
rect 298468 317416 298520 317422
rect 298468 317358 298520 317364
rect 298468 307828 298520 307834
rect 298468 307770 298520 307776
rect 298480 304314 298508 307770
rect 298388 304286 298508 304314
rect 298388 302002 298416 304286
rect 298388 301974 298600 302002
rect 298572 299470 298600 301974
rect 298560 299464 298612 299470
rect 298560 299406 298612 299412
rect 298468 289876 298520 289882
rect 298468 289818 298520 289824
rect 298480 282946 298508 289818
rect 298468 282940 298520 282946
rect 298468 282882 298520 282888
rect 298560 282804 298612 282810
rect 298560 282746 298612 282752
rect 298572 280158 298600 282746
rect 298560 280152 298612 280158
rect 298560 280094 298612 280100
rect 298468 270632 298520 270638
rect 298468 270574 298520 270580
rect 298480 263634 298508 270574
rect 298468 263628 298520 263634
rect 298468 263570 298520 263576
rect 298560 263492 298612 263498
rect 298560 263434 298612 263440
rect 298572 260846 298600 263434
rect 298560 260840 298612 260846
rect 298560 260782 298612 260788
rect 298468 251320 298520 251326
rect 298468 251262 298520 251268
rect 298480 251190 298508 251262
rect 298468 251184 298520 251190
rect 298468 251126 298520 251132
rect 298560 241528 298612 241534
rect 298560 241470 298612 241476
rect 298572 231878 298600 241470
rect 298560 231872 298612 231878
rect 298560 231814 298612 231820
rect 298560 231736 298612 231742
rect 298560 231678 298612 231684
rect 298572 229090 298600 231678
rect 298560 229084 298612 229090
rect 298560 229026 298612 229032
rect 298652 229084 298704 229090
rect 298652 229026 298704 229032
rect 298664 201550 298692 229026
rect 298560 201544 298612 201550
rect 298560 201486 298612 201492
rect 298652 201544 298704 201550
rect 298652 201486 298704 201492
rect 298572 196110 298600 201486
rect 298560 196104 298612 196110
rect 298560 196046 298612 196052
rect 298468 193248 298520 193254
rect 298468 193190 298520 193196
rect 298480 186266 298508 193190
rect 298480 186238 298600 186266
rect 298572 157332 298600 186238
rect 298480 157304 298600 157332
rect 298480 147642 298508 157304
rect 298480 147614 298600 147642
rect 298572 115954 298600 147614
rect 298480 115938 298600 115954
rect 298468 115932 298600 115938
rect 298520 115926 298600 115932
rect 298468 115874 298520 115880
rect 298480 115843 298508 115874
rect 298560 108860 298612 108866
rect 298560 108802 298612 108808
rect 298572 99482 298600 108802
rect 298560 99476 298612 99482
rect 298560 99418 298612 99424
rect 298468 99340 298520 99346
rect 298468 99282 298520 99288
rect 298480 86970 298508 99282
rect 298468 86964 298520 86970
rect 298468 86906 298520 86912
rect 298560 86964 298612 86970
rect 298560 86906 298612 86912
rect 298572 82090 298600 86906
rect 298480 82062 298600 82090
rect 298480 60602 298508 82062
rect 298480 60574 298600 60602
rect 298572 48362 298600 60574
rect 298480 48334 298600 48362
rect 298480 41154 298508 48334
rect 298480 41126 298600 41154
rect 298572 28966 298600 41126
rect 298560 28960 298612 28966
rect 298560 28902 298612 28908
rect 298652 28960 298704 28966
rect 298652 28902 298704 28908
rect 298284 13660 298336 13666
rect 298284 13602 298336 13608
rect 298664 11558 298692 28902
rect 298652 11552 298704 11558
rect 298652 11494 298704 11500
rect 298100 6044 298152 6050
rect 298100 5986 298152 5992
rect 299492 5982 299520 340054
rect 299676 13734 299704 340054
rect 300228 331242 300256 340054
rect 299860 331214 300256 331242
rect 299860 311930 299888 331214
rect 299768 311902 299888 311930
rect 299768 311794 299796 311902
rect 299768 311766 299888 311794
rect 299860 292618 299888 311766
rect 299768 292590 299888 292618
rect 299768 292482 299796 292590
rect 299768 292454 299888 292482
rect 299860 273222 299888 292454
rect 299848 273216 299900 273222
rect 299848 273158 299900 273164
rect 299848 273080 299900 273086
rect 299848 273022 299900 273028
rect 299860 253910 299888 273022
rect 299848 253904 299900 253910
rect 299848 253846 299900 253852
rect 299848 253768 299900 253774
rect 299848 253710 299900 253716
rect 299860 234598 299888 253710
rect 299848 234592 299900 234598
rect 299848 234534 299900 234540
rect 299848 234456 299900 234462
rect 299848 234398 299900 234404
rect 299860 215286 299888 234398
rect 299848 215280 299900 215286
rect 299848 215222 299900 215228
rect 299848 215144 299900 215150
rect 299848 215086 299900 215092
rect 299860 195974 299888 215086
rect 299848 195968 299900 195974
rect 299848 195910 299900 195916
rect 299848 195832 299900 195838
rect 299848 195774 299900 195780
rect 299860 174010 299888 195774
rect 299848 174004 299900 174010
rect 299848 173946 299900 173952
rect 299756 173936 299808 173942
rect 299756 173878 299808 173884
rect 299768 172514 299796 173878
rect 299756 172508 299808 172514
rect 299756 172450 299808 172456
rect 300032 172508 300084 172514
rect 300032 172450 300084 172456
rect 300044 157026 300072 172450
rect 299860 156998 300072 157026
rect 299860 118810 299888 156998
rect 299768 118782 299888 118810
rect 299768 118674 299796 118782
rect 299768 118646 299888 118674
rect 299860 80102 299888 118646
rect 299848 80096 299900 80102
rect 299848 80038 299900 80044
rect 299848 79960 299900 79966
rect 299848 79902 299900 79908
rect 299860 51202 299888 79902
rect 299848 51196 299900 51202
rect 299848 51138 299900 51144
rect 299848 48340 299900 48346
rect 299848 48282 299900 48288
rect 299860 45558 299888 48282
rect 299848 45552 299900 45558
rect 299848 45494 299900 45500
rect 299940 45552 299992 45558
rect 299940 45494 299992 45500
rect 299952 36009 299980 45494
rect 299754 36000 299810 36009
rect 299754 35935 299810 35944
rect 299938 36000 299994 36009
rect 299938 35935 299994 35944
rect 299768 35902 299796 35935
rect 299756 35896 299808 35902
rect 299756 35838 299808 35844
rect 300032 35896 300084 35902
rect 300032 35838 300084 35844
rect 300044 16726 300072 35838
rect 300032 16720 300084 16726
rect 300032 16662 300084 16668
rect 299848 15224 299900 15230
rect 299848 15166 299900 15172
rect 299664 13728 299716 13734
rect 299664 13670 299716 13676
rect 299860 11490 299888 15166
rect 299848 11484 299900 11490
rect 299848 11426 299900 11432
rect 299480 5976 299532 5982
rect 299480 5918 299532 5924
rect 300872 5914 300900 340068
rect 301056 340054 301346 340082
rect 301424 340054 301806 340082
rect 300952 332852 301004 332858
rect 300952 332794 301004 332800
rect 300964 11422 300992 332794
rect 301056 13802 301084 340054
rect 301424 332858 301452 340054
rect 301412 332852 301464 332858
rect 301412 332794 301464 332800
rect 301044 13796 301096 13802
rect 301044 13738 301096 13744
rect 300952 11416 301004 11422
rect 300952 11358 301004 11364
rect 300860 5908 300912 5914
rect 300860 5850 300912 5856
rect 302252 5846 302280 340068
rect 302436 340054 302726 340082
rect 302896 340054 303186 340082
rect 302332 335640 302384 335646
rect 302332 335582 302384 335588
rect 302344 11354 302372 335582
rect 302436 13054 302464 340054
rect 302896 335646 302924 340054
rect 303528 337340 303580 337346
rect 303528 337282 303580 337288
rect 302884 335640 302936 335646
rect 302884 335582 302936 335588
rect 302424 13048 302476 13054
rect 302424 12990 302476 12996
rect 302332 11348 302384 11354
rect 302332 11290 302384 11296
rect 302240 5840 302292 5846
rect 302240 5782 302292 5788
rect 298008 4276 298060 4282
rect 298008 4218 298060 4224
rect 296720 4140 296772 4146
rect 296720 4082 296772 4088
rect 297916 4140 297968 4146
rect 297916 4082 297968 4088
rect 295524 3120 295576 3126
rect 295524 3062 295576 3068
rect 295536 480 295564 3062
rect 296732 480 296760 4082
rect 298020 2122 298048 4218
rect 301412 4208 301464 4214
rect 301412 4150 301464 4156
rect 299112 3324 299164 3330
rect 299112 3266 299164 3272
rect 297928 2094 298048 2122
rect 297928 480 297956 2094
rect 299124 480 299152 3266
rect 300308 3052 300360 3058
rect 300308 2994 300360 3000
rect 300320 480 300348 2994
rect 301424 480 301452 4150
rect 303540 2922 303568 337282
rect 303632 5778 303660 340068
rect 303908 340054 304106 340082
rect 304184 340054 304566 340082
rect 304644 340054 304934 340082
rect 305104 340054 305394 340082
rect 303712 335708 303764 335714
rect 303712 335650 303764 335656
rect 303620 5772 303672 5778
rect 303620 5714 303672 5720
rect 303724 5710 303752 335650
rect 303804 335640 303856 335646
rect 303804 335582 303856 335588
rect 303816 11286 303844 335582
rect 303908 14074 303936 340054
rect 304184 335646 304212 340054
rect 304644 335714 304672 340054
rect 304632 335708 304684 335714
rect 304632 335650 304684 335656
rect 304172 335640 304224 335646
rect 304172 335582 304224 335588
rect 305000 118788 305052 118794
rect 305000 118730 305052 118736
rect 305012 113257 305040 118730
rect 304998 113248 305054 113257
rect 304998 113183 305054 113192
rect 305104 103630 305132 340054
rect 305840 337278 305868 340068
rect 306116 340054 306314 340082
rect 306576 340054 306774 340082
rect 306944 340054 307234 340082
rect 307312 340054 307694 340082
rect 307864 340054 308154 340082
rect 308232 340054 308522 340082
rect 308692 340054 308982 340082
rect 309244 340054 309442 340082
rect 309520 340054 309902 340082
rect 310164 340054 310362 340082
rect 310624 340054 310822 340082
rect 310992 340054 311282 340082
rect 311452 340054 311742 340082
rect 312004 340054 312110 340082
rect 312280 340054 312570 340082
rect 312648 340054 313030 340082
rect 305828 337272 305880 337278
rect 305828 337214 305880 337220
rect 306116 328506 306144 340054
rect 306472 335708 306524 335714
rect 306472 335650 306524 335656
rect 306380 335640 306432 335646
rect 306380 335582 306432 335588
rect 305368 328500 305420 328506
rect 305368 328442 305420 328448
rect 306104 328500 306156 328506
rect 306104 328442 306156 328448
rect 305380 312798 305408 328442
rect 305368 312792 305420 312798
rect 305368 312734 305420 312740
rect 305644 312792 305696 312798
rect 305644 312734 305696 312740
rect 305656 307850 305684 312734
rect 305564 307822 305684 307850
rect 305564 307766 305592 307822
rect 305552 307760 305604 307766
rect 305552 307702 305604 307708
rect 305460 298172 305512 298178
rect 305460 298114 305512 298120
rect 305472 289882 305500 298114
rect 305460 289876 305512 289882
rect 305460 289818 305512 289824
rect 305460 289740 305512 289746
rect 305460 289682 305512 289688
rect 305472 280158 305500 289682
rect 305460 280152 305512 280158
rect 305460 280094 305512 280100
rect 305276 280084 305328 280090
rect 305276 280026 305328 280032
rect 305288 278769 305316 280026
rect 305274 278760 305330 278769
rect 305274 278695 305330 278704
rect 305550 278760 305606 278769
rect 305550 278695 305606 278704
rect 305564 253722 305592 278695
rect 305288 253694 305592 253722
rect 305288 251190 305316 253694
rect 305276 251184 305328 251190
rect 305276 251126 305328 251132
rect 305184 241528 305236 241534
rect 305184 241470 305236 241476
rect 305196 231878 305224 241470
rect 305184 231872 305236 231878
rect 305184 231814 305236 231820
rect 305276 231872 305328 231878
rect 305276 231814 305328 231820
rect 305288 220810 305316 231814
rect 305288 220782 305408 220810
rect 305380 215354 305408 220782
rect 305368 215348 305420 215354
rect 305368 215290 305420 215296
rect 305276 215280 305328 215286
rect 305276 215222 305328 215228
rect 305288 205698 305316 215222
rect 305276 205692 305328 205698
rect 305276 205634 305328 205640
rect 305276 202904 305328 202910
rect 305276 202846 305328 202852
rect 305288 201482 305316 202846
rect 305276 201476 305328 201482
rect 305276 201418 305328 201424
rect 305276 195968 305328 195974
rect 305276 195910 305328 195916
rect 305288 188442 305316 195910
rect 305196 188414 305316 188442
rect 305196 183598 305224 188414
rect 305184 183592 305236 183598
rect 305184 183534 305236 183540
rect 305460 183592 305512 183598
rect 305460 183534 305512 183540
rect 305472 173942 305500 183534
rect 305368 173936 305420 173942
rect 305368 173878 305420 173884
rect 305460 173936 305512 173942
rect 305460 173878 305512 173884
rect 305380 162858 305408 173878
rect 305368 162852 305420 162858
rect 305368 162794 305420 162800
rect 305276 153264 305328 153270
rect 305276 153206 305328 153212
rect 305288 153134 305316 153206
rect 305276 153128 305328 153134
rect 305276 153070 305328 153076
rect 305368 142180 305420 142186
rect 305368 142122 305420 142128
rect 305380 132462 305408 142122
rect 305368 132456 305420 132462
rect 305368 132398 305420 132404
rect 305368 122868 305420 122874
rect 305368 122810 305420 122816
rect 305380 118794 305408 122810
rect 305368 118788 305420 118794
rect 305368 118730 305420 118736
rect 305274 113248 305330 113257
rect 305274 113183 305330 113192
rect 305288 106282 305316 113183
rect 305276 106276 305328 106282
rect 305276 106218 305328 106224
rect 305092 103624 305144 103630
rect 305092 103566 305144 103572
rect 305092 103488 305144 103494
rect 305092 103430 305144 103436
rect 303896 14068 303948 14074
rect 303896 14010 303948 14016
rect 303804 11280 303856 11286
rect 303804 11222 303856 11228
rect 305104 9586 305132 103430
rect 305276 102196 305328 102202
rect 305276 102138 305328 102144
rect 305288 97322 305316 102138
rect 305288 97294 305592 97322
rect 305564 87038 305592 97294
rect 305552 87032 305604 87038
rect 305552 86974 305604 86980
rect 305460 86964 305512 86970
rect 305460 86906 305512 86912
rect 305472 74594 305500 86906
rect 305276 74588 305328 74594
rect 305276 74530 305328 74536
rect 305460 74588 305512 74594
rect 305460 74530 305512 74536
rect 305288 74458 305316 74530
rect 305276 74452 305328 74458
rect 305276 74394 305328 74400
rect 305368 64932 305420 64938
rect 305368 64874 305420 64880
rect 305380 53122 305408 64874
rect 305380 53094 305500 53122
rect 305472 40746 305500 53094
rect 305380 40718 305500 40746
rect 305380 35902 305408 40718
rect 305368 35896 305420 35902
rect 305368 35838 305420 35844
rect 306286 29472 306342 29481
rect 306286 29407 306342 29416
rect 306300 29209 306328 29407
rect 306286 29200 306342 29209
rect 306286 29135 306342 29144
rect 305368 24880 305420 24886
rect 305368 24822 305420 24828
rect 305380 15201 305408 24822
rect 305182 15192 305238 15201
rect 305182 15127 305238 15136
rect 305366 15192 305422 15201
rect 305366 15127 305422 15136
rect 305092 9580 305144 9586
rect 305092 9522 305144 9528
rect 305000 6452 305052 6458
rect 305000 6394 305052 6400
rect 303712 5704 303764 5710
rect 303712 5646 303764 5652
rect 303804 2984 303856 2990
rect 303804 2926 303856 2932
rect 302608 2916 302660 2922
rect 302608 2858 302660 2864
rect 303528 2916 303580 2922
rect 303528 2858 303580 2864
rect 302620 480 302648 2858
rect 303816 480 303844 2926
rect 305012 480 305040 6394
rect 305196 5642 305224 15127
rect 305184 5636 305236 5642
rect 305184 5578 305236 5584
rect 306392 4865 306420 335582
rect 306484 5574 306512 335650
rect 306576 9654 306604 340054
rect 306944 335646 306972 340054
rect 307312 335714 307340 340054
rect 307300 335708 307352 335714
rect 307300 335650 307352 335656
rect 306932 335640 306984 335646
rect 306932 335582 306984 335588
rect 307760 335640 307812 335646
rect 307760 335582 307812 335588
rect 306564 9648 306616 9654
rect 306564 9590 306616 9596
rect 306472 5568 306524 5574
rect 306472 5510 306524 5516
rect 306378 4856 306434 4865
rect 306378 4791 306434 4800
rect 307772 4690 307800 335582
rect 307864 8906 307892 340054
rect 308232 335646 308260 340054
rect 308220 335640 308272 335646
rect 308220 335582 308272 335588
rect 308692 328506 308720 340054
rect 309140 335640 309192 335646
rect 309140 335582 309192 335588
rect 308128 328500 308180 328506
rect 308128 328442 308180 328448
rect 308680 328500 308732 328506
rect 308680 328442 308732 328448
rect 308140 311930 308168 328442
rect 308048 311902 308168 311930
rect 308048 309126 308076 311902
rect 308036 309120 308088 309126
rect 308036 309062 308088 309068
rect 308220 309120 308272 309126
rect 308220 309062 308272 309068
rect 308232 302954 308260 309062
rect 308140 302926 308260 302954
rect 308140 298110 308168 302926
rect 308128 298104 308180 298110
rect 308128 298046 308180 298052
rect 308220 298104 308272 298110
rect 308220 298046 308272 298052
rect 308232 278798 308260 298046
rect 307944 278792 307996 278798
rect 307944 278734 307996 278740
rect 308220 278792 308272 278798
rect 308220 278734 308272 278740
rect 307956 270502 307984 278734
rect 307944 270496 307996 270502
rect 307944 270438 307996 270444
rect 307944 258120 307996 258126
rect 307944 258062 307996 258068
rect 307956 251190 307984 258062
rect 307944 251184 307996 251190
rect 307944 251126 307996 251132
rect 308036 244248 308088 244254
rect 308036 244190 308088 244196
rect 308048 232014 308076 244190
rect 308036 232008 308088 232014
rect 308036 231950 308088 231956
rect 308036 231872 308088 231878
rect 308036 231814 308088 231820
rect 308048 217462 308076 231814
rect 308036 217456 308088 217462
rect 308036 217398 308088 217404
rect 308036 212560 308088 212566
rect 308034 212528 308036 212537
rect 308088 212528 308090 212537
rect 308034 212463 308090 212472
rect 308218 212528 308274 212537
rect 308218 212463 308274 212472
rect 308232 205562 308260 212463
rect 308036 205556 308088 205562
rect 308036 205498 308088 205504
rect 308220 205556 308272 205562
rect 308220 205498 308272 205504
rect 308048 196042 308076 205498
rect 308036 196036 308088 196042
rect 308036 195978 308088 195984
rect 308036 193248 308088 193254
rect 308034 193216 308036 193225
rect 308088 193216 308090 193225
rect 308034 193151 308090 193160
rect 308310 193216 308366 193225
rect 308310 193151 308366 193160
rect 308324 183598 308352 193151
rect 308128 183592 308180 183598
rect 308128 183534 308180 183540
rect 308312 183592 308364 183598
rect 308312 183534 308364 183540
rect 308140 178786 308168 183534
rect 309046 181112 309102 181121
rect 309046 181047 309048 181056
rect 309100 181047 309102 181056
rect 309048 181018 309100 181024
rect 308140 178758 308260 178786
rect 308232 173942 308260 178758
rect 308036 173936 308088 173942
rect 308036 173878 308088 173884
rect 308220 173936 308272 173942
rect 308220 173878 308272 173884
rect 308048 162874 308076 173878
rect 308048 162846 308168 162874
rect 308140 161430 308168 162846
rect 308128 161424 308180 161430
rect 308128 161366 308180 161372
rect 308036 151836 308088 151842
rect 308036 151778 308088 151784
rect 308048 148322 308076 151778
rect 308048 148294 308260 148322
rect 308232 133958 308260 148294
rect 309046 134056 309102 134065
rect 309046 133991 309102 134000
rect 308128 133952 308180 133958
rect 308128 133894 308180 133900
rect 308220 133952 308272 133958
rect 308220 133894 308272 133900
rect 308140 124250 308168 133894
rect 309060 133793 309088 133991
rect 309046 133784 309102 133793
rect 309046 133719 309102 133728
rect 308048 124222 308168 124250
rect 308048 108338 308076 124222
rect 308048 108310 308260 108338
rect 308232 104802 308260 108310
rect 308140 104774 308260 104802
rect 308140 103494 308168 104774
rect 308036 103488 308088 103494
rect 308036 103430 308088 103436
rect 308128 103488 308180 103494
rect 308128 103430 308180 103436
rect 308048 98546 308076 103430
rect 308048 98518 308168 98546
rect 308140 87009 308168 98518
rect 307942 87000 307998 87009
rect 307942 86935 307998 86944
rect 308126 87000 308182 87009
rect 308126 86935 308182 86944
rect 307956 84182 307984 86935
rect 307944 84176 307996 84182
rect 307944 84118 307996 84124
rect 308128 74588 308180 74594
rect 308128 74530 308180 74536
rect 308140 74474 308168 74530
rect 308048 74446 308168 74474
rect 308048 66298 308076 74446
rect 308036 66292 308088 66298
rect 308036 66234 308088 66240
rect 308036 64932 308088 64938
rect 308036 64874 308088 64880
rect 308048 64818 308076 64874
rect 308048 64790 308260 64818
rect 308232 56522 308260 64790
rect 308140 56494 308260 56522
rect 308140 50402 308168 56494
rect 308140 50374 308260 50402
rect 308232 44169 308260 50374
rect 307942 44160 307998 44169
rect 307942 44095 307998 44104
rect 308218 44160 308274 44169
rect 308218 44095 308274 44104
rect 307956 34542 307984 44095
rect 307944 34536 307996 34542
rect 307944 34478 307996 34484
rect 308128 34536 308180 34542
rect 308128 34478 308180 34484
rect 308140 19514 308168 34478
rect 308128 19508 308180 19514
rect 308128 19450 308180 19456
rect 307852 8900 307904 8906
rect 307852 8842 307904 8848
rect 309152 4706 309180 335582
rect 309244 8838 309272 340054
rect 309520 335646 309548 340054
rect 309508 335640 309560 335646
rect 309508 335582 309560 335588
rect 310164 328545 310192 340054
rect 310520 335640 310572 335646
rect 310520 335582 310572 335588
rect 310150 328536 310206 328545
rect 310150 328471 310206 328480
rect 309414 328400 309470 328409
rect 309414 328335 309470 328344
rect 309428 273222 309456 328335
rect 309416 273216 309468 273222
rect 309416 273158 309468 273164
rect 309416 267776 309468 267782
rect 309416 267718 309468 267724
rect 309428 253994 309456 267718
rect 309336 253966 309456 253994
rect 309336 253858 309364 253966
rect 309336 253830 309456 253858
rect 309428 215370 309456 253830
rect 309336 215342 309456 215370
rect 309336 215234 309364 215342
rect 309336 215206 309456 215234
rect 309428 205714 309456 215206
rect 309428 205686 309548 205714
rect 309520 201521 309548 205686
rect 309322 201512 309378 201521
rect 309322 201447 309324 201456
rect 309376 201447 309378 201456
rect 309506 201512 309562 201521
rect 309506 201447 309562 201456
rect 309324 201418 309376 201424
rect 309416 201408 309468 201414
rect 309416 201350 309468 201356
rect 309428 176746 309456 201350
rect 310428 185632 310480 185638
rect 310428 185574 310480 185580
rect 310440 180849 310468 185574
rect 310426 180840 310482 180849
rect 310426 180775 310482 180784
rect 309336 176718 309456 176746
rect 309336 176610 309364 176718
rect 309336 176582 309456 176610
rect 309428 150362 309456 176582
rect 309428 150334 309548 150362
rect 309520 149054 309548 150334
rect 309508 149048 309560 149054
rect 309508 148990 309560 148996
rect 309508 139460 309560 139466
rect 309508 139402 309560 139408
rect 309520 134570 309548 139402
rect 309508 134564 309560 134570
rect 309508 134506 309560 134512
rect 309692 134564 309744 134570
rect 309692 134506 309744 134512
rect 309704 120154 309732 134506
rect 309416 120148 309468 120154
rect 309416 120090 309468 120096
rect 309692 120148 309744 120154
rect 309692 120090 309744 120096
rect 309428 120034 309456 120090
rect 309336 120006 309456 120034
rect 309336 115258 309364 120006
rect 309324 115252 309376 115258
rect 309324 115194 309376 115200
rect 309324 102468 309376 102474
rect 309324 102410 309376 102416
rect 309336 97322 309364 102410
rect 309336 97294 309456 97322
rect 309428 89826 309456 97294
rect 309416 89820 309468 89826
rect 309416 89762 309468 89768
rect 309416 85604 309468 85610
rect 309416 85546 309468 85552
rect 309428 80186 309456 85546
rect 309428 80158 309548 80186
rect 309520 75868 309548 80158
rect 309336 75840 309548 75868
rect 309336 66230 309364 75840
rect 309324 66224 309376 66230
rect 309324 66166 309376 66172
rect 309416 66224 309468 66230
rect 309416 66166 309468 66172
rect 309428 56642 309456 66166
rect 309416 56636 309468 56642
rect 309416 56578 309468 56584
rect 309508 56500 309560 56506
rect 309508 56442 309560 56448
rect 309520 30954 309548 56442
rect 309336 30926 309548 30954
rect 309336 12918 309364 30926
rect 309324 12912 309376 12918
rect 309324 12854 309376 12860
rect 309232 8832 309284 8838
rect 309232 8774 309284 8780
rect 310532 4842 310560 335582
rect 310624 8770 310652 340054
rect 310992 335646 311020 340054
rect 310980 335640 311032 335646
rect 310980 335582 311032 335588
rect 311452 328506 311480 340054
rect 311900 335776 311952 335782
rect 311900 335718 311952 335724
rect 310888 328500 310940 328506
rect 310888 328442 310940 328448
rect 311440 328500 311492 328506
rect 311440 328442 311492 328448
rect 310900 318594 310928 328442
rect 310808 318566 310928 318594
rect 310808 316033 310836 318566
rect 310794 316024 310850 316033
rect 310794 315959 310850 315968
rect 310886 315888 310942 315897
rect 310886 315823 310942 315832
rect 310900 298178 310928 315823
rect 310888 298172 310940 298178
rect 310888 298114 310940 298120
rect 310796 296744 310848 296750
rect 310796 296686 310848 296692
rect 310808 295798 310836 296686
rect 310796 295792 310848 295798
rect 310796 295734 310848 295740
rect 310980 295792 311032 295798
rect 310980 295734 311032 295740
rect 310992 287042 311020 295734
rect 310808 287014 311020 287042
rect 310808 277438 310836 287014
rect 310704 277432 310756 277438
rect 310704 277374 310756 277380
rect 310796 277432 310848 277438
rect 310796 277374 310848 277380
rect 310716 273426 310744 277374
rect 310704 273420 310756 273426
rect 310704 273362 310756 273368
rect 310796 267844 310848 267850
rect 310796 267786 310848 267792
rect 310808 263702 310836 267786
rect 310796 263696 310848 263702
rect 310796 263638 310848 263644
rect 310796 263560 310848 263566
rect 310796 263502 310848 263508
rect 310808 258074 310836 263502
rect 310808 258046 310928 258074
rect 310900 256698 310928 258046
rect 310888 256692 310940 256698
rect 310888 256634 310940 256640
rect 310796 240032 310848 240038
rect 310796 239974 310848 239980
rect 310808 238746 310836 239974
rect 310704 238740 310756 238746
rect 310704 238682 310756 238688
rect 310796 238740 310848 238746
rect 310796 238682 310848 238688
rect 310716 229129 310744 238682
rect 310702 229120 310758 229129
rect 310702 229055 310758 229064
rect 310978 229120 311034 229129
rect 310978 229055 311034 229064
rect 310992 227066 311020 229055
rect 310900 227038 311020 227066
rect 310900 219434 310928 227038
rect 310888 219428 310940 219434
rect 310888 219370 310940 219376
rect 310888 214600 310940 214606
rect 310888 214542 310940 214548
rect 310900 201482 310928 214542
rect 310796 201476 310848 201482
rect 310796 201418 310848 201424
rect 310888 201476 310940 201482
rect 310888 201418 310940 201424
rect 310808 200122 310836 201418
rect 310796 200116 310848 200122
rect 310796 200058 310848 200064
rect 310794 180840 310850 180849
rect 310794 180775 310850 180784
rect 310808 179382 310836 180775
rect 310796 179376 310848 179382
rect 310796 179318 310848 179324
rect 310888 169788 310940 169794
rect 310888 169730 310940 169736
rect 310900 161430 310928 169730
rect 310888 161424 310940 161430
rect 310888 161366 310940 161372
rect 310980 161424 311032 161430
rect 310980 161366 311032 161372
rect 310992 149546 311020 161366
rect 310900 149518 311020 149546
rect 310900 133906 310928 149518
rect 310808 133890 310928 133906
rect 310796 133884 310928 133890
rect 310848 133878 310928 133884
rect 310796 133826 310848 133832
rect 310808 133795 310836 133826
rect 310796 124228 310848 124234
rect 310796 124170 310848 124176
rect 310808 114646 310836 124170
rect 310796 114640 310848 114646
rect 310796 114582 310848 114588
rect 310888 114504 310940 114510
rect 310888 114446 310940 114452
rect 310900 103494 310928 114446
rect 310888 103488 310940 103494
rect 310888 103430 310940 103436
rect 311072 103488 311124 103494
rect 311072 103430 311124 103436
rect 311084 93945 311112 103430
rect 311070 93936 311126 93945
rect 311070 93871 311126 93880
rect 310978 93800 311034 93809
rect 310978 93735 311034 93744
rect 310992 74474 311020 93735
rect 310900 74446 311020 74474
rect 310900 64938 310928 74446
rect 310888 64932 310940 64938
rect 310888 64874 310940 64880
rect 310980 64932 311032 64938
rect 310980 64874 311032 64880
rect 310992 58818 311020 64874
rect 310796 58812 310848 58818
rect 310796 58754 310848 58760
rect 310980 58812 311032 58818
rect 310980 58754 311032 58760
rect 310808 51762 310836 58754
rect 310808 51734 311020 51762
rect 310992 37346 311020 51734
rect 310808 37318 311020 37346
rect 310808 18086 310836 37318
rect 310796 18080 310848 18086
rect 310796 18022 310848 18028
rect 310704 18012 310756 18018
rect 310704 17954 310756 17960
rect 310716 12850 310744 17954
rect 310704 12844 310756 12850
rect 310704 12786 310756 12792
rect 310612 8764 310664 8770
rect 310612 8706 310664 8712
rect 310532 4814 310652 4842
rect 307760 4684 307812 4690
rect 307760 4626 307812 4632
rect 309060 4678 309180 4706
rect 310520 4684 310572 4690
rect 309060 4622 309088 4678
rect 310520 4626 310572 4632
rect 309048 4616 309100 4622
rect 309048 4558 309100 4564
rect 309140 4616 309192 4622
rect 309140 4558 309192 4564
rect 307392 4140 307444 4146
rect 307392 4082 307444 4088
rect 306196 3256 306248 3262
rect 306196 3198 306248 3204
rect 306208 480 306236 3198
rect 307404 480 307432 4082
rect 309152 2922 309180 4558
rect 310532 3602 310560 4626
rect 310624 4486 310652 4814
rect 311912 4570 311940 335718
rect 312004 8702 312032 340054
rect 312280 335782 312308 340054
rect 312268 335776 312320 335782
rect 312268 335718 312320 335724
rect 312648 334354 312676 340054
rect 313476 338042 313504 340068
rect 313384 338014 313504 338042
rect 313568 340054 313950 340082
rect 314028 340054 314410 340082
rect 314764 340054 314870 340082
rect 315040 340054 315330 340082
rect 315408 340054 315790 340082
rect 312728 337204 312780 337210
rect 312728 337146 312780 337152
rect 312176 334348 312228 334354
rect 312176 334290 312228 334296
rect 312636 334348 312688 334354
rect 312636 334290 312688 334296
rect 312082 181112 312138 181121
rect 312082 181047 312084 181056
rect 312136 181047 312138 181056
rect 312084 181018 312136 181024
rect 312188 12782 312216 334290
rect 312740 334234 312768 337146
rect 313280 335640 313332 335646
rect 313280 335582 313332 335588
rect 312556 334206 312768 334234
rect 312176 12776 312228 12782
rect 312176 12718 312228 12724
rect 311992 8696 312044 8702
rect 311992 8638 312044 8644
rect 311820 4554 311940 4570
rect 311808 4548 311940 4554
rect 311860 4542 311940 4548
rect 311808 4490 311860 4496
rect 310612 4480 310664 4486
rect 310612 4422 310664 4428
rect 310520 3596 310572 3602
rect 310520 3538 310572 3544
rect 312176 3596 312228 3602
rect 312176 3538 312228 3544
rect 309784 3324 309836 3330
rect 309784 3266 309836 3272
rect 309140 2916 309192 2922
rect 309140 2858 309192 2864
rect 308588 2848 308640 2854
rect 308588 2790 308640 2796
rect 308600 480 308628 2790
rect 309796 480 309824 3266
rect 310980 2916 311032 2922
rect 310980 2858 311032 2864
rect 310992 480 311020 2858
rect 312188 480 312216 3538
rect 312556 3126 312584 334206
rect 313188 4480 313240 4486
rect 313188 4422 313240 4428
rect 313200 3806 313228 4422
rect 313292 4418 313320 335582
rect 313384 8634 313412 338014
rect 313568 335646 313596 340054
rect 313556 335640 313608 335646
rect 313556 335582 313608 335588
rect 314028 328545 314056 340054
rect 314660 335300 314712 335306
rect 314660 335242 314712 335248
rect 314014 328536 314070 328545
rect 314014 328471 314070 328480
rect 313738 328400 313794 328409
rect 313738 328335 313794 328344
rect 313752 322266 313780 328335
rect 313660 322238 313780 322266
rect 313660 316033 313688 322238
rect 313462 316024 313518 316033
rect 313462 315959 313518 315968
rect 313646 316024 313702 316033
rect 313646 315959 313702 315968
rect 313476 306406 313504 315959
rect 313464 306400 313516 306406
rect 313464 306342 313516 306348
rect 313556 306400 313608 306406
rect 313556 306342 313608 306348
rect 313568 288538 313596 306342
rect 313568 288510 313688 288538
rect 313660 201482 313688 288510
rect 313556 201476 313608 201482
rect 313556 201418 313608 201424
rect 313648 201476 313700 201482
rect 313648 201418 313700 201424
rect 313568 190482 313596 201418
rect 313568 190454 313688 190482
rect 313660 180810 313688 190454
rect 313648 180804 313700 180810
rect 313648 180746 313700 180752
rect 313740 180804 313792 180810
rect 313740 180746 313792 180752
rect 313752 171170 313780 180746
rect 313568 171142 313780 171170
rect 313568 171086 313596 171142
rect 313556 171080 313608 171086
rect 313556 171022 313608 171028
rect 313832 161492 313884 161498
rect 313832 161434 313884 161440
rect 313844 150618 313872 161434
rect 313832 150612 313884 150618
rect 313832 150554 313884 150560
rect 313648 150476 313700 150482
rect 313648 150418 313700 150424
rect 313660 113150 313688 150418
rect 313648 113144 313700 113150
rect 313648 113086 313700 113092
rect 313464 102468 313516 102474
rect 313464 102410 313516 102416
rect 313476 85610 313504 102410
rect 313464 85604 313516 85610
rect 313464 85546 313516 85552
rect 313648 85604 313700 85610
rect 313648 85546 313700 85552
rect 313660 84182 313688 85546
rect 313648 84176 313700 84182
rect 313648 84118 313700 84124
rect 313740 74588 313792 74594
rect 313740 74530 313792 74536
rect 313752 56710 313780 74530
rect 313740 56704 313792 56710
rect 313740 56646 313792 56652
rect 313740 56568 313792 56574
rect 313740 56510 313792 56516
rect 313752 41478 313780 56510
rect 313556 41472 313608 41478
rect 313556 41414 313608 41420
rect 313740 41472 313792 41478
rect 313740 41414 313792 41420
rect 313568 12714 313596 41414
rect 313556 12708 313608 12714
rect 313556 12650 313608 12656
rect 313372 8628 313424 8634
rect 313372 8570 313424 8576
rect 314672 4758 314700 335242
rect 314764 8566 314792 340054
rect 315040 335306 315068 340054
rect 315028 335300 315080 335306
rect 315028 335242 315080 335248
rect 315408 330274 315436 340054
rect 316040 331016 316092 331022
rect 316040 330958 316092 330964
rect 314936 330268 314988 330274
rect 314936 330210 314988 330216
rect 315396 330268 315448 330274
rect 315396 330210 315448 330216
rect 314948 12646 314976 330210
rect 315946 29200 316002 29209
rect 315946 29135 316002 29144
rect 315960 29073 315988 29135
rect 315946 29064 316002 29073
rect 315946 28999 316002 29008
rect 314936 12640 314988 12646
rect 314936 12582 314988 12588
rect 314752 8560 314804 8566
rect 314752 8502 314804 8508
rect 316052 4826 316080 330958
rect 316144 8498 316172 340068
rect 316328 340054 316618 340082
rect 316696 340054 317078 340082
rect 316328 331022 316356 340054
rect 316696 333418 316724 340054
rect 316776 336932 316828 336938
rect 316776 336874 316828 336880
rect 316604 333390 316724 333418
rect 316316 331016 316368 331022
rect 316316 330958 316368 330964
rect 316604 328506 316632 333390
rect 316788 333282 316816 336874
rect 317420 335708 317472 335714
rect 317420 335650 317472 335656
rect 316696 333254 316816 333282
rect 316408 328500 316460 328506
rect 316408 328442 316460 328448
rect 316592 328500 316644 328506
rect 316592 328442 316644 328448
rect 316420 318918 316448 328442
rect 316408 318912 316460 318918
rect 316408 318854 316460 318860
rect 316316 318776 316368 318782
rect 316316 318718 316368 318724
rect 316328 307766 316356 318718
rect 316316 307760 316368 307766
rect 316316 307702 316368 307708
rect 316316 298172 316368 298178
rect 316316 298114 316368 298120
rect 316328 288522 316356 298114
rect 316316 288516 316368 288522
rect 316316 288458 316368 288464
rect 316224 287088 316276 287094
rect 316224 287030 316276 287036
rect 316236 278798 316264 287030
rect 316224 278792 316276 278798
rect 316224 278734 316276 278740
rect 316316 278792 316368 278798
rect 316316 278734 316368 278740
rect 316328 230466 316356 278734
rect 316236 230438 316356 230466
rect 316236 220862 316264 230438
rect 316224 220856 316276 220862
rect 316224 220798 316276 220804
rect 316316 220856 316368 220862
rect 316316 220798 316368 220804
rect 316328 211138 316356 220798
rect 316316 211132 316368 211138
rect 316316 211074 316368 211080
rect 316500 211132 316552 211138
rect 316500 211074 316552 211080
rect 316512 201521 316540 211074
rect 316314 201512 316370 201521
rect 316314 201447 316370 201456
rect 316498 201512 316554 201521
rect 316498 201447 316554 201456
rect 316328 191894 316356 201447
rect 316316 191888 316368 191894
rect 316316 191830 316368 191836
rect 316224 190528 316276 190534
rect 316224 190470 316276 190476
rect 316236 182238 316264 190470
rect 316224 182232 316276 182238
rect 316224 182174 316276 182180
rect 316316 182232 316368 182238
rect 316316 182174 316368 182180
rect 316328 154562 316356 182174
rect 316316 154556 316368 154562
rect 316316 154498 316368 154504
rect 316408 154556 316460 154562
rect 316408 154498 316460 154504
rect 316420 143562 316448 154498
rect 316328 143534 316448 143562
rect 316328 142118 316356 143534
rect 316316 142112 316368 142118
rect 316316 142054 316368 142060
rect 316316 132524 316368 132530
rect 316316 132466 316368 132472
rect 316328 124302 316356 132466
rect 316316 124296 316368 124302
rect 316316 124238 316368 124244
rect 316224 124228 316276 124234
rect 316224 124170 316276 124176
rect 316236 114578 316264 124170
rect 316224 114572 316276 114578
rect 316224 114514 316276 114520
rect 316316 114572 316368 114578
rect 316316 114514 316368 114520
rect 316328 20618 316356 114514
rect 316236 20590 316356 20618
rect 316236 12578 316264 20590
rect 316224 12572 316276 12578
rect 316224 12514 316276 12520
rect 316132 8492 316184 8498
rect 316132 8434 316184 8440
rect 316696 4978 316724 333254
rect 316604 4950 316724 4978
rect 316040 4820 316092 4826
rect 316040 4762 316092 4768
rect 314660 4752 314712 4758
rect 314660 4694 314712 4700
rect 315948 4752 316000 4758
rect 315948 4694 316000 4700
rect 314568 4548 314620 4554
rect 314568 4490 314620 4496
rect 313280 4412 313332 4418
rect 313280 4354 313332 4360
rect 314580 3874 314608 4490
rect 315960 4078 315988 4694
rect 315948 4072 316000 4078
rect 315948 4014 316000 4020
rect 314568 3868 314620 3874
rect 314568 3810 314620 3816
rect 313188 3800 313240 3806
rect 313188 3742 313240 3748
rect 315764 3800 315816 3806
rect 315764 3742 315816 3748
rect 314568 3460 314620 3466
rect 314568 3402 314620 3408
rect 312544 3120 312596 3126
rect 312544 3062 312596 3068
rect 313372 3052 313424 3058
rect 313372 2994 313424 3000
rect 313384 480 313412 2994
rect 314580 480 314608 3402
rect 315776 480 315804 3742
rect 316604 3194 316632 4950
rect 317432 4894 317460 335650
rect 317524 333282 317552 340068
rect 317616 340054 317998 340082
rect 318076 340054 318458 340082
rect 318918 340054 319024 340082
rect 317616 335714 317644 340054
rect 317604 335708 317656 335714
rect 317604 335650 317656 335656
rect 317524 333254 317644 333282
rect 317510 134056 317566 134065
rect 317510 133991 317512 134000
rect 317564 133991 317566 134000
rect 317512 133962 317564 133968
rect 317616 8430 317644 333254
rect 318076 328522 318104 340054
rect 318800 333192 318852 333198
rect 318800 333134 318852 333140
rect 317892 328494 318104 328522
rect 317892 318918 317920 328494
rect 317880 318912 317932 318918
rect 317880 318854 317932 318860
rect 317788 318844 317840 318850
rect 317788 318786 317840 318792
rect 317604 8424 317656 8430
rect 317604 8366 317656 8372
rect 317800 7614 317828 318786
rect 317788 7608 317840 7614
rect 317788 7550 317840 7556
rect 318812 5080 318840 333134
rect 318996 8974 319024 340054
rect 319088 340054 319378 340082
rect 319456 340054 319746 340082
rect 320206 340054 320404 340082
rect 319088 333198 319116 340054
rect 319456 334218 319484 340054
rect 319536 337000 319588 337006
rect 319536 336942 319588 336948
rect 319444 334212 319496 334218
rect 319444 334154 319496 334160
rect 319548 334098 319576 336942
rect 320272 335640 320324 335646
rect 320272 335582 320324 335588
rect 319456 334070 319576 334098
rect 319076 333192 319128 333198
rect 319076 333134 319128 333140
rect 319168 328500 319220 328506
rect 319168 328442 319220 328448
rect 318984 8968 319036 8974
rect 318984 8910 319036 8916
rect 319180 7682 319208 328442
rect 319168 7676 319220 7682
rect 319168 7618 319220 7624
rect 318720 5052 318840 5080
rect 318720 4962 318748 5052
rect 318708 4956 318760 4962
rect 318708 4898 318760 4904
rect 318800 4956 318852 4962
rect 318800 4898 318852 4904
rect 317420 4888 317472 4894
rect 317420 4830 317472 4836
rect 316684 4820 316736 4826
rect 316684 4762 316736 4768
rect 316592 3188 316644 3194
rect 316592 3130 316644 3136
rect 316696 2854 316724 4762
rect 317420 4412 317472 4418
rect 317420 4354 317472 4360
rect 317432 4010 317460 4354
rect 317420 4004 317472 4010
rect 317420 3946 317472 3952
rect 316960 3868 317012 3874
rect 316960 3810 317012 3816
rect 316684 2848 316736 2854
rect 316684 2790 316736 2796
rect 316972 480 317000 3810
rect 318812 3602 318840 4898
rect 319260 4072 319312 4078
rect 319260 4014 319312 4020
rect 318800 3596 318852 3602
rect 318800 3538 318852 3544
rect 318064 2848 318116 2854
rect 318064 2790 318116 2796
rect 318076 480 318104 2790
rect 319272 480 319300 4014
rect 319456 3126 319484 334070
rect 320284 7750 320312 335582
rect 320376 9042 320404 340054
rect 320468 340054 320666 340082
rect 320744 340054 321126 340082
rect 321586 340054 321784 340082
rect 320364 9036 320416 9042
rect 320364 8978 320416 8984
rect 320272 7744 320324 7750
rect 320272 7686 320324 7692
rect 320468 5030 320496 340054
rect 320744 335646 320772 340054
rect 321468 337136 321520 337142
rect 321468 337078 321520 337084
rect 320732 335640 320784 335646
rect 320732 335582 320784 335588
rect 320456 5024 320508 5030
rect 320456 4966 320508 4972
rect 320180 4888 320232 4894
rect 320180 4830 320232 4836
rect 320192 3806 320220 4830
rect 321480 4010 321508 337078
rect 321652 335640 321704 335646
rect 321652 335582 321704 335588
rect 321664 7818 321692 335582
rect 321756 8362 321784 340054
rect 321848 340054 322046 340082
rect 322216 340054 322506 340082
rect 322966 340054 323164 340082
rect 321744 8356 321796 8362
rect 321744 8298 321796 8304
rect 321652 7812 321704 7818
rect 321652 7754 321704 7760
rect 321848 5098 321876 340054
rect 322216 335646 322244 340054
rect 322296 336796 322348 336802
rect 322296 336738 322348 336744
rect 322204 335640 322256 335646
rect 322204 335582 322256 335588
rect 322308 334098 322336 336738
rect 323032 335708 323084 335714
rect 323032 335650 323084 335656
rect 322216 334070 322336 334098
rect 321836 5092 321888 5098
rect 321836 5034 321888 5040
rect 320456 4004 320508 4010
rect 320456 3946 320508 3952
rect 321468 4004 321520 4010
rect 321468 3946 321520 3952
rect 320180 3800 320232 3806
rect 320180 3742 320232 3748
rect 319444 3120 319496 3126
rect 319444 3062 319496 3068
rect 320468 480 320496 3946
rect 321652 3392 321704 3398
rect 321652 3334 321704 3340
rect 321664 480 321692 3334
rect 322216 2990 322244 334070
rect 323044 7886 323072 335650
rect 323136 9110 323164 340054
rect 323216 335640 323268 335646
rect 323216 335582 323268 335588
rect 323228 9178 323256 335582
rect 323216 9172 323268 9178
rect 323216 9114 323268 9120
rect 323124 9104 323176 9110
rect 323124 9046 323176 9052
rect 323032 7880 323084 7886
rect 323032 7822 323084 7828
rect 323320 5166 323348 340068
rect 323504 340054 323794 340082
rect 323872 340054 324254 340082
rect 324332 340054 324714 340082
rect 323504 335714 323532 340054
rect 323492 335708 323544 335714
rect 323492 335650 323544 335656
rect 323872 335646 323900 340054
rect 323860 335640 323912 335646
rect 323860 335582 323912 335588
rect 324332 5234 324360 340054
rect 325160 338337 325188 340068
rect 325344 340054 325634 340082
rect 325712 340054 326094 340082
rect 326264 340054 326554 340082
rect 326632 340054 326922 340082
rect 327092 340054 327382 340082
rect 325146 338328 325202 338337
rect 325146 338263 325202 338272
rect 324594 338192 324650 338201
rect 324650 338150 324728 338178
rect 324594 338127 324650 338136
rect 324700 336734 324728 338150
rect 324688 336728 324740 336734
rect 324688 336670 324740 336676
rect 325344 335034 325372 340054
rect 324412 335028 324464 335034
rect 324412 334970 324464 334976
rect 325332 335028 325384 335034
rect 325332 334970 325384 334976
rect 324424 6186 324452 334970
rect 324780 328364 324832 328370
rect 324780 328306 324832 328312
rect 324792 321450 324820 328306
rect 324608 321422 324820 321450
rect 324608 318714 324636 321422
rect 324596 318708 324648 318714
rect 324596 318650 324648 318656
rect 324780 318708 324832 318714
rect 324780 318650 324832 318656
rect 324792 311794 324820 318650
rect 324700 311766 324820 311794
rect 324700 299470 324728 311766
rect 324688 299464 324740 299470
rect 324688 299406 324740 299412
rect 324596 289944 324648 289950
rect 324596 289886 324648 289892
rect 324608 289814 324636 289886
rect 324596 289808 324648 289814
rect 324596 289750 324648 289756
rect 324780 289740 324832 289746
rect 324780 289682 324832 289688
rect 324792 280158 324820 289682
rect 324504 280152 324556 280158
rect 324504 280094 324556 280100
rect 324780 280152 324832 280158
rect 324780 280094 324832 280100
rect 324516 278730 324544 280094
rect 324504 278724 324556 278730
rect 324504 278666 324556 278672
rect 324688 263492 324740 263498
rect 324688 263434 324740 263440
rect 324700 260846 324728 263434
rect 324688 260840 324740 260846
rect 324688 260782 324740 260788
rect 324596 251252 324648 251258
rect 324596 251194 324648 251200
rect 324608 251161 324636 251194
rect 324594 251152 324650 251161
rect 324594 251087 324650 251096
rect 324778 251152 324834 251161
rect 324778 251087 324834 251096
rect 324792 241534 324820 251087
rect 324780 241528 324832 241534
rect 324780 241470 324832 241476
rect 324872 241528 324924 241534
rect 324872 241470 324924 241476
rect 324884 231878 324912 241470
rect 324596 231872 324648 231878
rect 324594 231840 324596 231849
rect 324872 231872 324924 231878
rect 324648 231840 324650 231849
rect 324594 231775 324650 231784
rect 324870 231840 324872 231849
rect 324924 231840 324926 231849
rect 324870 231775 324926 231784
rect 324884 212566 324912 231775
rect 324596 212560 324648 212566
rect 324596 212502 324648 212508
rect 324872 212560 324924 212566
rect 324872 212502 324924 212508
rect 324608 207754 324636 212502
rect 324608 207726 324728 207754
rect 324700 193254 324728 207726
rect 324596 193248 324648 193254
rect 324596 193190 324648 193196
rect 324688 193248 324740 193254
rect 324688 193190 324740 193196
rect 324608 186266 324636 193190
rect 324608 186238 324728 186266
rect 324700 182170 324728 186238
rect 324504 182164 324556 182170
rect 324504 182106 324556 182112
rect 324688 182164 324740 182170
rect 324688 182106 324740 182112
rect 324516 172553 324544 182106
rect 324502 172544 324558 172553
rect 324502 172479 324558 172488
rect 324686 172544 324742 172553
rect 324686 172479 324742 172488
rect 324700 164218 324728 172479
rect 324688 164212 324740 164218
rect 324688 164154 324740 164160
rect 324596 154624 324648 154630
rect 324596 154566 324648 154572
rect 324608 147762 324636 154566
rect 324596 147756 324648 147762
rect 324596 147698 324648 147704
rect 324596 147620 324648 147626
rect 324596 147562 324648 147568
rect 324608 144945 324636 147562
rect 324594 144936 324650 144945
rect 324594 144871 324650 144880
rect 324778 144936 324834 144945
rect 324778 144871 324834 144880
rect 324792 135425 324820 144871
rect 324778 135416 324834 135425
rect 324778 135351 324834 135360
rect 324594 135280 324650 135289
rect 324594 135215 324650 135224
rect 324608 131102 324636 135215
rect 324596 131096 324648 131102
rect 324596 131038 324648 131044
rect 324872 131096 324924 131102
rect 324872 131038 324924 131044
rect 324884 115977 324912 131038
rect 324686 115968 324742 115977
rect 324686 115903 324742 115912
rect 324870 115968 324926 115977
rect 324870 115903 324926 115912
rect 324700 106350 324728 115903
rect 324688 106344 324740 106350
rect 324688 106286 324740 106292
rect 324688 104916 324740 104922
rect 324688 104858 324740 104864
rect 324700 99482 324728 104858
rect 324688 99476 324740 99482
rect 324688 99418 324740 99424
rect 324596 99340 324648 99346
rect 324596 99282 324648 99288
rect 324608 82414 324636 99282
rect 324596 82408 324648 82414
rect 324596 82350 324648 82356
rect 324596 82272 324648 82278
rect 324596 82214 324648 82220
rect 324608 67794 324636 82214
rect 324596 67788 324648 67794
rect 324596 67730 324648 67736
rect 324596 67652 324648 67658
rect 324596 67594 324648 67600
rect 324608 66230 324636 67594
rect 324596 66224 324648 66230
rect 324596 66166 324648 66172
rect 324780 53100 324832 53106
rect 324780 53042 324832 53048
rect 324792 38622 324820 53042
rect 324780 38616 324832 38622
rect 324780 38558 324832 38564
rect 324780 38480 324832 38486
rect 324780 38422 324832 38428
rect 324792 33674 324820 38422
rect 324608 33646 324820 33674
rect 324608 28966 324636 33646
rect 325606 29608 325662 29617
rect 325606 29543 325662 29552
rect 325620 29345 325648 29543
rect 325606 29336 325662 29345
rect 325606 29271 325662 29280
rect 324596 28960 324648 28966
rect 324596 28902 324648 28908
rect 324596 19372 324648 19378
rect 324596 19314 324648 19320
rect 324608 7954 324636 19314
rect 324596 7948 324648 7954
rect 324596 7890 324648 7896
rect 324412 6180 324464 6186
rect 324412 6122 324464 6128
rect 324320 5228 324372 5234
rect 324320 5170 324372 5176
rect 323308 5160 323360 5166
rect 323308 5102 323360 5108
rect 325712 4622 325740 340054
rect 325792 335640 325844 335646
rect 326264 335594 326292 340054
rect 326344 336864 326396 336870
rect 326344 336806 326396 336812
rect 325792 335582 325844 335588
rect 325804 6254 325832 335582
rect 325988 335566 326292 335594
rect 325988 321638 326016 335566
rect 325976 321632 326028 321638
rect 325976 321574 326028 321580
rect 326068 321428 326120 321434
rect 326068 321370 326120 321376
rect 326080 294710 326108 321370
rect 326068 294704 326120 294710
rect 326068 294646 326120 294652
rect 325976 289876 326028 289882
rect 325976 289818 326028 289824
rect 325988 273222 326016 289818
rect 325976 273216 326028 273222
rect 325976 273158 326028 273164
rect 325976 273080 326028 273086
rect 325976 273022 326028 273028
rect 325988 253910 326016 273022
rect 325976 253904 326028 253910
rect 325976 253846 326028 253852
rect 325976 253768 326028 253774
rect 325976 253710 326028 253716
rect 325988 234598 326016 253710
rect 325976 234592 326028 234598
rect 325976 234534 326028 234540
rect 325976 234456 326028 234462
rect 325976 234398 326028 234404
rect 325988 215286 326016 234398
rect 325976 215280 326028 215286
rect 325976 215222 326028 215228
rect 325976 215144 326028 215150
rect 325976 215086 326028 215092
rect 325988 195974 326016 215086
rect 325976 195968 326028 195974
rect 325976 195910 326028 195916
rect 325976 195832 326028 195838
rect 325976 195774 326028 195780
rect 325988 176746 326016 195774
rect 325896 176718 326016 176746
rect 325896 176610 325924 176718
rect 325896 176582 326016 176610
rect 325988 157350 326016 176582
rect 325976 157344 326028 157350
rect 325976 157286 326028 157292
rect 325976 157208 326028 157214
rect 325976 157150 326028 157156
rect 325988 99498 326016 157150
rect 325896 99470 326016 99498
rect 325896 99362 325924 99470
rect 325896 99334 326016 99362
rect 325988 80102 326016 99334
rect 325976 80096 326028 80102
rect 325976 80038 326028 80044
rect 325976 79960 326028 79966
rect 325976 79902 326028 79908
rect 325988 67726 326016 79902
rect 325976 67720 326028 67726
rect 325976 67662 326028 67668
rect 325884 67652 325936 67658
rect 325884 67594 325936 67600
rect 325896 58070 325924 67594
rect 325884 58064 325936 58070
rect 325884 58006 325936 58012
rect 325884 57928 325936 57934
rect 325884 57870 325936 57876
rect 325896 46850 325924 57870
rect 325884 46844 325936 46850
rect 325884 46786 325936 46792
rect 326160 46844 326212 46850
rect 326160 46786 326212 46792
rect 326172 38570 326200 46786
rect 326080 38542 326200 38570
rect 326080 24426 326108 38542
rect 325988 24398 326108 24426
rect 325988 12510 326016 24398
rect 325976 12504 326028 12510
rect 325976 12446 326028 12452
rect 325884 12436 325936 12442
rect 325884 12378 325936 12384
rect 325896 8022 325924 12378
rect 325884 8016 325936 8022
rect 325884 7958 325936 7964
rect 325792 6248 325844 6254
rect 325792 6190 325844 6196
rect 326356 4740 326384 336806
rect 326632 335646 326660 340054
rect 326620 335640 326672 335646
rect 326620 335582 326672 335588
rect 326986 181384 327042 181393
rect 326986 181319 327042 181328
rect 327000 181121 327028 181319
rect 326986 181112 327042 181121
rect 326986 181047 327042 181056
rect 326896 134020 326948 134026
rect 326896 133962 326948 133968
rect 326908 133906 326936 133962
rect 326986 133920 327042 133929
rect 326908 133878 326986 133906
rect 326986 133855 327042 133864
rect 326986 87272 327042 87281
rect 326986 87207 327042 87216
rect 327000 87009 327028 87207
rect 326986 87000 327042 87009
rect 326986 86935 327042 86944
rect 326804 63776 326856 63782
rect 326802 63744 326804 63753
rect 326856 63744 326858 63753
rect 326802 63679 326858 63688
rect 326172 4712 326384 4740
rect 325700 4616 325752 4622
rect 325700 4558 325752 4564
rect 325240 3800 325292 3806
rect 325240 3742 325292 3748
rect 324044 3596 324096 3602
rect 324044 3538 324096 3544
rect 322204 2984 322256 2990
rect 322204 2926 322256 2932
rect 322848 2916 322900 2922
rect 322848 2858 322900 2864
rect 322860 480 322888 2858
rect 324056 480 324084 3538
rect 325252 480 325280 3742
rect 326172 2990 326200 4712
rect 327092 4690 327120 340054
rect 327172 335640 327224 335646
rect 327172 335582 327224 335588
rect 327184 6322 327212 335582
rect 327460 331226 327488 340190
rect 327920 340054 328302 340082
rect 327724 337000 327776 337006
rect 327724 336942 327776 336948
rect 327448 331220 327500 331226
rect 327448 331162 327500 331168
rect 327448 328500 327500 328506
rect 327448 328442 327500 328448
rect 327460 318782 327488 328442
rect 327448 318776 327500 318782
rect 327448 318718 327500 318724
rect 327448 309188 327500 309194
rect 327448 309130 327500 309136
rect 327460 299470 327488 309130
rect 327264 299464 327316 299470
rect 327264 299406 327316 299412
rect 327448 299464 327500 299470
rect 327448 299406 327500 299412
rect 327276 298110 327304 299406
rect 327264 298104 327316 298110
rect 327264 298046 327316 298052
rect 327540 288448 327592 288454
rect 327540 288390 327592 288396
rect 327552 280158 327580 288390
rect 327540 280152 327592 280158
rect 327540 280094 327592 280100
rect 327356 280084 327408 280090
rect 327356 280026 327408 280032
rect 327368 278769 327396 280026
rect 327354 278760 327410 278769
rect 327354 278695 327410 278704
rect 327630 278760 327686 278769
rect 327630 278695 327686 278704
rect 327644 253722 327672 278695
rect 327368 253694 327672 253722
rect 327368 251190 327396 253694
rect 327356 251184 327408 251190
rect 327356 251126 327408 251132
rect 327264 242684 327316 242690
rect 327264 242626 327316 242632
rect 327276 240106 327304 242626
rect 327264 240100 327316 240106
rect 327264 240042 327316 240048
rect 327356 240100 327408 240106
rect 327356 240042 327408 240048
rect 327368 230489 327396 240042
rect 327354 230480 327410 230489
rect 327354 230415 327410 230424
rect 327538 230480 327594 230489
rect 327538 230415 327594 230424
rect 327552 220862 327580 230415
rect 327356 220856 327408 220862
rect 327356 220798 327408 220804
rect 327540 220856 327592 220862
rect 327540 220798 327592 220804
rect 327368 215422 327396 220798
rect 327356 215416 327408 215422
rect 327356 215358 327408 215364
rect 327356 215280 327408 215286
rect 327356 215222 327408 215228
rect 327368 211138 327396 215222
rect 327356 211132 327408 211138
rect 327356 211074 327408 211080
rect 327540 211132 327592 211138
rect 327540 211074 327592 211080
rect 327552 201521 327580 211074
rect 327354 201512 327410 201521
rect 327354 201447 327410 201456
rect 327538 201512 327594 201521
rect 327538 201447 327594 201456
rect 327368 196110 327396 201447
rect 327356 196104 327408 196110
rect 327356 196046 327408 196052
rect 327356 195968 327408 195974
rect 327356 195910 327408 195916
rect 327368 186386 327396 195910
rect 327356 186380 327408 186386
rect 327356 186322 327408 186328
rect 327448 186244 327500 186250
rect 327448 186186 327500 186192
rect 327460 180810 327488 186186
rect 327448 180804 327500 180810
rect 327448 180746 327500 180752
rect 327356 171148 327408 171154
rect 327356 171090 327408 171096
rect 327368 153542 327396 171090
rect 327356 153536 327408 153542
rect 327356 153478 327408 153484
rect 327356 147620 327408 147626
rect 327356 147562 327408 147568
rect 327368 144922 327396 147562
rect 327368 144894 327488 144922
rect 327460 138281 327488 144894
rect 327446 138272 327502 138281
rect 327446 138207 327502 138216
rect 327354 135280 327410 135289
rect 327354 135215 327356 135224
rect 327408 135215 327410 135224
rect 327356 135186 327408 135192
rect 327264 133952 327316 133958
rect 327262 133920 327264 133929
rect 327316 133920 327318 133929
rect 327262 133855 327318 133864
rect 327356 128308 327408 128314
rect 327356 128250 327408 128256
rect 327368 125610 327396 128250
rect 327368 125582 327488 125610
rect 327460 120850 327488 125582
rect 327460 120822 327580 120850
rect 327552 106457 327580 120822
rect 327538 106448 327594 106457
rect 327538 106383 327594 106392
rect 327446 106312 327502 106321
rect 327446 106247 327502 106256
rect 327460 104854 327488 106247
rect 327448 104848 327500 104854
rect 327448 104790 327500 104796
rect 327356 95260 327408 95266
rect 327356 95202 327408 95208
rect 327368 86902 327396 95202
rect 327356 86896 327408 86902
rect 327356 86838 327408 86844
rect 327356 77308 327408 77314
rect 327356 77250 327408 77256
rect 327368 67658 327396 77250
rect 327356 67652 327408 67658
rect 327356 67594 327408 67600
rect 327356 66292 327408 66298
rect 327356 66234 327408 66240
rect 327368 53174 327396 66234
rect 327356 53168 327408 53174
rect 327356 53110 327408 53116
rect 327264 53100 327316 53106
rect 327264 53042 327316 53048
rect 327276 38706 327304 53042
rect 327276 38678 327396 38706
rect 327368 33810 327396 38678
rect 327276 33782 327396 33810
rect 327276 31634 327304 33782
rect 327276 31606 327488 31634
rect 327460 28966 327488 31606
rect 327264 28960 327316 28966
rect 327264 28902 327316 28908
rect 327448 28960 327500 28966
rect 327448 28902 327500 28908
rect 327276 19394 327304 28902
rect 327276 19366 327396 19394
rect 327368 19310 327396 19366
rect 327356 19304 327408 19310
rect 327356 19246 327408 19252
rect 327264 9716 327316 9722
rect 327264 9658 327316 9664
rect 327276 8090 327304 9658
rect 327264 8084 327316 8090
rect 327264 8026 327316 8032
rect 327172 6316 327224 6322
rect 327172 6258 327224 6264
rect 327080 4684 327132 4690
rect 327080 4626 327132 4632
rect 326436 3528 326488 3534
rect 326264 3476 326436 3482
rect 326264 3470 326488 3476
rect 326264 3454 326476 3470
rect 326264 3398 326292 3454
rect 326252 3392 326304 3398
rect 326252 3334 326304 3340
rect 327632 3188 327684 3194
rect 327632 3130 327684 3136
rect 326160 2984 326212 2990
rect 326160 2926 326212 2932
rect 326436 2848 326488 2854
rect 326436 2790 326488 2796
rect 326448 480 326476 2790
rect 327644 480 327672 3130
rect 327736 2922 327764 336942
rect 327816 336796 327868 336802
rect 327816 336738 327868 336744
rect 327828 4010 327856 336738
rect 327920 335646 327948 340054
rect 327908 335640 327960 335646
rect 327908 335582 327960 335588
rect 328748 331242 328776 340068
rect 328656 331214 328776 331242
rect 328840 340054 329222 340082
rect 328552 328500 328604 328506
rect 328552 328442 328604 328448
rect 328564 318782 328592 328442
rect 328552 318776 328604 318782
rect 328552 318718 328604 318724
rect 328656 311914 328684 331214
rect 328840 328506 328868 340054
rect 329668 337754 329696 340068
rect 330036 340054 330142 340082
rect 330312 340054 330602 340082
rect 330680 340054 330970 340082
rect 329656 337748 329708 337754
rect 329656 337690 329708 337696
rect 329932 335640 329984 335646
rect 329932 335582 329984 335588
rect 328828 328500 328880 328506
rect 328828 328442 328880 328448
rect 328736 318776 328788 318782
rect 328736 318718 328788 318724
rect 328644 311908 328696 311914
rect 328644 311850 328696 311856
rect 328644 311704 328696 311710
rect 328644 311646 328696 311652
rect 328552 292596 328604 292602
rect 328552 292538 328604 292544
rect 328564 282962 328592 292538
rect 328472 282934 328592 282962
rect 328472 282826 328500 282934
rect 328472 282798 328592 282826
rect 328564 263650 328592 282798
rect 328472 263622 328592 263650
rect 328472 263514 328500 263622
rect 328472 263486 328592 263514
rect 328564 244338 328592 263486
rect 328472 244310 328592 244338
rect 328472 244202 328500 244310
rect 328472 244174 328592 244202
rect 328564 225026 328592 244174
rect 328472 224998 328592 225026
rect 328472 224890 328500 224998
rect 328472 224862 328592 224890
rect 328564 205714 328592 224862
rect 328472 205686 328592 205714
rect 328472 205578 328500 205686
rect 328472 205550 328592 205578
rect 328564 186402 328592 205550
rect 328472 186374 328592 186402
rect 328472 186266 328500 186374
rect 328472 186238 328592 186266
rect 328564 167090 328592 186238
rect 328472 167062 328592 167090
rect 328472 166954 328500 167062
rect 328472 166926 328592 166954
rect 328564 147778 328592 166926
rect 328472 147750 328592 147778
rect 328472 147642 328500 147750
rect 328472 147614 328592 147642
rect 328564 135250 328592 147614
rect 328552 135244 328604 135250
rect 328552 135186 328604 135192
rect 328458 125624 328514 125633
rect 328458 125559 328460 125568
rect 328512 125559 328514 125568
rect 328460 125530 328512 125536
rect 328552 118652 328604 118658
rect 328552 118594 328604 118600
rect 328564 109154 328592 118594
rect 328472 109126 328592 109154
rect 328472 109018 328500 109126
rect 328472 108990 328592 109018
rect 328564 89842 328592 108990
rect 328472 89814 328592 89842
rect 328472 89706 328500 89814
rect 328472 89678 328592 89706
rect 328564 70514 328592 89678
rect 328552 70508 328604 70514
rect 328552 70450 328604 70456
rect 328552 70372 328604 70378
rect 328552 70314 328604 70320
rect 328564 51082 328592 70314
rect 328472 51054 328592 51082
rect 328472 50946 328500 51054
rect 328472 50918 328592 50946
rect 328366 40624 328422 40633
rect 328366 40559 328422 40568
rect 328380 40225 328408 40559
rect 328366 40216 328422 40225
rect 328366 40151 328422 40160
rect 328564 31890 328592 50918
rect 328552 31884 328604 31890
rect 328552 31826 328604 31832
rect 328552 27668 328604 27674
rect 328552 27610 328604 27616
rect 328564 22778 328592 27610
rect 328552 22772 328604 22778
rect 328552 22714 328604 22720
rect 328552 12368 328604 12374
rect 328552 12310 328604 12316
rect 328564 9602 328592 12310
rect 328472 9574 328592 9602
rect 328472 8158 328500 9574
rect 328460 8152 328512 8158
rect 328460 8094 328512 8100
rect 328656 4486 328684 311646
rect 328748 292602 328776 318718
rect 328736 292596 328788 292602
rect 328736 292538 328788 292544
rect 328736 135244 328788 135250
rect 328736 135186 328788 135192
rect 328748 125633 328776 135186
rect 328734 125624 328790 125633
rect 328734 125559 328790 125568
rect 329944 8226 329972 335582
rect 329932 8220 329984 8226
rect 329932 8162 329984 8168
rect 330036 4554 330064 340054
rect 330312 335646 330340 340054
rect 330680 337770 330708 340054
rect 330404 337742 330708 337770
rect 331128 337748 331180 337754
rect 330404 337618 330432 337742
rect 331128 337690 331180 337696
rect 330392 337612 330444 337618
rect 330392 337554 330444 337560
rect 330484 337612 330536 337618
rect 330484 337554 330536 337560
rect 330300 335640 330352 335646
rect 330300 335582 330352 335588
rect 330024 4548 330076 4554
rect 330024 4490 330076 4496
rect 328644 4480 328696 4486
rect 328644 4422 328696 4428
rect 327816 4004 327868 4010
rect 327816 3946 327868 3952
rect 330024 4004 330076 4010
rect 330024 3946 330076 3952
rect 328828 3732 328880 3738
rect 328828 3674 328880 3680
rect 327724 2916 327776 2922
rect 327724 2858 327776 2864
rect 328840 480 328868 3674
rect 330036 480 330064 3946
rect 330496 3806 330524 337554
rect 331140 4010 331168 337690
rect 331416 4758 331444 340068
rect 331876 337482 331904 340068
rect 331864 337476 331916 337482
rect 331864 337418 331916 337424
rect 332336 337385 332364 340068
rect 332322 337376 332378 337385
rect 332322 337311 332378 337320
rect 331404 4752 331456 4758
rect 331404 4694 331456 4700
rect 332796 4418 332824 340068
rect 333256 337550 333284 340068
rect 333716 337686 333744 340068
rect 333704 337680 333756 337686
rect 333704 337622 333756 337628
rect 333244 337544 333296 337550
rect 333244 337486 333296 337492
rect 333888 337476 333940 337482
rect 333888 337418 333940 337424
rect 332784 4412 332836 4418
rect 332784 4354 332836 4360
rect 331128 4004 331180 4010
rect 331128 3946 331180 3952
rect 330484 3800 330536 3806
rect 330484 3742 330536 3748
rect 332416 3392 332468 3398
rect 332416 3334 332468 3340
rect 331220 2916 331272 2922
rect 331220 2858 331272 2864
rect 331232 480 331260 2858
rect 332428 480 332456 3334
rect 333900 626 333928 337418
rect 334176 6390 334204 340068
rect 334544 337958 334572 340068
rect 334636 340054 335018 340082
rect 335478 340054 335584 340082
rect 334532 337952 334584 337958
rect 334532 337894 334584 337900
rect 334636 337770 334664 340054
rect 334716 337952 334768 337958
rect 334716 337894 334768 337900
rect 334544 337742 334664 337770
rect 334544 337414 334572 337742
rect 334624 337544 334676 337550
rect 334624 337486 334676 337492
rect 334532 337408 334584 337414
rect 334532 337350 334584 337356
rect 334164 6384 334216 6390
rect 334164 6326 334216 6332
rect 334636 3738 334664 337486
rect 334624 3732 334676 3738
rect 334624 3674 334676 3680
rect 334728 3074 334756 337894
rect 334808 337408 334860 337414
rect 334808 337350 334860 337356
rect 334820 3534 334848 337350
rect 335266 63880 335322 63889
rect 335266 63815 335322 63824
rect 335280 63782 335308 63815
rect 335268 63776 335320 63782
rect 335268 63718 335320 63724
rect 335556 5302 335584 340054
rect 335924 338026 335952 340068
rect 335912 338020 335964 338026
rect 335912 337962 335964 337968
rect 336384 337414 336412 340068
rect 336372 337408 336424 337414
rect 336372 337350 336424 337356
rect 336646 134192 336702 134201
rect 336646 134127 336702 134136
rect 336660 133958 336688 134127
rect 336648 133952 336700 133958
rect 336648 133894 336700 133900
rect 336646 87272 336702 87281
rect 336646 87207 336702 87216
rect 336660 87009 336688 87207
rect 336646 87000 336702 87009
rect 336646 86935 336702 86944
rect 336844 5370 336872 340068
rect 337304 337822 337332 340068
rect 337292 337816 337344 337822
rect 337292 337758 337344 337764
rect 337396 337634 337424 340190
rect 363892 340134 363920 340190
rect 363052 340128 363104 340134
rect 338146 340054 338252 340082
rect 336936 337606 337424 337634
rect 336936 60722 336964 337606
rect 338028 337340 338080 337346
rect 338028 337282 338080 337288
rect 338040 180946 338068 337282
rect 338028 180940 338080 180946
rect 338028 180882 338080 180888
rect 338028 180804 338080 180810
rect 338028 180746 338080 180752
rect 336924 60716 336976 60722
rect 336924 60658 336976 60664
rect 337108 60716 337160 60722
rect 337108 60658 337160 60664
rect 337120 57934 337148 60658
rect 337108 57928 337160 57934
rect 337108 57870 337160 57876
rect 336924 48340 336976 48346
rect 336924 48282 336976 48288
rect 336936 48249 336964 48282
rect 336922 48240 336978 48249
rect 336922 48175 336978 48184
rect 337014 48104 337070 48113
rect 337014 48039 337070 48048
rect 337028 22114 337056 48039
rect 337934 40624 337990 40633
rect 337934 40559 337990 40568
rect 337948 40089 337976 40559
rect 337934 40080 337990 40089
rect 337934 40015 337990 40024
rect 336936 22086 337056 22114
rect 336832 5364 336884 5370
rect 336832 5306 336884 5312
rect 335544 5296 335596 5302
rect 335544 5238 335596 5244
rect 334808 3528 334860 3534
rect 334808 3470 334860 3476
rect 336936 3262 336964 22086
rect 338040 3738 338068 180746
rect 338224 5438 338252 340054
rect 338316 340054 338606 340082
rect 338212 5432 338264 5438
rect 338212 5374 338264 5380
rect 337108 3732 337160 3738
rect 337108 3674 337160 3680
rect 338028 3732 338080 3738
rect 338028 3674 338080 3680
rect 336924 3256 336976 3262
rect 336924 3198 336976 3204
rect 334636 3046 334756 3074
rect 334636 2990 334664 3046
rect 334624 2984 334676 2990
rect 334624 2926 334676 2932
rect 334716 2984 334768 2990
rect 334716 2926 334768 2932
rect 333624 598 333928 626
rect 333624 480 333652 598
rect 334728 480 334756 2926
rect 335912 2848 335964 2854
rect 335912 2790 335964 2796
rect 335924 480 335952 2790
rect 337120 480 337148 3674
rect 338316 3670 338344 340054
rect 339052 337074 339080 340068
rect 339526 340054 339632 340082
rect 339040 337068 339092 337074
rect 339040 337010 339092 337016
rect 338764 336864 338816 336870
rect 338764 336806 338816 336812
rect 338304 3664 338356 3670
rect 338304 3606 338356 3612
rect 338776 3330 338804 336806
rect 339604 5506 339632 340054
rect 339972 337890 340000 340068
rect 340156 340054 340446 340082
rect 340906 340054 341012 340082
rect 339960 337884 340012 337890
rect 339960 337826 340012 337832
rect 340156 337736 340184 340054
rect 339696 337708 340184 337736
rect 339592 5500 339644 5506
rect 339592 5442 339644 5448
rect 339696 3942 339724 337708
rect 340788 337680 340840 337686
rect 340788 337622 340840 337628
rect 340800 4876 340828 337622
rect 340708 4848 340828 4876
rect 339684 3936 339736 3942
rect 339684 3878 339736 3884
rect 339500 3732 339552 3738
rect 339500 3674 339552 3680
rect 338764 3324 338816 3330
rect 338764 3266 338816 3272
rect 338304 3256 338356 3262
rect 338304 3198 338356 3204
rect 338316 480 338344 3198
rect 339512 480 339540 3674
rect 340708 480 340736 4848
rect 340984 4350 341012 340054
rect 341352 337210 341380 340068
rect 341812 338094 341840 340068
rect 341904 340054 342194 340082
rect 341800 338088 341852 338094
rect 341800 338030 341852 338036
rect 341340 337204 341392 337210
rect 341340 337146 341392 337152
rect 341904 335594 341932 340054
rect 341984 337000 342036 337006
rect 341984 336942 342036 336948
rect 341076 335566 341932 335594
rect 340972 4344 341024 4350
rect 340972 4286 341024 4292
rect 341076 4282 341104 335566
rect 341996 335458 342024 336942
rect 342640 336802 342668 340068
rect 343100 337142 343128 340068
rect 343284 340054 343574 340082
rect 343088 337136 343140 337142
rect 343088 337078 343140 337084
rect 342628 336796 342680 336802
rect 342628 336738 342680 336744
rect 343284 335594 343312 340054
rect 344020 337822 344048 340068
rect 344480 338026 344508 340068
rect 344572 340054 344954 340082
rect 344468 338020 344520 338026
rect 344468 337962 344520 337968
rect 344008 337816 344060 337822
rect 344008 337758 344060 337764
rect 341536 335430 342024 335458
rect 342548 335566 343312 335594
rect 344572 335578 344600 340054
rect 345204 339108 345256 339114
rect 345204 339050 345256 339056
rect 344928 337816 344980 337822
rect 344928 337758 344980 337764
rect 344744 336932 344796 336938
rect 344744 336874 344796 336880
rect 344652 336864 344704 336870
rect 344652 336806 344704 336812
rect 344560 335572 344612 335578
rect 341064 4276 341116 4282
rect 341064 4218 341116 4224
rect 341536 3126 341564 335430
rect 342548 321722 342576 335566
rect 344560 335514 344612 335520
rect 344664 335458 344692 336806
rect 344296 335430 344692 335458
rect 343824 328500 343876 328506
rect 343824 328442 343876 328448
rect 342548 321694 342668 321722
rect 342640 318866 342668 321694
rect 342548 318838 342668 318866
rect 342548 318782 342576 318838
rect 342536 318776 342588 318782
rect 342536 318718 342588 318724
rect 342536 309188 342588 309194
rect 342456 309148 342536 309176
rect 342456 307766 342484 309148
rect 342536 309130 342588 309136
rect 342444 307760 342496 307766
rect 342444 307702 342496 307708
rect 342536 298172 342588 298178
rect 342536 298114 342588 298120
rect 342548 292670 342576 298114
rect 342536 292664 342588 292670
rect 342536 292606 342588 292612
rect 342536 292528 342588 292534
rect 342536 292470 342588 292476
rect 342548 280158 342576 292470
rect 343836 282962 343864 328442
rect 343744 282934 343864 282962
rect 343744 282826 343772 282934
rect 343744 282798 343864 282826
rect 342536 280152 342588 280158
rect 342536 280094 342588 280100
rect 342536 270564 342588 270570
rect 342536 270506 342588 270512
rect 342548 260846 342576 270506
rect 343836 263650 343864 282798
rect 343744 263622 343864 263650
rect 343744 263514 343772 263622
rect 343744 263486 343864 263514
rect 342536 260840 342588 260846
rect 342536 260782 342588 260788
rect 342536 251252 342588 251258
rect 342536 251194 342588 251200
rect 342548 241505 342576 251194
rect 343836 244338 343864 263486
rect 343744 244310 343864 244338
rect 343744 244202 343772 244310
rect 343744 244174 343864 244202
rect 342350 241496 342406 241505
rect 342350 241431 342406 241440
rect 342534 241496 342590 241505
rect 342534 241431 342590 241440
rect 342364 231878 342392 241431
rect 342352 231872 342404 231878
rect 342352 231814 342404 231820
rect 342536 231872 342588 231878
rect 342536 231814 342588 231820
rect 342548 222193 342576 231814
rect 343836 225026 343864 244174
rect 343744 224998 343864 225026
rect 343744 224890 343772 224998
rect 343744 224862 343864 224890
rect 342350 222184 342406 222193
rect 342350 222119 342406 222128
rect 342534 222184 342590 222193
rect 342534 222119 342590 222128
rect 342364 212566 342392 222119
rect 343836 212566 343864 224862
rect 342352 212560 342404 212566
rect 342352 212502 342404 212508
rect 342536 212560 342588 212566
rect 342536 212502 342588 212508
rect 343824 212560 343876 212566
rect 343824 212502 343876 212508
rect 342548 196058 342576 212502
rect 343732 212492 343784 212498
rect 343732 212434 343784 212440
rect 343744 211138 343772 212434
rect 343732 211132 343784 211138
rect 343732 211074 343784 211080
rect 343732 202836 343784 202842
rect 343732 202778 343784 202784
rect 343744 196058 343772 202778
rect 342456 196030 342576 196058
rect 343652 196030 343772 196058
rect 342456 195922 342484 196030
rect 342456 195894 342576 195922
rect 342548 193225 342576 195894
rect 342350 193216 342406 193225
rect 342350 193151 342406 193160
rect 342534 193216 342590 193225
rect 343652 193202 343680 196030
rect 343652 193174 343864 193202
rect 342534 193151 342590 193160
rect 342364 183598 342392 193151
rect 342352 183592 342404 183598
rect 342352 183534 342404 183540
rect 342536 183592 342588 183598
rect 342536 183534 342588 183540
rect 342548 164393 342576 183534
rect 343836 183530 343864 193174
rect 343824 183524 343876 183530
rect 343824 183466 343876 183472
rect 343916 183524 343968 183530
rect 343916 183466 343968 183472
rect 343928 182170 343956 183466
rect 343916 182164 343968 182170
rect 343916 182106 343968 182112
rect 344100 182164 344152 182170
rect 344100 182106 344152 182112
rect 344112 172553 344140 182106
rect 343914 172544 343970 172553
rect 343914 172479 343970 172488
rect 344098 172544 344154 172553
rect 344098 172479 344154 172488
rect 343928 164393 343956 172479
rect 342534 164384 342590 164393
rect 342534 164319 342590 164328
rect 343914 164384 343970 164393
rect 343914 164319 343970 164328
rect 342534 164248 342590 164257
rect 342534 164183 342590 164192
rect 343914 164248 343970 164257
rect 343914 164183 343970 164192
rect 342548 162858 342576 164183
rect 343928 162858 343956 164183
rect 342536 162852 342588 162858
rect 342536 162794 342588 162800
rect 342628 162852 342680 162858
rect 342628 162794 342680 162800
rect 343916 162852 343968 162858
rect 343916 162794 343968 162800
rect 342640 135266 342668 162794
rect 343916 153264 343968 153270
rect 343916 153206 343968 153212
rect 343928 148374 343956 153206
rect 343916 148368 343968 148374
rect 343916 148310 343968 148316
rect 342548 135238 342668 135266
rect 343824 135312 343876 135318
rect 343824 135254 343876 135260
rect 342548 119082 342576 135238
rect 342548 119054 342760 119082
rect 342732 114617 342760 119054
rect 342534 114608 342590 114617
rect 342534 114543 342590 114552
rect 342718 114608 342774 114617
rect 342718 114543 342774 114552
rect 342548 114510 342576 114543
rect 342536 114504 342588 114510
rect 342536 114446 342588 114452
rect 343836 109154 343864 135254
rect 343744 109126 343864 109154
rect 343744 109018 343772 109126
rect 343744 108990 343864 109018
rect 342536 104984 342588 104990
rect 342536 104926 342588 104932
rect 342548 104854 342576 104926
rect 342536 104848 342588 104854
rect 342536 104790 342588 104796
rect 342536 95260 342588 95266
rect 342536 95202 342588 95208
rect 342548 80170 342576 95202
rect 343836 86970 343864 108990
rect 343732 86964 343784 86970
rect 343732 86906 343784 86912
rect 343824 86964 343876 86970
rect 343824 86906 343876 86912
rect 343744 85542 343772 86906
rect 343732 85536 343784 85542
rect 343732 85478 343784 85484
rect 342536 80164 342588 80170
rect 342536 80106 342588 80112
rect 342536 80028 342588 80034
rect 342536 79970 342588 79976
rect 342548 51202 342576 79970
rect 343732 76016 343784 76022
rect 343732 75958 343784 75964
rect 343744 75886 343772 75958
rect 343732 75880 343784 75886
rect 343732 75822 343784 75828
rect 343916 66292 343968 66298
rect 343916 66234 343968 66240
rect 343928 60738 343956 66234
rect 343836 60710 343956 60738
rect 342536 51196 342588 51202
rect 342536 51138 342588 51144
rect 342536 46980 342588 46986
rect 342536 46922 342588 46928
rect 342548 46866 342576 46922
rect 342456 46838 342576 46866
rect 342456 29102 342484 46838
rect 343836 41426 343864 60710
rect 343744 41398 343864 41426
rect 343744 41290 343772 41398
rect 343744 41262 343864 41290
rect 342444 29096 342496 29102
rect 342444 29038 342496 29044
rect 342536 29028 342588 29034
rect 342536 28970 342588 28976
rect 342548 27606 342576 28970
rect 342536 27600 342588 27606
rect 342536 27542 342588 27548
rect 343836 12458 343864 41262
rect 343744 12430 343864 12458
rect 342444 9716 342496 9722
rect 342444 9658 342496 9664
rect 342456 4214 342484 9658
rect 343744 6458 343772 12430
rect 343732 6452 343784 6458
rect 343732 6394 343784 6400
rect 344296 4298 344324 335430
rect 344756 335322 344784 336874
rect 344204 4270 344324 4298
rect 344388 335294 344784 335322
rect 342444 4208 342496 4214
rect 342444 4150 342496 4156
rect 343088 3936 343140 3942
rect 343088 3878 343140 3884
rect 341892 3664 341944 3670
rect 341892 3606 341944 3612
rect 341524 3120 341576 3126
rect 341524 3062 341576 3068
rect 341904 480 341932 3606
rect 343100 480 343128 3878
rect 344204 3874 344232 4270
rect 344284 4140 344336 4146
rect 344284 4082 344336 4088
rect 344192 3868 344244 3874
rect 344192 3810 344244 3816
rect 344296 480 344324 4082
rect 344388 4078 344416 335294
rect 344940 4146 344968 337758
rect 345112 335640 345164 335646
rect 345112 335582 345164 335588
rect 345124 193322 345152 335582
rect 345216 329066 345244 339050
rect 345400 337958 345428 340068
rect 345768 339114 345796 340068
rect 345952 340054 346242 340082
rect 345756 339108 345808 339114
rect 345756 339050 345808 339056
rect 345388 337952 345440 337958
rect 345388 337894 345440 337900
rect 345756 337952 345808 337958
rect 345756 337894 345808 337900
rect 345664 337204 345716 337210
rect 345664 337146 345716 337152
rect 345216 329038 345336 329066
rect 345308 328522 345336 329038
rect 345216 328494 345336 328522
rect 345216 318782 345244 328494
rect 345204 318776 345256 318782
rect 345204 318718 345256 318724
rect 345296 309188 345348 309194
rect 345216 309148 345296 309176
rect 345216 289814 345244 309148
rect 345296 309130 345348 309136
rect 345204 289808 345256 289814
rect 345204 289750 345256 289756
rect 345204 280288 345256 280294
rect 345204 280230 345256 280236
rect 345216 280140 345244 280230
rect 345216 280112 345336 280140
rect 345308 270586 345336 280112
rect 345216 270558 345336 270586
rect 345216 270502 345244 270558
rect 345204 270496 345256 270502
rect 345204 270438 345256 270444
rect 345204 260976 345256 260982
rect 345204 260918 345256 260924
rect 345216 260828 345244 260918
rect 345216 260800 345336 260828
rect 345308 251433 345336 260800
rect 345294 251424 345350 251433
rect 345294 251359 345350 251368
rect 345202 251288 345258 251297
rect 345202 251223 345258 251232
rect 345216 251190 345244 251223
rect 345204 251184 345256 251190
rect 345204 251126 345256 251132
rect 345216 241534 345244 241565
rect 345204 241528 345256 241534
rect 345256 241476 345428 241482
rect 345204 241470 345428 241476
rect 345216 241454 345428 241470
rect 345400 231946 345428 241454
rect 345388 231940 345440 231946
rect 345388 231882 345440 231888
rect 345296 231872 345348 231878
rect 345296 231814 345348 231820
rect 345216 222222 345244 222253
rect 345308 222222 345336 231814
rect 345204 222216 345256 222222
rect 345296 222216 345348 222222
rect 345256 222164 345296 222170
rect 345348 222164 345428 222170
rect 345204 222158 345428 222164
rect 345216 222142 345428 222158
rect 345400 212634 345428 222142
rect 345388 212628 345440 212634
rect 345388 212570 345440 212576
rect 345296 212560 345348 212566
rect 345296 212502 345348 212508
rect 345308 202892 345336 212502
rect 345216 202864 345336 202892
rect 345216 201482 345244 202864
rect 345204 201476 345256 201482
rect 345204 201418 345256 201424
rect 345112 193316 345164 193322
rect 345112 193258 345164 193264
rect 345112 193180 345164 193186
rect 345112 193122 345164 193128
rect 345020 192772 345072 192778
rect 345020 192714 345072 192720
rect 345032 190670 345060 192714
rect 345020 190664 345072 190670
rect 345020 190606 345072 190612
rect 345018 172544 345074 172553
rect 345018 172479 345074 172488
rect 345032 171086 345060 172479
rect 345020 171080 345072 171086
rect 345020 171022 345072 171028
rect 345124 4826 345152 193122
rect 345296 190664 345348 190670
rect 345296 190606 345348 190612
rect 345308 172553 345336 190606
rect 345294 172544 345350 172553
rect 345294 172479 345350 172488
rect 345204 171080 345256 171086
rect 345204 171022 345256 171028
rect 345216 162858 345244 171022
rect 345204 162852 345256 162858
rect 345204 162794 345256 162800
rect 345296 144968 345348 144974
rect 345216 144916 345296 144922
rect 345216 144910 345348 144916
rect 345216 144894 345336 144910
rect 345216 143546 345244 144894
rect 345204 143540 345256 143546
rect 345204 143482 345256 143488
rect 345388 143540 345440 143546
rect 345388 143482 345440 143488
rect 345400 125662 345428 143482
rect 345204 125656 345256 125662
rect 345204 125598 345256 125604
rect 345388 125656 345440 125662
rect 345388 125598 345440 125604
rect 345216 124166 345244 125598
rect 345204 124160 345256 124166
rect 345204 124102 345256 124108
rect 345204 114572 345256 114578
rect 345204 114514 345256 114520
rect 345216 104854 345244 114514
rect 345204 104848 345256 104854
rect 345204 104790 345256 104796
rect 345388 98728 345440 98734
rect 345388 98670 345440 98676
rect 345400 93838 345428 98670
rect 345388 93832 345440 93838
rect 345388 93774 345440 93780
rect 345204 75948 345256 75954
rect 345204 75890 345256 75896
rect 345216 66230 345244 75890
rect 345204 66224 345256 66230
rect 345204 66166 345256 66172
rect 345204 56636 345256 56642
rect 345204 56578 345256 56584
rect 345216 46918 345244 56578
rect 345204 46912 345256 46918
rect 345204 46854 345256 46860
rect 345296 29028 345348 29034
rect 345296 28970 345348 28976
rect 345308 27606 345336 28970
rect 345296 27600 345348 27606
rect 345296 27542 345348 27548
rect 345204 9716 345256 9722
rect 345204 9658 345256 9664
rect 345112 4820 345164 4826
rect 345112 4762 345164 4768
rect 345216 4146 345244 9658
rect 344928 4140 344980 4146
rect 344928 4082 344980 4088
rect 345204 4140 345256 4146
rect 345204 4082 345256 4088
rect 345480 4140 345532 4146
rect 345480 4082 345532 4088
rect 344376 4072 344428 4078
rect 344376 4014 344428 4020
rect 345492 480 345520 4082
rect 345676 2922 345704 337146
rect 345768 3058 345796 337894
rect 345952 335646 345980 340054
rect 346688 337142 346716 340068
rect 347148 337346 347176 340068
rect 347332 340054 347622 340082
rect 347136 337340 347188 337346
rect 347136 337282 347188 337288
rect 346676 337136 346728 337142
rect 346676 337078 346728 337084
rect 345940 335640 345992 335646
rect 345940 335582 345992 335588
rect 347332 328506 347360 340054
rect 348068 337006 348096 340068
rect 348252 340054 348542 340082
rect 348712 340054 349002 340082
rect 348252 338094 348280 340054
rect 348240 338088 348292 338094
rect 348240 338030 348292 338036
rect 348424 337544 348476 337550
rect 348424 337486 348476 337492
rect 348056 337000 348108 337006
rect 348056 336942 348108 336948
rect 347872 333328 347924 333334
rect 347872 333270 347924 333276
rect 346584 328500 346636 328506
rect 346584 328442 346636 328448
rect 347320 328500 347372 328506
rect 347320 328442 347372 328448
rect 346596 282962 346624 328442
rect 347780 289808 347832 289814
rect 347780 289750 347832 289756
rect 346504 282934 346624 282962
rect 346504 282826 346532 282934
rect 346504 282798 346624 282826
rect 346596 263650 346624 282798
rect 347792 280265 347820 289750
rect 347778 280256 347834 280265
rect 347778 280191 347834 280200
rect 346504 263622 346624 263650
rect 346504 263514 346532 263622
rect 346504 263486 346624 263514
rect 346596 244338 346624 263486
rect 346504 244310 346624 244338
rect 346504 244202 346532 244310
rect 346504 244174 346624 244202
rect 346596 225026 346624 244174
rect 346504 224998 346624 225026
rect 346504 224890 346532 224998
rect 346504 224862 346624 224890
rect 346596 205714 346624 224862
rect 346504 205686 346624 205714
rect 346504 205578 346532 205686
rect 346504 205550 346624 205578
rect 346596 186386 346624 205550
rect 346584 186380 346636 186386
rect 346584 186322 346636 186328
rect 346676 186244 346728 186250
rect 346676 186186 346728 186192
rect 346688 167074 346716 186186
rect 346492 167068 346544 167074
rect 346492 167010 346544 167016
rect 346676 167068 346728 167074
rect 346676 167010 346728 167016
rect 346504 166954 346532 167010
rect 346504 166926 346716 166954
rect 346688 135318 346716 166926
rect 346584 135312 346636 135318
rect 346584 135254 346636 135260
rect 346676 135312 346728 135318
rect 346676 135254 346728 135260
rect 346596 109154 346624 135254
rect 346504 109126 346624 109154
rect 346504 109018 346532 109126
rect 346504 108990 346624 109018
rect 346596 70514 346624 108990
rect 346584 70508 346636 70514
rect 346584 70450 346636 70456
rect 346584 70372 346636 70378
rect 346584 70314 346636 70320
rect 346596 51202 346624 70314
rect 346584 51196 346636 51202
rect 346584 51138 346636 51144
rect 346584 45620 346636 45626
rect 346584 45562 346636 45568
rect 346596 40746 346624 45562
rect 346504 40718 346624 40746
rect 346504 32450 346532 40718
rect 346504 32422 346624 32450
rect 346596 26246 346624 32422
rect 346584 26240 346636 26246
rect 346584 26182 346636 26188
rect 346400 16652 346452 16658
rect 346400 16594 346452 16600
rect 346412 4962 346440 16594
rect 346400 4956 346452 4962
rect 346400 4898 346452 4904
rect 347884 4894 347912 333270
rect 347964 328500 348016 328506
rect 347964 328442 348016 328448
rect 347976 328370 348004 328442
rect 347964 328364 348016 328370
rect 347964 328306 348016 328312
rect 347964 318844 348016 318850
rect 347964 318786 348016 318792
rect 347976 309330 348004 318786
rect 347964 309324 348016 309330
rect 347964 309266 348016 309272
rect 347964 309188 348016 309194
rect 347964 309130 348016 309136
rect 347976 309058 348004 309130
rect 347964 309052 348016 309058
rect 347964 308994 348016 309000
rect 347964 299600 348016 299606
rect 347964 299542 348016 299548
rect 347976 299470 348004 299542
rect 347964 299464 348016 299470
rect 347964 299406 348016 299412
rect 348056 299464 348108 299470
rect 348056 299406 348108 299412
rect 348068 289898 348096 299406
rect 347976 289870 348096 289898
rect 347976 289814 348004 289870
rect 347964 289808 348016 289814
rect 347964 289750 348016 289756
rect 347962 280256 348018 280265
rect 347962 280191 348018 280200
rect 347976 280158 348004 280191
rect 347964 280152 348016 280158
rect 347964 280094 348016 280100
rect 348056 280152 348108 280158
rect 348056 280094 348108 280100
rect 348068 270586 348096 280094
rect 347976 270558 348096 270586
rect 347976 270502 348004 270558
rect 347964 270496 348016 270502
rect 347964 270438 348016 270444
rect 347964 260976 348016 260982
rect 347964 260918 348016 260924
rect 347976 260846 348004 260918
rect 347964 260840 348016 260846
rect 347964 260782 348016 260788
rect 348056 260772 348108 260778
rect 348056 260714 348108 260720
rect 348068 251274 348096 260714
rect 347976 251246 348096 251274
rect 347976 251190 348004 251246
rect 347964 251184 348016 251190
rect 347964 251126 348016 251132
rect 347964 241528 348016 241534
rect 347964 241470 348016 241476
rect 347976 231849 348004 241470
rect 347962 231840 348018 231849
rect 347962 231775 348018 231784
rect 348146 231840 348202 231849
rect 348146 231775 348202 231784
rect 348160 222222 348188 231775
rect 347964 222216 348016 222222
rect 347964 222158 348016 222164
rect 348148 222216 348200 222222
rect 348148 222158 348200 222164
rect 347976 212537 348004 222158
rect 347962 212528 348018 212537
rect 347962 212463 348018 212472
rect 348146 212528 348202 212537
rect 348146 212463 348202 212472
rect 348160 202910 348188 212463
rect 347964 202904 348016 202910
rect 347964 202846 348016 202852
rect 348148 202904 348200 202910
rect 348148 202846 348200 202852
rect 347976 193225 348004 202846
rect 347962 193216 348018 193225
rect 347962 193151 348018 193160
rect 348146 193216 348202 193225
rect 348146 193151 348202 193160
rect 348160 183598 348188 193151
rect 347964 183592 348016 183598
rect 347964 183534 348016 183540
rect 348148 183592 348200 183598
rect 348148 183534 348200 183540
rect 347976 173913 348004 183534
rect 347962 173904 348018 173913
rect 347962 173839 348018 173848
rect 348146 173904 348202 173913
rect 348146 173839 348202 173848
rect 348160 164257 348188 173839
rect 347962 164248 348018 164257
rect 347962 164183 348018 164192
rect 348146 164248 348202 164257
rect 348146 164183 348202 164192
rect 347976 154562 348004 164183
rect 347964 154556 348016 154562
rect 347964 154498 348016 154504
rect 348148 154556 348200 154562
rect 348148 154498 348200 154504
rect 348160 144945 348188 154498
rect 347962 144936 348018 144945
rect 347962 144871 348018 144880
rect 348146 144936 348202 144945
rect 348146 144871 348202 144880
rect 347976 135250 348004 144871
rect 347964 135244 348016 135250
rect 347964 135186 348016 135192
rect 348148 135244 348200 135250
rect 348148 135186 348200 135192
rect 348160 125633 348188 135186
rect 347962 125624 348018 125633
rect 347962 125559 347964 125568
rect 348016 125559 348018 125568
rect 348146 125624 348202 125633
rect 348146 125559 348202 125568
rect 347964 125530 348016 125536
rect 347964 116068 348016 116074
rect 347964 116010 348016 116016
rect 347976 115938 348004 116010
rect 347964 115932 348016 115938
rect 347964 115874 348016 115880
rect 348148 115932 348200 115938
rect 348148 115874 348200 115880
rect 348160 106321 348188 115874
rect 347962 106312 348018 106321
rect 347962 106247 347964 106256
rect 348016 106247 348018 106256
rect 348146 106312 348202 106321
rect 348146 106247 348202 106256
rect 347964 106218 348016 106224
rect 347964 96756 348016 96762
rect 347964 96698 348016 96704
rect 347976 96626 348004 96698
rect 347964 96620 348016 96626
rect 347964 96562 348016 96568
rect 348056 96620 348108 96626
rect 348056 96562 348108 96568
rect 348068 89706 348096 96562
rect 347976 89678 348096 89706
rect 347976 86986 348004 89678
rect 347976 86958 348096 86986
rect 348068 80186 348096 86958
rect 348068 80158 348188 80186
rect 348160 74610 348188 80158
rect 348068 74582 348188 74610
rect 348068 74526 348096 74582
rect 348056 74520 348108 74526
rect 348056 74462 348108 74468
rect 347964 64932 348016 64938
rect 347964 64874 348016 64880
rect 347976 55214 348004 64874
rect 348330 64016 348386 64025
rect 348330 63951 348386 63960
rect 348344 63753 348372 63951
rect 348330 63744 348386 63753
rect 348330 63679 348386 63688
rect 347964 55208 348016 55214
rect 347964 55150 348016 55156
rect 347964 45688 348016 45694
rect 347964 45630 348016 45636
rect 347976 45529 348004 45630
rect 347962 45520 348018 45529
rect 347962 45455 348018 45464
rect 348054 45384 348110 45393
rect 348054 45319 348110 45328
rect 348068 26217 348096 45319
rect 348054 26208 348110 26217
rect 348054 26143 348110 26152
rect 348238 26208 348294 26217
rect 348238 26143 348294 26152
rect 348252 24857 348280 26143
rect 348054 24848 348110 24857
rect 348054 24783 348110 24792
rect 348238 24848 348294 24857
rect 348238 24783 348294 24792
rect 348068 16266 348096 24783
rect 348068 16238 348280 16266
rect 348252 6934 348280 16238
rect 348056 6928 348108 6934
rect 348056 6870 348108 6876
rect 348240 6928 348292 6934
rect 348240 6870 348292 6876
rect 347872 4888 347924 4894
rect 347872 4830 347924 4836
rect 346676 4072 346728 4078
rect 346676 4014 346728 4020
rect 345756 3052 345808 3058
rect 345756 2994 345808 3000
rect 345664 2916 345716 2922
rect 345664 2858 345716 2864
rect 346688 480 346716 4014
rect 347872 3596 347924 3602
rect 347872 3538 347924 3544
rect 347884 480 347912 3538
rect 348068 3466 348096 6870
rect 348056 3460 348108 3466
rect 348056 3402 348108 3408
rect 348436 3262 348464 337486
rect 348712 333334 348740 340054
rect 349068 338020 349120 338026
rect 349068 337962 349120 337968
rect 348700 333328 348752 333334
rect 348700 333270 348752 333276
rect 349080 3602 349108 337962
rect 349356 336870 349384 340068
rect 349448 340054 349830 340082
rect 349448 337890 349476 340054
rect 349804 338088 349856 338094
rect 349804 338030 349856 338036
rect 349436 337884 349488 337890
rect 349436 337826 349488 337832
rect 349344 336864 349396 336870
rect 349344 336806 349396 336812
rect 349816 4146 349844 338030
rect 350276 336938 350304 340068
rect 350736 337278 350764 340068
rect 350828 340054 351210 340082
rect 350724 337272 350776 337278
rect 350724 337214 350776 337220
rect 350264 336932 350316 336938
rect 350264 336874 350316 336880
rect 349804 4140 349856 4146
rect 349804 4082 349856 4088
rect 350828 3806 350856 340054
rect 351656 337958 351684 340068
rect 351644 337952 351696 337958
rect 351644 337894 351696 337900
rect 351828 337952 351880 337958
rect 351828 337894 351880 337900
rect 351184 337340 351236 337346
rect 351184 337282 351236 337288
rect 350816 3800 350868 3806
rect 350816 3742 350868 3748
rect 349068 3596 349120 3602
rect 349068 3538 349120 3544
rect 350264 3460 350316 3466
rect 350264 3402 350316 3408
rect 349068 3324 349120 3330
rect 349068 3266 349120 3272
rect 348424 3256 348476 3262
rect 348424 3198 348476 3204
rect 349080 480 349108 3266
rect 350276 480 350304 3402
rect 351196 3330 351224 337282
rect 351840 3534 351868 337894
rect 352012 337884 352064 337890
rect 352012 337826 352064 337832
rect 352024 4010 352052 337826
rect 352012 4004 352064 4010
rect 352012 3946 352064 3952
rect 352116 3942 352144 340068
rect 352208 340054 352590 340082
rect 352760 340054 353050 340082
rect 352208 337414 352236 340054
rect 352760 337890 352788 340054
rect 352748 337884 352800 337890
rect 352748 337826 352800 337832
rect 353404 337754 353432 340068
rect 352564 337748 352616 337754
rect 352564 337690 352616 337696
rect 353392 337748 353444 337754
rect 353392 337690 353444 337696
rect 352196 337408 352248 337414
rect 352196 337350 352248 337356
rect 352104 3936 352156 3942
rect 352104 3878 352156 3884
rect 352576 3618 352604 337690
rect 353208 337544 353260 337550
rect 353208 337486 353260 337492
rect 352484 3590 352604 3618
rect 351368 3528 351420 3534
rect 351368 3470 351420 3476
rect 351828 3528 351880 3534
rect 351828 3470 351880 3476
rect 351184 3324 351236 3330
rect 351184 3266 351236 3272
rect 351380 480 351408 3470
rect 352484 3194 352512 3590
rect 353220 3534 353248 337486
rect 353864 337074 353892 340068
rect 353852 337068 353904 337074
rect 353852 337010 353904 337016
rect 354324 336802 354352 340068
rect 354784 337210 354812 340068
rect 354876 340054 355258 340082
rect 354772 337204 354824 337210
rect 354772 337146 354824 337152
rect 354312 336796 354364 336802
rect 354312 336738 354364 336744
rect 353760 3596 353812 3602
rect 353760 3538 353812 3544
rect 352564 3528 352616 3534
rect 352564 3470 352616 3476
rect 353208 3528 353260 3534
rect 353208 3470 353260 3476
rect 352472 3188 352524 3194
rect 352472 3130 352524 3136
rect 352576 480 352604 3470
rect 353772 480 353800 3538
rect 354876 3398 354904 340054
rect 355324 337884 355376 337890
rect 355324 337826 355376 337832
rect 355336 4146 355364 337826
rect 355704 337482 355732 340068
rect 356178 340054 356468 340082
rect 355692 337476 355744 337482
rect 355692 337418 355744 337424
rect 355968 337408 356020 337414
rect 355968 337350 356020 337356
rect 355324 4140 355376 4146
rect 355324 4082 355376 4088
rect 355980 3534 356008 337350
rect 356060 87168 356112 87174
rect 356058 87136 356060 87145
rect 356112 87136 356114 87145
rect 356058 87071 356114 87080
rect 356058 40216 356114 40225
rect 356058 40151 356114 40160
rect 356072 40118 356100 40151
rect 356060 40112 356112 40118
rect 356060 40054 356112 40060
rect 354956 3528 355008 3534
rect 354956 3470 355008 3476
rect 355968 3528 356020 3534
rect 355968 3470 356020 3476
rect 354864 3392 354916 3398
rect 354864 3334 354916 3340
rect 354968 480 354996 3470
rect 356152 3324 356204 3330
rect 356152 3266 356204 3272
rect 356164 480 356192 3266
rect 356440 2990 356468 340054
rect 356532 340054 356638 340082
rect 356428 2984 356480 2990
rect 356428 2926 356480 2932
rect 356532 2854 356560 340054
rect 356704 337748 356756 337754
rect 356704 337690 356756 337696
rect 356716 4078 356744 337690
rect 356992 337618 357020 340068
rect 357452 338094 357480 340068
rect 357636 340054 357926 340082
rect 357440 338088 357492 338094
rect 357440 338030 357492 338036
rect 356980 337612 357032 337618
rect 356980 337554 357032 337560
rect 357440 134088 357492 134094
rect 357438 134056 357440 134065
rect 357492 134056 357494 134065
rect 357438 133991 357494 134000
rect 356704 4072 356756 4078
rect 356704 4014 356756 4020
rect 357636 3738 357664 340054
rect 358372 337686 358400 340068
rect 358360 337680 358412 337686
rect 358360 337622 358412 337628
rect 358084 337612 358136 337618
rect 358084 337554 358136 337560
rect 357624 3732 357676 3738
rect 357624 3674 357676 3680
rect 358096 3602 358124 337554
rect 358728 337136 358780 337142
rect 358728 337078 358780 337084
rect 358084 3596 358136 3602
rect 358084 3538 358136 3544
rect 357348 3120 357400 3126
rect 357348 3062 357400 3068
rect 356520 2848 356572 2854
rect 356520 2790 356572 2796
rect 357360 480 357388 3062
rect 358740 610 358768 337078
rect 358832 3670 358860 340068
rect 359292 337890 359320 340068
rect 359280 337884 359332 337890
rect 359280 337826 359332 337832
rect 359752 337822 359780 340068
rect 360212 338026 360240 340068
rect 360200 338020 360252 338026
rect 360200 337962 360252 337968
rect 359740 337816 359792 337822
rect 359740 337758 359792 337764
rect 360580 337754 360608 340068
rect 361040 337958 361068 340068
rect 361028 337952 361080 337958
rect 361028 337894 361080 337900
rect 360568 337748 360620 337754
rect 360568 337690 360620 337696
rect 361500 337346 361528 340068
rect 361776 340054 361974 340082
rect 363052 340070 363104 340076
rect 363880 340128 363932 340134
rect 363880 340070 363932 340076
rect 361488 337340 361540 337346
rect 361488 337282 361540 337288
rect 359464 337068 359516 337074
rect 359464 337010 359516 337016
rect 358820 3664 358872 3670
rect 358820 3606 358872 3612
rect 359476 3126 359504 337010
rect 360108 337000 360160 337006
rect 360108 336942 360160 336948
rect 359554 63744 359610 63753
rect 359554 63679 359556 63688
rect 359608 63679 359610 63688
rect 359556 63650 359608 63656
rect 360014 16824 360070 16833
rect 360014 16759 360016 16768
rect 360068 16759 360070 16768
rect 360016 16730 360068 16736
rect 359464 3120 359516 3126
rect 359464 3062 359516 3068
rect 360120 626 360148 336942
rect 361120 134088 361172 134094
rect 361118 134056 361120 134065
rect 361172 134056 361174 134065
rect 361118 133991 361174 134000
rect 361118 16824 361174 16833
rect 361118 16759 361120 16768
rect 361172 16759 361174 16768
rect 361120 16730 361172 16736
rect 360936 4004 360988 4010
rect 360936 3946 360988 3952
rect 358544 604 358596 610
rect 358544 546 358596 552
rect 358728 604 358780 610
rect 358728 546 358780 552
rect 359752 598 360148 626
rect 358556 480 358584 546
rect 359752 480 359780 598
rect 360948 480 360976 3946
rect 361776 3534 361804 340054
rect 362420 337550 362448 340068
rect 362408 337544 362460 337550
rect 362408 337486 362460 337492
rect 362880 337482 362908 340068
rect 363064 338094 363092 340070
rect 363052 338088 363104 338094
rect 363052 338030 363104 338036
rect 363144 338088 363196 338094
rect 363144 338030 363196 338036
rect 362868 337476 362920 337482
rect 362868 337418 362920 337424
rect 363156 337396 363184 338030
rect 363340 337618 363368 340068
rect 363328 337612 363380 337618
rect 363328 337554 363380 337560
rect 363800 337414 363828 340068
rect 363788 337408 363840 337414
rect 363156 337368 363276 337396
rect 362224 336864 362276 336870
rect 362224 336806 362276 336812
rect 362130 181520 362186 181529
rect 362130 181455 362186 181464
rect 362144 180849 362172 181455
rect 362130 180840 362186 180849
rect 362130 180775 362186 180784
rect 362132 4140 362184 4146
rect 362132 4082 362184 4088
rect 361764 3528 361816 3534
rect 361764 3470 361816 3476
rect 362144 480 362172 4082
rect 362236 4010 362264 336806
rect 362868 336796 362920 336802
rect 362868 336738 362920 336744
rect 362880 4146 362908 336738
rect 363248 328438 363276 337368
rect 363788 337350 363840 337356
rect 364628 337074 364656 340068
rect 365088 337142 365116 340068
rect 365548 337210 365576 340068
rect 365536 337204 365588 337210
rect 365536 337146 365588 337152
rect 365076 337136 365128 337142
rect 365076 337078 365128 337084
rect 364616 337068 364668 337074
rect 364616 337010 364668 337016
rect 364248 337000 364300 337006
rect 364248 336942 364300 336948
rect 363236 328432 363288 328438
rect 363236 328374 363288 328380
rect 363328 318844 363380 318850
rect 363328 318786 363380 318792
rect 363340 309194 363368 318786
rect 362960 309188 363012 309194
rect 362960 309130 363012 309136
rect 363328 309188 363380 309194
rect 363328 309130 363380 309136
rect 362972 302122 363000 309130
rect 362960 302116 363012 302122
rect 362960 302058 363012 302064
rect 363236 302116 363288 302122
rect 363236 302058 363288 302064
rect 363248 285002 363276 302058
rect 363156 284974 363276 285002
rect 363156 280158 363184 284974
rect 363144 280152 363196 280158
rect 363144 280094 363196 280100
rect 363236 270564 363288 270570
rect 363236 270506 363288 270512
rect 363248 263514 363276 270506
rect 363156 263486 363276 263514
rect 363156 260846 363184 263486
rect 363144 260840 363196 260846
rect 363144 260782 363196 260788
rect 363236 251252 363288 251258
rect 363236 251194 363288 251200
rect 363248 244202 363276 251194
rect 363156 244174 363276 244202
rect 363156 241505 363184 244174
rect 362958 241496 363014 241505
rect 362958 241431 363014 241440
rect 363142 241496 363198 241505
rect 363142 241431 363198 241440
rect 362972 231878 363000 241431
rect 362960 231872 363012 231878
rect 362960 231814 363012 231820
rect 363236 231872 363288 231878
rect 363236 231814 363288 231820
rect 363248 224890 363276 231814
rect 363156 224862 363276 224890
rect 363156 222193 363184 224862
rect 362958 222184 363014 222193
rect 362958 222119 363014 222128
rect 363142 222184 363198 222193
rect 363142 222119 363198 222128
rect 362972 212566 363000 222119
rect 362960 212560 363012 212566
rect 362960 212502 363012 212508
rect 363236 212560 363288 212566
rect 363236 212502 363288 212508
rect 363248 205578 363276 212502
rect 363156 205550 363276 205578
rect 363156 202881 363184 205550
rect 362958 202872 363014 202881
rect 362958 202807 363014 202816
rect 363142 202872 363198 202881
rect 363142 202807 363198 202816
rect 362972 193254 363000 202807
rect 362960 193248 363012 193254
rect 362960 193190 363012 193196
rect 363236 193248 363288 193254
rect 363236 193190 363288 193196
rect 363248 186266 363276 193190
rect 363156 186238 363276 186266
rect 363156 183569 363184 186238
rect 362958 183560 363014 183569
rect 362958 183495 363014 183504
rect 363142 183560 363198 183569
rect 363142 183495 363198 183504
rect 362972 173942 363000 183495
rect 362960 173936 363012 173942
rect 362960 173878 363012 173884
rect 363236 173936 363288 173942
rect 363236 173878 363288 173884
rect 363248 166954 363276 173878
rect 363156 166926 363276 166954
rect 363156 164218 363184 166926
rect 362960 164212 363012 164218
rect 362960 164154 363012 164160
rect 363144 164212 363196 164218
rect 363144 164154 363196 164160
rect 362972 154601 363000 164154
rect 362958 154592 363014 154601
rect 362958 154527 363014 154536
rect 363234 154592 363290 154601
rect 363234 154527 363290 154536
rect 363248 147642 363276 154527
rect 363156 147614 363276 147642
rect 363156 140026 363184 147614
rect 362972 139998 363184 140026
rect 362972 135289 363000 139998
rect 362958 135280 363014 135289
rect 362958 135215 363014 135224
rect 363234 135280 363290 135289
rect 363234 135215 363290 135224
rect 363248 128330 363276 135215
rect 363156 128302 363276 128330
rect 363156 120714 363184 128302
rect 362972 120686 363184 120714
rect 362972 115977 363000 120686
rect 362958 115968 363014 115977
rect 362958 115903 363014 115912
rect 363234 115968 363290 115977
rect 363234 115903 363290 115912
rect 363248 109018 363276 115903
rect 363156 108990 363276 109018
rect 363156 101402 363184 108990
rect 362972 101374 363184 101402
rect 362972 96665 363000 101374
rect 362958 96656 363014 96665
rect 362958 96591 363014 96600
rect 363234 96656 363290 96665
rect 363234 96591 363290 96600
rect 363248 89706 363276 96591
rect 363064 89678 363276 89706
rect 363064 86970 363092 89678
rect 363052 86964 363104 86970
rect 363052 86906 363104 86912
rect 362960 77308 363012 77314
rect 362960 77250 363012 77256
rect 362972 77178 363000 77250
rect 362960 77172 363012 77178
rect 362960 77114 363012 77120
rect 363052 70304 363104 70310
rect 363052 70246 363104 70252
rect 363064 60722 363092 70246
rect 363052 60716 363104 60722
rect 363052 60658 363104 60664
rect 363236 60716 363288 60722
rect 363236 60658 363288 60664
rect 363248 57934 363276 60658
rect 363236 57928 363288 57934
rect 363236 57870 363288 57876
rect 363144 48340 363196 48346
rect 363144 48282 363196 48288
rect 363156 41426 363184 48282
rect 363064 41410 363184 41426
rect 363052 41404 363184 41410
rect 363104 41398 363184 41404
rect 363236 41404 363288 41410
rect 363052 41346 363104 41352
rect 363236 41346 363288 41352
rect 363248 38622 363276 41346
rect 363236 38616 363288 38622
rect 363236 38558 363288 38564
rect 363144 29028 363196 29034
rect 363144 28970 363196 28976
rect 363156 22114 363184 28970
rect 363064 22098 363184 22114
rect 363052 22092 363184 22098
rect 363104 22086 363184 22092
rect 363236 22092 363288 22098
rect 363052 22034 363104 22040
rect 363236 22034 363288 22040
rect 363248 19310 363276 22034
rect 363236 19304 363288 19310
rect 363236 19246 363288 19252
rect 363236 9716 363288 9722
rect 363236 9658 363288 9664
rect 362868 4140 362920 4146
rect 362868 4082 362920 4088
rect 362224 4004 362276 4010
rect 362224 3946 362276 3952
rect 363248 3330 363276 9658
rect 364260 3534 364288 336942
rect 366008 336870 366036 340068
rect 366364 336932 366416 336938
rect 366364 336874 366416 336880
rect 365996 336864 366048 336870
rect 365996 336806 366048 336812
rect 365626 87408 365682 87417
rect 365626 87343 365682 87352
rect 365640 87174 365668 87343
rect 365628 87168 365680 87174
rect 365628 87110 365680 87116
rect 365628 63708 365680 63714
rect 365628 63650 365680 63656
rect 365640 63617 365668 63650
rect 365626 63608 365682 63617
rect 365626 63543 365682 63552
rect 365628 40112 365680 40118
rect 365626 40080 365628 40089
rect 365680 40080 365682 40089
rect 365626 40015 365682 40024
rect 366376 4146 366404 336874
rect 366468 336802 366496 340068
rect 366928 337006 366956 340068
rect 366916 337000 366968 337006
rect 366916 336942 366968 336948
rect 367388 336938 367416 340068
rect 367376 336932 367428 336938
rect 367376 336874 367428 336880
rect 367848 336870 367876 340068
rect 366916 336864 366968 336870
rect 366916 336806 366968 336812
rect 367836 336864 367888 336870
rect 367836 336806 367888 336812
rect 366456 336796 366508 336802
rect 366456 336738 366508 336744
rect 364524 4140 364576 4146
rect 364524 4082 364576 4088
rect 366364 4140 366416 4146
rect 366364 4082 366416 4088
rect 363328 3528 363380 3534
rect 363328 3470 363380 3476
rect 364248 3528 364300 3534
rect 364248 3470 364300 3476
rect 363236 3324 363288 3330
rect 363236 3266 363288 3272
rect 363340 480 363368 3470
rect 364536 480 364564 4082
rect 366928 3330 366956 336806
rect 368216 336802 368244 340068
rect 368492 340054 368690 340082
rect 368860 340054 369150 340082
rect 369610 340054 369808 340082
rect 367008 336796 367060 336802
rect 367008 336738 367060 336744
rect 368204 336796 368256 336802
rect 368204 336738 368256 336744
rect 365720 3324 365772 3330
rect 365720 3266 365772 3272
rect 366916 3324 366968 3330
rect 366916 3266 366968 3272
rect 365732 480 365760 3266
rect 367020 3210 367048 336738
rect 368492 4146 368520 340054
rect 368860 335594 368888 340054
rect 369780 337770 369808 340054
rect 370056 337890 370084 340068
rect 370044 337884 370096 337890
rect 370044 337826 370096 337832
rect 369780 337742 370084 337770
rect 368584 335566 368888 335594
rect 368584 4146 368612 335566
rect 368020 4140 368072 4146
rect 368020 4082 368072 4088
rect 368480 4140 368532 4146
rect 368480 4082 368532 4088
rect 368572 4140 368624 4146
rect 368572 4082 368624 4088
rect 369216 4140 369268 4146
rect 369216 4082 369268 4088
rect 366928 3182 367048 3210
rect 366928 480 366956 3182
rect 368032 480 368060 4082
rect 369228 480 369256 4082
rect 370056 3346 370084 337742
rect 370516 337210 370544 340068
rect 370990 340054 371188 340082
rect 371056 337884 371108 337890
rect 371056 337826 371108 337832
rect 370504 337204 370556 337210
rect 370504 337146 370556 337152
rect 371068 3534 371096 337826
rect 371160 4146 371188 340054
rect 371436 337550 371464 340068
rect 371424 337544 371476 337550
rect 371424 337486 371476 337492
rect 371804 337074 371832 340068
rect 372264 337754 372292 340068
rect 372252 337748 372304 337754
rect 372252 337690 372304 337696
rect 372724 337686 372752 340068
rect 372712 337680 372764 337686
rect 372712 337622 372764 337628
rect 373184 337482 373212 340068
rect 373264 337748 373316 337754
rect 373264 337690 373316 337696
rect 373172 337476 373224 337482
rect 373172 337418 373224 337424
rect 372712 337204 372764 337210
rect 372712 337146 372764 337152
rect 371792 337068 371844 337074
rect 371792 337010 371844 337016
rect 371148 4140 371200 4146
rect 371148 4082 371200 4088
rect 371056 3528 371108 3534
rect 371056 3470 371108 3476
rect 371608 3528 371660 3534
rect 371608 3470 371660 3476
rect 372724 3482 372752 337146
rect 373276 3534 373304 337690
rect 373644 336938 373672 340068
rect 374104 337754 374132 340068
rect 374564 337822 374592 340068
rect 374552 337816 374604 337822
rect 374552 337758 374604 337764
rect 374092 337748 374144 337754
rect 374092 337690 374144 337696
rect 373908 337680 373960 337686
rect 373908 337622 373960 337628
rect 373632 336932 373684 336938
rect 373632 336874 373684 336880
rect 373264 3528 373316 3534
rect 370056 3318 370452 3346
rect 370424 480 370452 3318
rect 371620 480 371648 3470
rect 372724 3454 372844 3482
rect 373264 3470 373316 3476
rect 373920 3466 373948 337622
rect 374092 337544 374144 337550
rect 374092 337486 374144 337492
rect 374000 4140 374052 4146
rect 374000 4082 374052 4088
rect 372816 480 372844 3454
rect 373908 3460 373960 3466
rect 373908 3402 373960 3408
rect 374012 480 374040 4082
rect 374104 3346 374132 337486
rect 375024 337346 375052 340068
rect 375288 337748 375340 337754
rect 375288 337690 375340 337696
rect 375012 337340 375064 337346
rect 375012 337282 375064 337288
rect 374644 336932 374696 336938
rect 374644 336874 374696 336880
rect 374656 3806 374684 336874
rect 374644 3800 374696 3806
rect 374644 3742 374696 3748
rect 374104 3318 375236 3346
rect 375300 3330 375328 337690
rect 375392 337618 375420 340068
rect 375852 337686 375880 340068
rect 376312 338026 376340 340068
rect 376300 338020 376352 338026
rect 376300 337962 376352 337968
rect 376024 337816 376076 337822
rect 376024 337758 376076 337764
rect 375840 337680 375892 337686
rect 375840 337622 375892 337628
rect 375380 337612 375432 337618
rect 375380 337554 375432 337560
rect 375656 337068 375708 337074
rect 375656 337010 375708 337016
rect 375668 3346 375696 337010
rect 376036 3874 376064 337758
rect 376668 337612 376720 337618
rect 376668 337554 376720 337560
rect 376024 3868 376076 3874
rect 376024 3810 376076 3816
rect 376680 3738 376708 337554
rect 376772 337482 376800 340068
rect 377232 337754 377260 340068
rect 377692 338094 377720 340068
rect 377680 338088 377732 338094
rect 377680 338030 377732 338036
rect 377220 337748 377272 337754
rect 377220 337690 377272 337696
rect 377956 337748 378008 337754
rect 377956 337690 378008 337696
rect 377404 337680 377456 337686
rect 377404 337622 377456 337628
rect 376760 337476 376812 337482
rect 376760 337418 376812 337424
rect 376668 3732 376720 3738
rect 376668 3674 376720 3680
rect 377416 3670 377444 337622
rect 377404 3664 377456 3670
rect 377404 3606 377456 3612
rect 377968 3534 377996 337690
rect 378152 337550 378180 340068
rect 378612 337686 378640 340068
rect 378600 337680 378652 337686
rect 378600 337622 378652 337628
rect 379072 337618 379100 340068
rect 379440 337958 379468 340068
rect 379428 337952 379480 337958
rect 379428 337894 379480 337900
rect 379900 337754 379928 340068
rect 379888 337748 379940 337754
rect 379888 337690 379940 337696
rect 380360 337686 380388 340068
rect 380820 337890 380848 340068
rect 380808 337884 380860 337890
rect 380808 337826 380860 337832
rect 381280 337754 381308 340068
rect 380808 337748 380860 337754
rect 380808 337690 380860 337696
rect 381268 337748 381320 337754
rect 381268 337690 381320 337696
rect 380164 337680 380216 337686
rect 380164 337622 380216 337628
rect 380348 337680 380400 337686
rect 380348 337622 380400 337628
rect 379060 337612 379112 337618
rect 379060 337554 379112 337560
rect 378140 337544 378192 337550
rect 378140 337486 378192 337492
rect 378048 337476 378100 337482
rect 378048 337418 378100 337424
rect 378060 3602 378088 337418
rect 379612 337408 379664 337414
rect 379612 337350 379664 337356
rect 378048 3596 378100 3602
rect 378048 3538 378100 3544
rect 377588 3528 377640 3534
rect 377588 3470 377640 3476
rect 377956 3528 378008 3534
rect 377956 3470 378008 3476
rect 375208 480 375236 3318
rect 375288 3324 375340 3330
rect 375668 3318 376432 3346
rect 375288 3266 375340 3272
rect 376404 480 376432 3318
rect 377600 480 377628 3470
rect 378784 3460 378836 3466
rect 378784 3402 378836 3408
rect 378796 480 378824 3402
rect 379624 610 379652 337350
rect 380176 3466 380204 337622
rect 380164 3460 380216 3466
rect 380164 3402 380216 3408
rect 380820 3058 380848 337690
rect 381636 337612 381688 337618
rect 381636 337554 381688 337560
rect 381544 337340 381596 337346
rect 381544 337282 381596 337288
rect 381556 4146 381584 337282
rect 381544 4140 381596 4146
rect 381544 4082 381596 4088
rect 381176 3800 381228 3806
rect 381176 3742 381228 3748
rect 380808 3052 380860 3058
rect 380808 2994 380860 3000
rect 379612 604 379664 610
rect 379612 546 379664 552
rect 379980 604 380032 610
rect 379980 546 380032 552
rect 379992 480 380020 546
rect 381188 480 381216 3742
rect 381648 2990 381676 337554
rect 381740 337482 381768 340068
rect 382108 340054 382214 340082
rect 381728 337476 381780 337482
rect 381728 337418 381780 337424
rect 382108 3194 382136 340054
rect 382660 337822 382688 340068
rect 382648 337816 382700 337822
rect 382648 337758 382700 337764
rect 382188 337748 382240 337754
rect 382188 337690 382240 337696
rect 382096 3188 382148 3194
rect 382096 3130 382148 3136
rect 382200 3126 382228 337690
rect 383028 337414 383056 340068
rect 383502 340054 383608 340082
rect 383016 337408 383068 337414
rect 383016 337350 383068 337356
rect 383476 3868 383528 3874
rect 383476 3810 383528 3816
rect 382372 3324 382424 3330
rect 382372 3266 382424 3272
rect 382188 3120 382240 3126
rect 382188 3062 382240 3068
rect 381636 2984 381688 2990
rect 381636 2926 381688 2932
rect 382384 480 382412 3266
rect 383488 3210 383516 3810
rect 383580 3330 383608 340054
rect 383948 337754 383976 340068
rect 384776 337770 384804 340190
rect 384868 338094 384896 340068
rect 384856 338088 384908 338094
rect 384856 338030 384908 338036
rect 383936 337748 383988 337754
rect 384776 337742 384896 337770
rect 383936 337690 383988 337696
rect 384304 337544 384356 337550
rect 384304 337486 384356 337492
rect 383568 3324 383620 3330
rect 383568 3266 383620 3272
rect 384316 3262 384344 337486
rect 384672 4140 384724 4146
rect 384672 4082 384724 4088
rect 384304 3256 384356 3262
rect 383488 3182 383608 3210
rect 384304 3198 384356 3204
rect 383580 480 383608 3182
rect 384684 480 384712 4082
rect 384868 3806 384896 337742
rect 384948 337748 385000 337754
rect 384948 337690 385000 337696
rect 384960 3942 384988 337690
rect 385328 337346 385356 340068
rect 385802 340054 386092 340082
rect 386262 340054 386368 340082
rect 386064 337770 386092 340054
rect 386064 337742 386276 337770
rect 385316 337340 385368 337346
rect 385316 337282 385368 337288
rect 386248 4622 386276 337742
rect 386236 4616 386288 4622
rect 386236 4558 386288 4564
rect 384948 3936 385000 3942
rect 384948 3878 385000 3884
rect 384856 3800 384908 3806
rect 384856 3742 384908 3748
rect 386340 3738 386368 340054
rect 386616 337618 386644 340068
rect 387090 340054 387472 340082
rect 387550 340054 387748 340082
rect 387444 337770 387472 340054
rect 387444 337742 387656 337770
rect 386604 337612 386656 337618
rect 386604 337554 386656 337560
rect 387524 337612 387576 337618
rect 387524 337554 387576 337560
rect 387064 337544 387116 337550
rect 387064 337486 387116 337492
rect 387076 3874 387104 337486
rect 387536 4690 387564 337554
rect 387524 4684 387576 4690
rect 387524 4626 387576 4632
rect 387628 4078 387656 337742
rect 387720 4146 387748 340054
rect 387996 337550 388024 340068
rect 388444 337884 388496 337890
rect 388444 337826 388496 337832
rect 387984 337544 388036 337550
rect 387984 337486 388036 337492
rect 387708 4140 387760 4146
rect 387708 4082 387760 4088
rect 387616 4072 387668 4078
rect 387616 4014 387668 4020
rect 387064 3868 387116 3874
rect 387064 3810 387116 3816
rect 385868 3732 385920 3738
rect 385868 3674 385920 3680
rect 386328 3732 386380 3738
rect 386328 3674 386380 3680
rect 385880 480 385908 3674
rect 387064 3664 387116 3670
rect 387064 3606 387116 3612
rect 387076 480 387104 3606
rect 388456 3534 388484 337826
rect 388824 337770 388852 340190
rect 388930 340054 389128 340082
rect 388824 337742 389036 337770
rect 389008 3942 389036 337742
rect 389100 4010 389128 340054
rect 389376 337754 389404 340068
rect 389364 337748 389416 337754
rect 389364 337690 389416 337696
rect 389836 337074 389864 340068
rect 390296 338026 390324 340068
rect 390284 338020 390336 338026
rect 390284 337962 390336 337968
rect 390468 337748 390520 337754
rect 390468 337690 390520 337696
rect 389824 337068 389876 337074
rect 389824 337010 389876 337016
rect 390376 337068 390428 337074
rect 390376 337010 390428 337016
rect 390388 5506 390416 337010
rect 390376 5500 390428 5506
rect 390376 5442 390428 5448
rect 390480 4758 390508 337690
rect 390664 337618 390692 340068
rect 391138 340054 391520 340082
rect 391598 340054 391888 340082
rect 391492 337770 391520 340054
rect 391492 337742 391796 337770
rect 390652 337612 390704 337618
rect 390652 337554 390704 337560
rect 391664 337612 391716 337618
rect 391664 337554 391716 337560
rect 391480 8220 391532 8226
rect 391480 8162 391532 8168
rect 390468 4752 390520 4758
rect 390468 4694 390520 4700
rect 389088 4004 389140 4010
rect 389088 3946 389140 3952
rect 388996 3936 389048 3942
rect 388996 3878 389048 3884
rect 389456 3596 389508 3602
rect 389456 3538 389508 3544
rect 388444 3528 388496 3534
rect 388444 3470 388496 3476
rect 388260 3256 388312 3262
rect 388260 3198 388312 3204
rect 388272 480 388300 3198
rect 389468 480 389496 3538
rect 391492 3398 391520 8162
rect 391676 5438 391704 337554
rect 391768 8226 391796 337742
rect 391756 8220 391808 8226
rect 391756 8162 391808 8168
rect 391860 8106 391888 340054
rect 392044 337618 392072 340068
rect 392518 340054 392900 340082
rect 392978 340054 393268 340082
rect 392872 337770 392900 340054
rect 392872 337742 393176 337770
rect 392032 337612 392084 337618
rect 392032 337554 392084 337560
rect 393044 337612 393096 337618
rect 393044 337554 393096 337560
rect 392584 337272 392636 337278
rect 392584 337214 392636 337220
rect 391768 8078 391888 8106
rect 391664 5432 391716 5438
rect 391664 5374 391716 5380
rect 391768 3602 391796 8078
rect 391756 3596 391808 3602
rect 391756 3538 391808 3544
rect 391848 3528 391900 3534
rect 391848 3470 391900 3476
rect 390652 3392 390704 3398
rect 390652 3334 390704 3340
rect 391480 3392 391532 3398
rect 391480 3334 391532 3340
rect 390664 480 390692 3334
rect 391860 480 391888 3470
rect 392596 2922 392624 337214
rect 393056 5370 393084 337554
rect 393044 5364 393096 5370
rect 393044 5306 393096 5312
rect 393044 3868 393096 3874
rect 393044 3810 393096 3816
rect 392584 2916 392636 2922
rect 392584 2858 392636 2864
rect 393056 480 393084 3810
rect 393148 3738 393176 337742
rect 393136 3732 393188 3738
rect 393136 3674 393188 3680
rect 393240 3602 393268 340054
rect 393424 337142 393452 340068
rect 393884 337822 393912 340068
rect 394266 340054 394648 340082
rect 393964 337952 394016 337958
rect 393964 337894 394016 337900
rect 393872 337816 393924 337822
rect 393872 337758 393924 337764
rect 393412 337136 393464 337142
rect 393412 337078 393464 337084
rect 393228 3596 393280 3602
rect 393228 3538 393280 3544
rect 393976 2854 394004 337894
rect 394424 337816 394476 337822
rect 394424 337758 394476 337764
rect 394436 5234 394464 337758
rect 394516 337136 394568 337142
rect 394516 337078 394568 337084
rect 394528 5302 394556 337078
rect 394516 5296 394568 5302
rect 394516 5238 394568 5244
rect 394424 5228 394476 5234
rect 394424 5170 394476 5176
rect 394620 3534 394648 340054
rect 394712 337482 394740 340068
rect 395186 340054 395568 340082
rect 395646 340054 396028 340082
rect 395344 337884 395396 337890
rect 395344 337826 395396 337832
rect 394700 337476 394752 337482
rect 394700 337418 394752 337424
rect 394608 3528 394660 3534
rect 394608 3470 394660 3476
rect 395356 3466 395384 337826
rect 395540 337736 395568 340054
rect 395540 337708 395936 337736
rect 395804 337476 395856 337482
rect 395804 337418 395856 337424
rect 395816 5166 395844 337418
rect 395804 5160 395856 5166
rect 395804 5102 395856 5108
rect 395908 5098 395936 337708
rect 395896 5092 395948 5098
rect 395896 5034 395948 5040
rect 394240 3460 394292 3466
rect 394240 3402 394292 3408
rect 395344 3460 395396 3466
rect 395344 3402 395396 3408
rect 393964 2848 394016 2854
rect 393964 2790 394016 2796
rect 394252 480 394280 3402
rect 396000 2990 396028 340054
rect 396092 337686 396120 340068
rect 396552 337754 396580 340068
rect 397012 338026 397040 340068
rect 397000 338020 397052 338026
rect 397000 337962 397052 337968
rect 396540 337748 396592 337754
rect 396540 337690 396592 337696
rect 397276 337748 397328 337754
rect 397276 337690 397328 337696
rect 396080 337680 396132 337686
rect 396080 337622 396132 337628
rect 397288 4894 397316 337690
rect 397472 337686 397500 340068
rect 397840 337754 397868 340068
rect 398300 337890 398328 340068
rect 398288 337884 398340 337890
rect 398288 337826 398340 337832
rect 397828 337748 397880 337754
rect 397828 337690 397880 337696
rect 398564 337748 398616 337754
rect 398564 337690 398616 337696
rect 397368 337680 397420 337686
rect 397368 337622 397420 337628
rect 397460 337680 397512 337686
rect 397460 337622 397512 337628
rect 397380 5030 397408 337622
rect 398472 181008 398524 181014
rect 398470 180976 398472 180985
rect 398524 180976 398526 180985
rect 398470 180911 398526 180920
rect 398472 134088 398524 134094
rect 398470 134056 398472 134065
rect 398524 134056 398526 134065
rect 398470 133991 398526 134000
rect 398470 87136 398526 87145
rect 398470 87071 398472 87080
rect 398524 87071 398526 87080
rect 398472 87042 398524 87048
rect 398472 63776 398524 63782
rect 398470 63744 398472 63753
rect 398524 63744 398526 63753
rect 398470 63679 398526 63688
rect 398472 40248 398524 40254
rect 398470 40216 398472 40225
rect 398524 40216 398526 40225
rect 398470 40151 398526 40160
rect 398472 29232 398524 29238
rect 398470 29200 398472 29209
rect 398524 29200 398526 29209
rect 398470 29135 398526 29144
rect 398472 16856 398524 16862
rect 398470 16824 398472 16833
rect 398524 16824 398526 16833
rect 398470 16759 398526 16768
rect 398576 7138 398604 337690
rect 398656 337680 398708 337686
rect 398656 337622 398708 337628
rect 398564 7132 398616 7138
rect 398564 7074 398616 7080
rect 397368 5024 397420 5030
rect 397368 4966 397420 4972
rect 398668 4962 398696 337622
rect 398656 4956 398708 4962
rect 398656 4898 398708 4904
rect 397276 4888 397328 4894
rect 397276 4830 397328 4836
rect 398760 4826 398788 340068
rect 399116 337816 399168 337822
rect 399116 337758 399168 337764
rect 399024 181008 399076 181014
rect 399022 180976 399024 180985
rect 399076 180976 399078 180985
rect 399022 180911 399078 180920
rect 399024 134088 399076 134094
rect 399022 134056 399024 134065
rect 399076 134056 399078 134065
rect 399022 133991 399078 134000
rect 398838 87136 398894 87145
rect 398838 87071 398840 87080
rect 398892 87071 398894 87080
rect 398840 87042 398892 87048
rect 399024 63776 399076 63782
rect 399022 63744 399024 63753
rect 399076 63744 399078 63753
rect 399022 63679 399078 63688
rect 399024 40248 399076 40254
rect 399022 40216 399024 40225
rect 399076 40216 399078 40225
rect 399022 40151 399078 40160
rect 399024 29232 399076 29238
rect 399022 29200 399024 29209
rect 399076 29200 399078 29209
rect 399022 29135 399078 29144
rect 399024 16856 399076 16862
rect 399022 16824 399024 16833
rect 399076 16824 399078 16833
rect 399022 16759 399078 16768
rect 398748 4820 398800 4826
rect 398748 4762 398800 4768
rect 397828 3052 397880 3058
rect 397828 2994 397880 3000
rect 395436 2984 395488 2990
rect 395436 2926 395488 2932
rect 395988 2984 396040 2990
rect 395988 2926 396040 2932
rect 395448 480 395476 2926
rect 396632 2916 396684 2922
rect 396632 2858 396684 2864
rect 396644 480 396672 2858
rect 397840 480 397868 2994
rect 399128 626 399156 337758
rect 399220 337754 399248 340068
rect 399484 337952 399536 337958
rect 399484 337894 399536 337900
rect 399208 337748 399260 337754
rect 399208 337690 399260 337696
rect 399496 2922 399524 337894
rect 399680 337142 399708 340068
rect 400036 337748 400088 337754
rect 400036 337690 400088 337696
rect 399668 337136 399720 337142
rect 399668 337078 399720 337084
rect 400048 8974 400076 337690
rect 400036 8968 400088 8974
rect 400036 8910 400088 8916
rect 400140 4214 400168 340068
rect 400600 337754 400628 340068
rect 400588 337748 400640 337754
rect 400588 337690 400640 337696
rect 401060 337686 401088 340068
rect 401416 337748 401468 337754
rect 401416 337690 401468 337696
rect 401048 337680 401100 337686
rect 401048 337622 401100 337628
rect 401428 8770 401456 337690
rect 401416 8764 401468 8770
rect 401416 8706 401468 8712
rect 401520 5642 401548 340068
rect 401888 337754 401916 340068
rect 401876 337748 401928 337754
rect 401876 337690 401928 337696
rect 402244 337476 402296 337482
rect 402244 337418 402296 337424
rect 401876 337340 401928 337346
rect 401876 337282 401928 337288
rect 401508 5636 401560 5642
rect 401508 5578 401560 5584
rect 400128 4208 400180 4214
rect 400128 4150 400180 4156
rect 400220 3460 400272 3466
rect 400220 3402 400272 3408
rect 399484 2916 399536 2922
rect 399484 2858 399536 2864
rect 399036 598 399156 626
rect 399036 480 399064 598
rect 400232 480 400260 3402
rect 401888 3346 401916 337282
rect 402256 4978 402284 337418
rect 402348 336938 402376 340068
rect 402822 340054 402928 340082
rect 402796 337748 402848 337754
rect 402796 337690 402848 337696
rect 402336 336932 402388 336938
rect 402336 336874 402388 336880
rect 402808 8838 402836 337690
rect 402796 8832 402848 8838
rect 402796 8774 402848 8780
rect 402900 5710 402928 340054
rect 403268 337754 403296 340068
rect 403728 337822 403756 340068
rect 404202 340054 404308 340082
rect 403716 337816 403768 337822
rect 403716 337758 403768 337764
rect 403256 337748 403308 337754
rect 403256 337690 403308 337696
rect 404176 337748 404228 337754
rect 404176 337690 404228 337696
rect 404188 8906 404216 337690
rect 404176 8900 404228 8906
rect 404176 8842 404228 8848
rect 404280 5778 404308 340054
rect 404648 337754 404676 340068
rect 405122 340054 405412 340082
rect 405490 340054 405688 340082
rect 404636 337748 404688 337754
rect 404636 337690 404688 337696
rect 405096 337544 405148 337550
rect 405096 337486 405148 337492
rect 405004 337408 405056 337414
rect 405004 337350 405056 337356
rect 404268 5772 404320 5778
rect 404268 5714 404320 5720
rect 402888 5704 402940 5710
rect 402888 5646 402940 5652
rect 402256 4950 402652 4978
rect 401888 3318 402560 3346
rect 401324 3120 401376 3126
rect 401324 3062 401376 3068
rect 401336 480 401364 3062
rect 402532 480 402560 3318
rect 402624 3058 402652 4950
rect 405016 3398 405044 337350
rect 405004 3392 405056 3398
rect 405004 3334 405056 3340
rect 403716 3188 403768 3194
rect 403716 3130 403768 3136
rect 402612 3052 402664 3058
rect 402612 2994 402664 3000
rect 403728 480 403756 3130
rect 405108 3126 405136 337486
rect 405384 336938 405412 340054
rect 405556 337748 405608 337754
rect 405556 337690 405608 337696
rect 405372 336932 405424 336938
rect 405372 336874 405424 336880
rect 405568 9654 405596 337690
rect 405556 9648 405608 9654
rect 405556 9590 405608 9596
rect 405660 5846 405688 340054
rect 405936 337754 405964 340068
rect 406410 340054 406792 340082
rect 406870 340054 407068 340082
rect 406384 338020 406436 338026
rect 406384 337962 406436 337968
rect 405924 337748 405976 337754
rect 405924 337690 405976 337696
rect 405648 5840 405700 5846
rect 405648 5782 405700 5788
rect 406108 3392 406160 3398
rect 406108 3334 406160 3340
rect 405096 3120 405148 3126
rect 405096 3062 405148 3068
rect 404912 2848 404964 2854
rect 404912 2790 404964 2796
rect 404924 480 404952 2790
rect 406120 480 406148 3334
rect 406396 2854 406424 337962
rect 406764 337958 406792 340054
rect 406752 337952 406804 337958
rect 406752 337894 406804 337900
rect 406936 337748 406988 337754
rect 406936 337690 406988 337696
rect 406948 9586 406976 337690
rect 406936 9580 406988 9586
rect 406936 9522 406988 9528
rect 407040 5914 407068 340054
rect 407316 337754 407344 340068
rect 407790 340054 408080 340082
rect 408250 340054 408448 340082
rect 407304 337748 407356 337754
rect 407304 337690 407356 337696
rect 407764 337612 407816 337618
rect 407764 337554 407816 337560
rect 407028 5908 407080 5914
rect 407028 5850 407080 5856
rect 407776 3330 407804 337554
rect 408052 337278 408080 340054
rect 408316 337748 408368 337754
rect 408316 337690 408368 337696
rect 408040 337272 408092 337278
rect 408040 337214 408092 337220
rect 408328 9518 408356 337690
rect 408316 9512 408368 9518
rect 408316 9454 408368 9460
rect 408420 5982 408448 340054
rect 408696 337618 408724 340068
rect 409064 337754 409092 340068
rect 409538 340054 409828 340082
rect 409144 337884 409196 337890
rect 409144 337826 409196 337832
rect 409052 337748 409104 337754
rect 409052 337690 409104 337696
rect 408684 337612 408736 337618
rect 408684 337554 408736 337560
rect 408408 5976 408460 5982
rect 408408 5918 408460 5924
rect 407304 3324 407356 3330
rect 407304 3266 407356 3272
rect 407764 3324 407816 3330
rect 407764 3266 407816 3272
rect 406384 2848 406436 2854
rect 406384 2790 406436 2796
rect 407316 480 407344 3266
rect 409156 3262 409184 337826
rect 409800 6050 409828 340054
rect 409984 337074 410012 340068
rect 410444 337142 410472 340068
rect 410918 340054 411208 340082
rect 410524 337680 410576 337686
rect 410524 337622 410576 337628
rect 410432 337136 410484 337142
rect 410432 337078 410484 337084
rect 409972 337068 410024 337074
rect 409972 337010 410024 337016
rect 409788 6044 409840 6050
rect 409788 5986 409840 5992
rect 408500 3256 408552 3262
rect 408500 3198 408552 3204
rect 409144 3256 409196 3262
rect 409144 3198 409196 3204
rect 408512 480 408540 3198
rect 409696 3188 409748 3194
rect 409696 3130 409748 3136
rect 409708 480 409736 3130
rect 410536 2990 410564 337622
rect 411180 6118 411208 340054
rect 411364 337414 411392 340068
rect 411824 337550 411852 340068
rect 412298 340054 412588 340082
rect 411904 337816 411956 337822
rect 411904 337758 411956 337764
rect 411812 337544 411864 337550
rect 411812 337486 411864 337492
rect 411352 337408 411404 337414
rect 411352 337350 411404 337356
rect 411168 6112 411220 6118
rect 411168 6054 411220 6060
rect 411916 3194 411944 337758
rect 412560 7206 412588 340054
rect 412652 337686 412680 340068
rect 412640 337680 412692 337686
rect 412640 337622 412692 337628
rect 413112 337210 413140 340068
rect 413586 340054 413876 340082
rect 413100 337204 413152 337210
rect 413100 337146 413152 337152
rect 413848 7274 413876 340054
rect 414032 337754 414060 340068
rect 414020 337748 414072 337754
rect 414020 337690 414072 337696
rect 414492 337686 414520 340068
rect 414966 340054 415256 340082
rect 413928 337680 413980 337686
rect 413928 337622 413980 337628
rect 414480 337680 414532 337686
rect 414480 337622 414532 337628
rect 413836 7268 413888 7274
rect 413836 7210 413888 7216
rect 412548 7200 412600 7206
rect 412548 7142 412600 7148
rect 413940 6866 413968 337622
rect 415228 7342 415256 340054
rect 415308 337748 415360 337754
rect 415308 337690 415360 337696
rect 415216 7336 415268 7342
rect 415216 7278 415268 7284
rect 413928 6860 413980 6866
rect 413928 6802 413980 6808
rect 415320 6798 415348 337690
rect 415412 337482 415440 340068
rect 415872 337958 415900 340068
rect 416346 340054 416544 340082
rect 415860 337952 415912 337958
rect 415860 337894 415912 337900
rect 415400 337476 415452 337482
rect 415400 337418 415452 337424
rect 416516 7410 416544 340054
rect 416596 337476 416648 337482
rect 416596 337418 416648 337424
rect 416504 7404 416556 7410
rect 416504 7346 416556 7352
rect 415308 6792 415360 6798
rect 415308 6734 415360 6740
rect 416608 6730 416636 337418
rect 416596 6724 416648 6730
rect 416596 6666 416648 6672
rect 416700 6662 416728 340068
rect 417160 337686 417188 340068
rect 417634 340054 418016 340082
rect 417424 337884 417476 337890
rect 417424 337826 417476 337832
rect 417148 337680 417200 337686
rect 417148 337622 417200 337628
rect 416688 6656 416740 6662
rect 416688 6598 416740 6604
rect 415676 4684 415728 4690
rect 415676 4626 415728 4632
rect 413284 4616 413336 4622
rect 413284 4558 413336 4564
rect 412548 3256 412600 3262
rect 412548 3198 412600 3204
rect 411904 3188 411956 3194
rect 411904 3130 411956 3136
rect 412088 3120 412140 3126
rect 412088 3062 412140 3068
rect 410524 2984 410576 2990
rect 410524 2926 410576 2932
rect 410892 2916 410944 2922
rect 410892 2858 410944 2864
rect 410904 480 410932 2858
rect 412100 480 412128 3062
rect 412560 2990 412588 3198
rect 412548 2984 412600 2990
rect 412548 2926 412600 2932
rect 413296 480 413324 4558
rect 414480 4072 414532 4078
rect 414480 4014 414532 4020
rect 414492 480 414520 4014
rect 415688 480 415716 4626
rect 416872 4004 416924 4010
rect 416872 3946 416924 3952
rect 416884 480 416912 3946
rect 417436 3194 417464 337826
rect 417884 181008 417936 181014
rect 417882 180976 417884 180985
rect 417936 180976 417938 180985
rect 417882 180911 417938 180920
rect 417884 134088 417936 134094
rect 417882 134056 417884 134065
rect 417936 134056 417938 134065
rect 417882 133991 417938 134000
rect 417884 87168 417936 87174
rect 417882 87136 417884 87145
rect 417936 87136 417938 87145
rect 417882 87071 417938 87080
rect 417882 63744 417938 63753
rect 417882 63679 417884 63688
rect 417936 63679 417938 63688
rect 417884 63650 417936 63656
rect 417884 40248 417936 40254
rect 417882 40216 417884 40225
rect 417936 40216 417938 40225
rect 417882 40151 417938 40160
rect 417882 29200 417938 29209
rect 417882 29135 417884 29144
rect 417936 29135 417938 29144
rect 417884 29106 417936 29112
rect 417882 16824 417938 16833
rect 417882 16759 417938 16768
rect 417896 16425 417924 16759
rect 417882 16416 417938 16425
rect 417882 16351 417938 16360
rect 417988 7478 418016 340054
rect 417976 7472 418028 7478
rect 417976 7414 418028 7420
rect 418080 6594 418108 340068
rect 418540 338094 418568 340068
rect 419014 340054 419396 340082
rect 418528 338088 418580 338094
rect 418528 338030 418580 338036
rect 418344 181008 418396 181014
rect 418342 180976 418344 180985
rect 418396 180976 418398 180985
rect 418342 180911 418398 180920
rect 418344 134088 418396 134094
rect 418342 134056 418344 134065
rect 418396 134056 418398 134065
rect 418342 133991 418398 134000
rect 418344 87168 418396 87174
rect 418342 87136 418344 87145
rect 418396 87136 418398 87145
rect 418342 87071 418398 87080
rect 418344 40248 418396 40254
rect 418342 40216 418344 40225
rect 418396 40216 418398 40225
rect 418342 40151 418398 40160
rect 418158 29200 418214 29209
rect 418158 29135 418160 29144
rect 418212 29135 418214 29144
rect 418160 29106 418212 29112
rect 419368 7546 419396 340054
rect 419356 7540 419408 7546
rect 419356 7482 419408 7488
rect 418068 6588 418120 6594
rect 418068 6530 418120 6536
rect 419460 6526 419488 340068
rect 419920 337278 419948 340068
rect 420184 337816 420236 337822
rect 420184 337758 420236 337764
rect 420656 337770 420684 340190
rect 420762 340054 420868 340082
rect 419908 337272 419960 337278
rect 419908 337214 419960 337220
rect 419630 63744 419686 63753
rect 419630 63679 419632 63688
rect 419684 63679 419686 63688
rect 419632 63650 419684 63656
rect 419448 6520 419500 6526
rect 419448 6462 419500 6468
rect 417976 4140 418028 4146
rect 417976 4082 418028 4088
rect 417424 3188 417476 3194
rect 417424 3130 417476 3136
rect 417988 480 418016 4082
rect 420196 3330 420224 337758
rect 420656 337742 420776 337770
rect 420748 8294 420776 337742
rect 420736 8288 420788 8294
rect 420736 8230 420788 8236
rect 420840 6458 420868 340054
rect 421208 338026 421236 340068
rect 421682 340054 421972 340082
rect 422142 340054 422248 340082
rect 421196 338020 421248 338026
rect 421196 337962 421248 337968
rect 421944 337770 421972 340054
rect 421944 337742 422156 337770
rect 421564 337272 421616 337278
rect 421564 337214 421616 337220
rect 420828 6452 420880 6458
rect 420828 6394 420880 6400
rect 421576 4146 421604 337214
rect 422128 8226 422156 337742
rect 422116 8220 422168 8226
rect 422116 8162 422168 8168
rect 422220 6390 422248 340054
rect 422588 337822 422616 340068
rect 422576 337816 422628 337822
rect 422576 337758 422628 337764
rect 423048 337754 423076 340068
rect 423036 337748 423088 337754
rect 423036 337690 423088 337696
rect 422208 6384 422260 6390
rect 422208 6326 422260 6332
rect 423508 6322 423536 340068
rect 423876 337890 423904 340068
rect 423864 337884 423916 337890
rect 423864 337826 423916 337832
rect 424336 337754 424364 340068
rect 424810 340054 424916 340082
rect 423588 337748 423640 337754
rect 423588 337690 423640 337696
rect 424324 337748 424376 337754
rect 424324 337690 424376 337696
rect 423496 6316 423548 6322
rect 423496 6258 423548 6264
rect 422760 4752 422812 4758
rect 422760 4694 422812 4700
rect 421564 4140 421616 4146
rect 421564 4082 421616 4088
rect 420368 3936 420420 3942
rect 420368 3878 420420 3884
rect 419172 3324 419224 3330
rect 419172 3266 419224 3272
rect 420184 3324 420236 3330
rect 420184 3266 420236 3272
rect 419184 480 419212 3266
rect 420380 480 420408 3878
rect 421564 3868 421616 3874
rect 421564 3810 421616 3816
rect 421576 480 421604 3810
rect 422772 480 422800 4694
rect 423600 4282 423628 337690
rect 424888 6254 424916 340054
rect 424968 337748 425020 337754
rect 424968 337690 425020 337696
rect 424876 6248 424928 6254
rect 424876 6190 424928 6196
rect 423956 5500 424008 5506
rect 423956 5442 424008 5448
rect 423588 4276 423640 4282
rect 423588 4218 423640 4224
rect 423968 480 423996 5442
rect 424980 4350 425008 337690
rect 425256 337686 425284 340068
rect 425716 337754 425744 340068
rect 426190 340054 426296 340082
rect 425704 337748 425756 337754
rect 425704 337690 425756 337696
rect 425244 337680 425296 337686
rect 425244 337622 425296 337628
rect 425150 87272 425206 87281
rect 425150 87207 425206 87216
rect 425058 87000 425114 87009
rect 425164 86986 425192 87207
rect 425114 86958 425192 86986
rect 425058 86935 425114 86944
rect 425060 16720 425112 16726
rect 425058 16688 425060 16697
rect 425112 16688 425114 16697
rect 425058 16623 425114 16632
rect 426268 6186 426296 340054
rect 426636 337822 426664 340068
rect 426624 337816 426676 337822
rect 426624 337758 426676 337764
rect 427096 337754 427124 340068
rect 427570 340054 427676 340082
rect 427176 337952 427228 337958
rect 427176 337894 427228 337900
rect 426348 337748 426400 337754
rect 426348 337690 426400 337696
rect 426992 337748 427044 337754
rect 426992 337690 427044 337696
rect 427084 337748 427136 337754
rect 427084 337690 427136 337696
rect 426256 6180 426308 6186
rect 426256 6122 426308 6128
rect 426360 5658 426388 337690
rect 427004 337634 427032 337690
rect 427188 337634 427216 337894
rect 427004 337606 427216 337634
rect 427648 8158 427676 340054
rect 427924 337754 427952 340068
rect 427728 337748 427780 337754
rect 427728 337690 427780 337696
rect 427912 337748 427964 337754
rect 427912 337690 427964 337696
rect 427636 8152 427688 8158
rect 427636 8094 427688 8100
rect 426268 5630 426388 5658
rect 426268 4418 426296 5630
rect 426348 5432 426400 5438
rect 426348 5374 426400 5380
rect 426256 4412 426308 4418
rect 426256 4354 426308 4360
rect 424968 4344 425020 4350
rect 424968 4286 425020 4292
rect 425152 3052 425204 3058
rect 425152 2994 425204 3000
rect 425164 480 425192 2994
rect 426360 480 426388 5374
rect 427740 4486 427768 337690
rect 428384 337414 428412 340068
rect 428858 340054 429056 340082
rect 428464 337952 428516 337958
rect 428464 337894 428516 337900
rect 428372 337408 428424 337414
rect 428372 337350 428424 337356
rect 427728 4480 427780 4486
rect 427728 4422 427780 4428
rect 428476 4078 428504 337894
rect 429028 8090 429056 340054
rect 429108 337952 429160 337958
rect 429108 337894 429160 337900
rect 429120 337754 429148 337894
rect 429304 337754 429332 340068
rect 429108 337748 429160 337754
rect 429108 337690 429160 337696
rect 429292 337748 429344 337754
rect 429292 337690 429344 337696
rect 429764 337414 429792 340068
rect 430238 340054 430436 340082
rect 430698 340054 431080 340082
rect 429844 337680 429896 337686
rect 429844 337622 429896 337628
rect 429108 337408 429160 337414
rect 429108 337350 429160 337356
rect 429752 337408 429804 337414
rect 429752 337350 429804 337356
rect 429016 8084 429068 8090
rect 429016 8026 429068 8032
rect 429120 4554 429148 337350
rect 429108 4548 429160 4554
rect 429108 4490 429160 4496
rect 428464 4072 428516 4078
rect 428464 4014 428516 4020
rect 429856 4010 429884 337622
rect 430408 8022 430436 340054
rect 431052 338162 431080 340054
rect 431040 338156 431092 338162
rect 431040 338098 431092 338104
rect 431144 337414 431172 340068
rect 431526 340054 431816 340082
rect 431224 338088 431276 338094
rect 431224 338030 431276 338036
rect 430488 337408 430540 337414
rect 430488 337350 430540 337356
rect 431132 337408 431184 337414
rect 431132 337350 431184 337356
rect 430396 8016 430448 8022
rect 430396 7958 430448 7964
rect 429936 5364 429988 5370
rect 429936 5306 429988 5312
rect 429844 4004 429896 4010
rect 429844 3946 429896 3952
rect 427544 3800 427596 3806
rect 427544 3742 427596 3748
rect 427556 480 427584 3742
rect 428740 3732 428792 3738
rect 428740 3674 428792 3680
rect 428752 480 428780 3674
rect 429948 480 429976 5306
rect 430500 4622 430528 337350
rect 430488 4616 430540 4622
rect 430488 4558 430540 4564
rect 431132 3664 431184 3670
rect 431132 3606 431184 3612
rect 431144 480 431172 3606
rect 431236 3398 431264 338030
rect 431788 7954 431816 340054
rect 431972 337754 432000 340068
rect 431960 337748 432012 337754
rect 431960 337690 432012 337696
rect 432432 337414 432460 340068
rect 432906 340054 433196 340082
rect 431868 337408 431920 337414
rect 431868 337350 431920 337356
rect 432420 337408 432472 337414
rect 432420 337350 432472 337356
rect 431776 7948 431828 7954
rect 431776 7890 431828 7896
rect 431880 4690 431908 337350
rect 433168 7886 433196 340054
rect 433352 337482 433380 340068
rect 433340 337476 433392 337482
rect 433340 337418 433392 337424
rect 433812 337414 433840 340068
rect 434286 340054 434484 340082
rect 434746 340054 435036 340082
rect 435114 340054 435496 340082
rect 435574 340054 435956 340082
rect 434076 338156 434128 338162
rect 434076 338098 434128 338104
rect 433984 337544 434036 337550
rect 433984 337486 434036 337492
rect 433248 337408 433300 337414
rect 433248 337350 433300 337356
rect 433800 337408 433852 337414
rect 433800 337350 433852 337356
rect 433156 7880 433208 7886
rect 433156 7822 433208 7828
rect 433260 4758 433288 337350
rect 433524 5296 433576 5302
rect 433524 5238 433576 5244
rect 433248 4752 433300 4758
rect 433248 4694 433300 4700
rect 431868 4684 431920 4690
rect 431868 4626 431920 4632
rect 432328 3596 432380 3602
rect 432328 3538 432380 3544
rect 431224 3392 431276 3398
rect 431224 3334 431276 3340
rect 432340 480 432368 3538
rect 433536 480 433564 5238
rect 433996 3058 434024 337486
rect 434088 3942 434116 338098
rect 434456 318850 434484 340054
rect 435008 337929 435036 340054
rect 434994 337920 435050 337929
rect 434994 337855 435050 337864
rect 435088 337476 435140 337482
rect 435088 337418 435140 337424
rect 434628 337408 434680 337414
rect 434628 337350 434680 337356
rect 434352 318844 434404 318850
rect 434352 318786 434404 318792
rect 434444 318844 434496 318850
rect 434444 318786 434496 318792
rect 434364 311930 434392 318786
rect 434364 311902 434576 311930
rect 434548 309126 434576 311902
rect 434536 309120 434588 309126
rect 434536 309062 434588 309068
rect 434260 299532 434312 299538
rect 434260 299474 434312 299480
rect 434272 299418 434300 299474
rect 434350 299432 434406 299441
rect 434272 299390 434350 299418
rect 434350 299367 434406 299376
rect 434350 289912 434406 289921
rect 434350 289847 434406 289856
rect 434364 289814 434392 289847
rect 434352 289808 434404 289814
rect 434352 289750 434404 289756
rect 434260 280220 434312 280226
rect 434260 280162 434312 280168
rect 434272 280106 434300 280162
rect 434350 280120 434406 280129
rect 434272 280078 434350 280106
rect 434350 280055 434406 280064
rect 434350 270600 434406 270609
rect 434350 270535 434406 270544
rect 434364 270502 434392 270535
rect 434352 270496 434404 270502
rect 434352 270438 434404 270444
rect 434260 260908 434312 260914
rect 434260 260850 434312 260856
rect 434272 260794 434300 260850
rect 434350 260808 434406 260817
rect 434272 260766 434350 260794
rect 434350 260743 434406 260752
rect 434350 251288 434406 251297
rect 434350 251223 434406 251232
rect 434364 251190 434392 251223
rect 434352 251184 434404 251190
rect 434352 251126 434404 251132
rect 434260 241528 434312 241534
rect 434260 241470 434312 241476
rect 434272 234666 434300 241470
rect 434260 234660 434312 234666
rect 434260 234602 434312 234608
rect 434352 234524 434404 234530
rect 434352 234466 434404 234472
rect 434364 225078 434392 234466
rect 434352 225072 434404 225078
rect 434352 225014 434404 225020
rect 434260 224936 434312 224942
rect 434260 224878 434312 224884
rect 434272 220794 434300 224878
rect 434260 220788 434312 220794
rect 434260 220730 434312 220736
rect 434260 215280 434312 215286
rect 434260 215222 434312 215228
rect 434272 211154 434300 215222
rect 434272 211126 434392 211154
rect 434364 202910 434392 211126
rect 434548 202910 434576 202941
rect 434352 202904 434404 202910
rect 434536 202904 434588 202910
rect 434352 202846 434404 202852
rect 434456 202852 434536 202858
rect 434456 202846 434588 202852
rect 434456 202830 434576 202846
rect 434456 196042 434484 202830
rect 434444 196036 434496 196042
rect 434444 195978 434496 195984
rect 434444 193248 434496 193254
rect 434444 193190 434496 193196
rect 434456 183666 434484 193190
rect 434444 183660 434496 183666
rect 434444 183602 434496 183608
rect 434260 183592 434312 183598
rect 434260 183534 434312 183540
rect 434272 173890 434300 183534
rect 434350 173904 434406 173913
rect 434272 173862 434350 173890
rect 434350 173839 434406 173848
rect 434442 164248 434498 164257
rect 434442 164183 434498 164192
rect 434456 159186 434484 164183
rect 434444 159180 434496 159186
rect 434444 159122 434496 159128
rect 434444 154624 434496 154630
rect 434444 154566 434496 154572
rect 434456 147626 434484 154566
rect 434444 147620 434496 147626
rect 434444 147562 434496 147568
rect 434534 143576 434590 143585
rect 434456 143546 434534 143562
rect 434444 143540 434534 143546
rect 434496 143534 434534 143540
rect 434534 143511 434590 143520
rect 434444 143482 434496 143488
rect 434536 137964 434588 137970
rect 434536 137906 434588 137912
rect 434548 128602 434576 137906
rect 434456 128574 434576 128602
rect 434456 120714 434484 128574
rect 434364 120686 434484 120714
rect 434364 109070 434392 120686
rect 434352 109064 434404 109070
rect 434352 109006 434404 109012
rect 434444 108996 434496 109002
rect 434444 108938 434496 108944
rect 434456 104854 434484 108938
rect 434444 104848 434496 104854
rect 434444 104790 434496 104796
rect 434352 95260 434404 95266
rect 434352 95202 434404 95208
rect 434364 91798 434392 95202
rect 434352 91792 434404 91798
rect 434352 91734 434404 91740
rect 434640 87378 434668 337350
rect 435100 321586 435128 337418
rect 435364 336728 435416 336734
rect 435364 336670 435416 336676
rect 435376 335458 435404 336670
rect 435468 335646 435496 340054
rect 435456 335640 435508 335646
rect 435456 335582 435508 335588
rect 435376 335430 435496 335458
rect 435100 321558 435404 321586
rect 435376 316742 435404 321558
rect 435364 316736 435416 316742
rect 435364 316678 435416 316684
rect 435364 302252 435416 302258
rect 435364 302194 435416 302200
rect 435376 297430 435404 302194
rect 435364 297424 435416 297430
rect 435364 297366 435416 297372
rect 435364 282940 435416 282946
rect 435364 282882 435416 282888
rect 435376 278118 435404 282882
rect 435364 278112 435416 278118
rect 435364 278054 435416 278060
rect 435364 263628 435416 263634
rect 435364 263570 435416 263576
rect 435376 263514 435404 263570
rect 435284 263486 435404 263514
rect 435284 260846 435312 263486
rect 435272 260840 435324 260846
rect 435272 260782 435324 260788
rect 435272 251320 435324 251326
rect 435192 251268 435272 251274
rect 435192 251262 435324 251268
rect 435192 251246 435312 251262
rect 435192 251190 435220 251246
rect 435180 251184 435232 251190
rect 435180 251126 435232 251132
rect 435088 241528 435140 241534
rect 435088 241470 435140 241476
rect 435100 234666 435128 241470
rect 435088 234660 435140 234666
rect 435088 234602 435140 234608
rect 435180 234524 435232 234530
rect 435180 234466 435232 234472
rect 435192 231826 435220 234466
rect 435100 231798 435220 231826
rect 435100 225010 435128 231798
rect 435088 225004 435140 225010
rect 435088 224946 435140 224952
rect 435088 222216 435140 222222
rect 435088 222158 435140 222164
rect 435100 215354 435128 222158
rect 435088 215348 435140 215354
rect 435088 215290 435140 215296
rect 435180 215212 435232 215218
rect 435180 215154 435232 215160
rect 435192 212537 435220 215154
rect 435178 212528 435234 212537
rect 435178 212463 435234 212472
rect 435362 212528 435418 212537
rect 435362 212463 435418 212472
rect 435376 202892 435404 212463
rect 435192 202881 435404 202892
rect 435178 202872 435418 202881
rect 435234 202864 435362 202872
rect 435178 202807 435234 202816
rect 435362 202807 435418 202816
rect 435376 195906 435404 202807
rect 435180 195900 435232 195906
rect 435180 195842 435232 195848
rect 435364 195900 435416 195906
rect 435364 195842 435416 195848
rect 435192 186266 435220 195842
rect 435192 186238 435404 186266
rect 435376 167074 435404 186238
rect 435180 167068 435232 167074
rect 435180 167010 435232 167016
rect 435364 167068 435416 167074
rect 435364 167010 435416 167016
rect 435192 165102 435220 167010
rect 435180 165096 435232 165102
rect 435180 165038 435232 165044
rect 435468 147762 435496 335430
rect 435548 316736 435600 316742
rect 435548 316678 435600 316684
rect 435560 302258 435588 316678
rect 435548 302252 435600 302258
rect 435548 302194 435600 302200
rect 435548 297424 435600 297430
rect 435548 297366 435600 297372
rect 435560 282946 435588 297366
rect 435548 282940 435600 282946
rect 435548 282882 435600 282888
rect 435548 278112 435600 278118
rect 435548 278054 435600 278060
rect 435560 263634 435588 278054
rect 435548 263628 435600 263634
rect 435548 263570 435600 263576
rect 435548 165096 435600 165102
rect 435548 165038 435600 165044
rect 435560 147830 435588 165038
rect 435548 147824 435600 147830
rect 435548 147766 435600 147772
rect 435456 147756 435508 147762
rect 435456 147698 435508 147704
rect 434720 147620 434772 147626
rect 434720 147562 434772 147568
rect 435456 147620 435508 147626
rect 435456 147562 435508 147568
rect 435548 147620 435600 147626
rect 435548 147562 435600 147568
rect 434732 143585 434760 147562
rect 434718 143576 434774 143585
rect 434718 143511 434774 143520
rect 435364 138032 435416 138038
rect 435364 137974 435416 137980
rect 435376 125594 435404 137974
rect 435364 125588 435416 125594
rect 435364 125530 435416 125536
rect 435364 109064 435416 109070
rect 435284 109012 435364 109018
rect 435284 109006 435416 109012
rect 435284 108990 435404 109006
rect 435284 99498 435312 108990
rect 435284 99470 435404 99498
rect 435376 99226 435404 99470
rect 435192 99198 435404 99226
rect 434628 87372 434680 87378
rect 434628 87314 434680 87320
rect 434536 87168 434588 87174
rect 434536 87110 434588 87116
rect 434628 87168 434680 87174
rect 435192 87145 435220 99198
rect 434628 87110 434680 87116
rect 435178 87136 435234 87145
rect 434548 80050 434576 87110
rect 434364 80022 434576 80050
rect 434364 75886 434392 80022
rect 434352 75880 434404 75886
rect 434352 75822 434404 75828
rect 434260 66360 434312 66366
rect 434260 66302 434312 66308
rect 434272 66230 434300 66302
rect 434260 66224 434312 66230
rect 434260 66166 434312 66172
rect 434444 66156 434496 66162
rect 434444 66098 434496 66104
rect 434456 60602 434484 66098
rect 434364 60574 434484 60602
rect 434364 51134 434392 60574
rect 434352 51128 434404 51134
rect 434352 51070 434404 51076
rect 434260 51060 434312 51066
rect 434260 51002 434312 51008
rect 434272 48249 434300 51002
rect 434258 48240 434314 48249
rect 434258 48175 434314 48184
rect 434442 41304 434498 41313
rect 434442 41239 434498 41248
rect 434456 35086 434484 41239
rect 434444 35080 434496 35086
rect 434444 35022 434496 35028
rect 434536 29096 434588 29102
rect 434536 29038 434588 29044
rect 434548 27606 434576 29038
rect 434536 27600 434588 27606
rect 434536 27542 434588 27548
rect 434536 18012 434588 18018
rect 434536 17954 434588 17960
rect 434548 17066 434576 17954
rect 434640 17066 434668 87110
rect 435178 87071 435234 87080
rect 435178 87000 435234 87009
rect 435178 86935 435234 86944
rect 435192 85542 435220 86935
rect 435180 85536 435232 85542
rect 435180 85478 435232 85484
rect 435180 75948 435232 75954
rect 435180 75890 435232 75896
rect 435192 67794 435220 75890
rect 435180 67788 435232 67794
rect 435180 67730 435232 67736
rect 435180 67652 435232 67658
rect 435180 67594 435232 67600
rect 435192 66230 435220 67594
rect 435180 66224 435232 66230
rect 435180 66166 435232 66172
rect 435180 51060 435232 51066
rect 435180 51002 435232 51008
rect 435192 48362 435220 51002
rect 435192 48334 435312 48362
rect 435284 48278 435312 48334
rect 435272 48272 435324 48278
rect 435272 48214 435324 48220
rect 435364 38684 435416 38690
rect 435364 38626 435416 38632
rect 435376 28966 435404 38626
rect 435364 28960 435416 28966
rect 435364 28902 435416 28908
rect 435272 19372 435324 19378
rect 435272 19314 435324 19320
rect 434536 17060 434588 17066
rect 434536 17002 434588 17008
rect 434628 17060 434680 17066
rect 434628 17002 434680 17008
rect 434626 16960 434682 16969
rect 434456 16918 434626 16946
rect 434456 16726 434484 16918
rect 434626 16895 434682 16904
rect 434536 16856 434588 16862
rect 434536 16798 434588 16804
rect 434628 16856 434680 16862
rect 434628 16798 434680 16804
rect 434444 16720 434496 16726
rect 434444 16662 434496 16668
rect 434548 7818 434576 16798
rect 434536 7812 434588 7818
rect 434536 7754 434588 7760
rect 434640 5506 434668 16798
rect 435284 12458 435312 19314
rect 435192 12430 435312 12458
rect 434628 5500 434680 5506
rect 434628 5442 434680 5448
rect 434628 5228 434680 5234
rect 434628 5170 434680 5176
rect 434076 3936 434128 3942
rect 434076 3878 434128 3884
rect 433984 3052 434036 3058
rect 433984 2994 434036 3000
rect 434640 480 434668 5170
rect 435192 3806 435220 12430
rect 435180 3800 435232 3806
rect 435180 3742 435232 3748
rect 435468 3602 435496 147562
rect 435560 138038 435588 147562
rect 435548 138032 435600 138038
rect 435548 137974 435600 137980
rect 435548 125588 435600 125594
rect 435548 125530 435600 125536
rect 435560 109070 435588 125530
rect 435548 109064 435600 109070
rect 435548 109006 435600 109012
rect 435928 7750 435956 340054
rect 436020 337414 436048 340068
rect 436480 337686 436508 340068
rect 436954 340054 437336 340082
rect 436376 337680 436428 337686
rect 436376 337622 436428 337628
rect 436468 337680 436520 337686
rect 436468 337622 436520 337628
rect 436008 337408 436060 337414
rect 436008 337350 436060 337356
rect 436008 335640 436060 335646
rect 436008 335582 436060 335588
rect 436388 335594 436416 337622
rect 436836 337408 436888 337414
rect 436836 337350 436888 337356
rect 435916 7744 435968 7750
rect 435916 7686 435968 7692
rect 436020 5438 436048 335582
rect 436388 335566 436784 335594
rect 436008 5432 436060 5438
rect 436008 5374 436060 5380
rect 436756 3874 436784 335566
rect 436744 3868 436796 3874
rect 436744 3810 436796 3816
rect 436848 3738 436876 337350
rect 437308 7682 437336 340054
rect 437400 337890 437428 340068
rect 437388 337884 437440 337890
rect 437388 337826 437440 337832
rect 437388 337680 437440 337686
rect 437388 337622 437440 337628
rect 437296 7676 437348 7682
rect 437296 7618 437348 7624
rect 437400 5370 437428 337622
rect 437860 337414 437888 340068
rect 438334 340054 438716 340082
rect 438214 337920 438270 337929
rect 438214 337855 438270 337864
rect 438228 337618 438256 337855
rect 438216 337612 438268 337618
rect 438216 337554 438268 337560
rect 437848 337408 437900 337414
rect 437848 337350 437900 337356
rect 438124 336660 438176 336666
rect 438124 336602 438176 336608
rect 437388 5364 437440 5370
rect 437388 5306 437440 5312
rect 437020 5160 437072 5166
rect 437020 5102 437072 5108
rect 436836 3732 436888 3738
rect 436836 3674 436888 3680
rect 435456 3596 435508 3602
rect 435456 3538 435508 3544
rect 435824 3528 435876 3534
rect 435824 3470 435876 3476
rect 435836 480 435864 3470
rect 437032 480 437060 5102
rect 438136 3534 438164 336602
rect 438688 7614 438716 340054
rect 438780 337754 438808 340068
rect 438768 337748 438820 337754
rect 438768 337690 438820 337696
rect 439148 337414 439176 340068
rect 439622 340054 440004 340082
rect 440082 340054 440188 340082
rect 438768 337408 438820 337414
rect 438768 337350 438820 337356
rect 439136 337408 439188 337414
rect 439136 337350 439188 337356
rect 438676 7608 438728 7614
rect 438676 7550 438728 7556
rect 438780 5302 438808 337350
rect 439976 9450 440004 340054
rect 440056 337408 440108 337414
rect 440056 337350 440108 337356
rect 439964 9444 440016 9450
rect 439964 9386 440016 9392
rect 438768 5296 438820 5302
rect 438768 5238 438820 5244
rect 440068 5234 440096 337350
rect 440056 5228 440108 5234
rect 440056 5170 440108 5176
rect 438216 5092 438268 5098
rect 438216 5034 438268 5040
rect 438124 3528 438176 3534
rect 438124 3470 438176 3476
rect 438228 480 438256 5034
rect 440160 3670 440188 340054
rect 440528 337414 440556 340068
rect 441002 340054 441292 340082
rect 440516 337408 440568 337414
rect 440516 337350 440568 337356
rect 441264 335594 441292 340054
rect 441448 337686 441476 340068
rect 441436 337680 441488 337686
rect 441436 337622 441488 337628
rect 441908 337414 441936 340068
rect 442382 340054 442580 340082
rect 442750 340054 442948 340082
rect 441528 337408 441580 337414
rect 441528 337350 441580 337356
rect 441896 337408 441948 337414
rect 441896 337350 441948 337356
rect 441264 335566 441476 335594
rect 441448 9382 441476 335566
rect 441436 9376 441488 9382
rect 441436 9318 441488 9324
rect 441540 5166 441568 337350
rect 442264 336524 442316 336530
rect 442264 336466 442316 336472
rect 441528 5160 441580 5166
rect 441528 5102 441580 5108
rect 440608 5024 440660 5030
rect 440608 4966 440660 4972
rect 440148 3664 440200 3670
rect 440148 3606 440200 3612
rect 439412 3460 439464 3466
rect 439412 3402 439464 3408
rect 439424 480 439452 3402
rect 440620 480 440648 4966
rect 441804 4888 441856 4894
rect 441804 4830 441856 4836
rect 441816 480 441844 4830
rect 442276 2922 442304 336466
rect 442552 333282 442580 340054
rect 442816 337408 442868 337414
rect 442816 337350 442868 337356
rect 442552 333254 442764 333282
rect 442736 9314 442764 333254
rect 442724 9308 442776 9314
rect 442724 9250 442776 9256
rect 442828 5098 442856 337350
rect 442816 5092 442868 5098
rect 442816 5034 442868 5040
rect 442920 3602 442948 340054
rect 443196 337414 443224 340068
rect 443670 340054 443960 340082
rect 443184 337408 443236 337414
rect 443184 337350 443236 337356
rect 443932 335594 443960 340054
rect 444116 337754 444144 340068
rect 444104 337748 444156 337754
rect 444104 337690 444156 337696
rect 444576 337414 444604 340068
rect 445050 340054 445340 340082
rect 445510 340054 445708 340082
rect 444840 337680 444892 337686
rect 444840 337622 444892 337628
rect 444852 337550 444880 337622
rect 444840 337544 444892 337550
rect 444840 337486 444892 337492
rect 444288 337408 444340 337414
rect 444288 337350 444340 337356
rect 444564 337408 444616 337414
rect 444564 337350 444616 337356
rect 443932 335566 444236 335594
rect 444208 318850 444236 335566
rect 444104 318844 444156 318850
rect 444104 318786 444156 318792
rect 444196 318844 444248 318850
rect 444196 318786 444248 318792
rect 444116 311982 444144 318786
rect 444104 311976 444156 311982
rect 444104 311918 444156 311924
rect 444196 311976 444248 311982
rect 444196 311918 444248 311924
rect 444208 302258 444236 311918
rect 444012 302252 444064 302258
rect 444012 302194 444064 302200
rect 444196 302252 444248 302258
rect 444196 302194 444248 302200
rect 444024 302138 444052 302194
rect 444024 302110 444144 302138
rect 444116 292618 444144 302110
rect 444116 292590 444236 292618
rect 444208 282946 444236 292590
rect 444012 282940 444064 282946
rect 444012 282882 444064 282888
rect 444196 282940 444248 282946
rect 444196 282882 444248 282888
rect 444024 282826 444052 282882
rect 444024 282798 444144 282826
rect 444116 273306 444144 282798
rect 444116 273278 444236 273306
rect 444208 263634 444236 273278
rect 444012 263628 444064 263634
rect 444012 263570 444064 263576
rect 444196 263628 444248 263634
rect 444196 263570 444248 263576
rect 444024 263514 444052 263570
rect 444024 263486 444144 263514
rect 444116 253994 444144 263486
rect 444116 253966 444236 253994
rect 444208 244322 444236 253966
rect 444012 244316 444064 244322
rect 444012 244258 444064 244264
rect 444196 244316 444248 244322
rect 444196 244258 444248 244264
rect 444024 244202 444052 244258
rect 444024 244174 444144 244202
rect 444116 234682 444144 244174
rect 444116 234654 444236 234682
rect 444208 225010 444236 234654
rect 444012 225004 444064 225010
rect 444012 224946 444064 224952
rect 444196 225004 444248 225010
rect 444196 224946 444248 224952
rect 444024 224890 444052 224946
rect 444024 224862 444144 224890
rect 444116 215370 444144 224862
rect 444116 215342 444236 215370
rect 444208 205698 444236 215342
rect 444012 205692 444064 205698
rect 444012 205634 444064 205640
rect 444196 205692 444248 205698
rect 444196 205634 444248 205640
rect 444024 205578 444052 205634
rect 444024 205550 444144 205578
rect 444116 196058 444144 205550
rect 444116 196030 444236 196058
rect 444208 186386 444236 196030
rect 444012 186380 444064 186386
rect 444012 186322 444064 186328
rect 444196 186380 444248 186386
rect 444196 186322 444248 186328
rect 444024 186266 444052 186322
rect 444024 186238 444144 186266
rect 444116 183569 444144 186238
rect 443918 183560 443974 183569
rect 443918 183495 443974 183504
rect 444102 183560 444158 183569
rect 444102 183495 444158 183504
rect 443932 173942 443960 183495
rect 443920 173936 443972 173942
rect 443920 173878 443972 173884
rect 444104 173936 444156 173942
rect 444104 173878 444156 173884
rect 444116 167090 444144 173878
rect 444024 167062 444144 167090
rect 444024 166954 444052 167062
rect 444024 166926 444144 166954
rect 444116 164218 444144 166926
rect 444104 164212 444156 164218
rect 444104 164154 444156 164160
rect 444104 157344 444156 157350
rect 444104 157286 444156 157292
rect 444116 154578 444144 157286
rect 444116 154562 444236 154578
rect 444116 154556 444248 154562
rect 444116 154550 444196 154556
rect 444196 154498 444248 154504
rect 444208 154467 444236 154498
rect 444104 145036 444156 145042
rect 444104 144978 444156 144984
rect 444116 143546 444144 144978
rect 444104 143540 444156 143546
rect 444104 143482 444156 143488
rect 444104 128308 444156 128314
rect 444104 128250 444156 128256
rect 444116 125594 444144 128250
rect 444104 125588 444156 125594
rect 444104 125530 444156 125536
rect 444196 118652 444248 118658
rect 444196 118594 444248 118600
rect 444208 109070 444236 118594
rect 444012 109064 444064 109070
rect 444196 109064 444248 109070
rect 444064 109012 444144 109018
rect 444012 109006 444144 109012
rect 444196 109006 444248 109012
rect 444024 108990 444144 109006
rect 444116 106282 444144 108990
rect 444104 106276 444156 106282
rect 444104 106218 444156 106224
rect 444104 99340 444156 99346
rect 444104 99282 444156 99288
rect 444116 96642 444144 99282
rect 444116 96614 444236 96642
rect 444208 89758 444236 96614
rect 444012 89752 444064 89758
rect 444196 89752 444248 89758
rect 444064 89700 444144 89706
rect 444012 89694 444144 89700
rect 444196 89694 444248 89700
rect 444024 89678 444144 89694
rect 444116 86970 444144 89678
rect 444104 86964 444156 86970
rect 444104 86906 444156 86912
rect 444196 77308 444248 77314
rect 444196 77250 444248 77256
rect 444208 67658 444236 77250
rect 444104 67652 444156 67658
rect 444104 67594 444156 67600
rect 444196 67652 444248 67658
rect 444196 67594 444248 67600
rect 444116 60858 444144 67594
rect 444104 60852 444156 60858
rect 444104 60794 444156 60800
rect 444012 60716 444064 60722
rect 444012 60658 444064 60664
rect 444024 51066 444052 60658
rect 444012 51060 444064 51066
rect 444012 51002 444064 51008
rect 444196 51060 444248 51066
rect 444196 51002 444248 51008
rect 444208 48278 444236 51002
rect 444196 48272 444248 48278
rect 444196 48214 444248 48220
rect 444104 38684 444156 38690
rect 444104 38626 444156 38632
rect 444116 31890 444144 38626
rect 444104 31884 444156 31890
rect 444104 31826 444156 31832
rect 444104 29028 444156 29034
rect 444104 28970 444156 28976
rect 444116 22114 444144 28970
rect 444116 22086 444236 22114
rect 444208 12458 444236 22086
rect 444024 12430 444236 12458
rect 444024 9246 444052 12430
rect 444012 9240 444064 9246
rect 444012 9182 444064 9188
rect 444300 5030 444328 337350
rect 445312 331922 445340 340054
rect 445576 337408 445628 337414
rect 445576 337350 445628 337356
rect 445312 331894 445524 331922
rect 444380 87032 444432 87038
rect 444378 87000 444380 87009
rect 444432 87000 444434 87009
rect 444378 86935 444434 86944
rect 444380 29096 444432 29102
rect 444378 29064 444380 29073
rect 444432 29064 444434 29073
rect 444378 28999 444434 29008
rect 444380 16720 444432 16726
rect 444378 16688 444380 16697
rect 444432 16688 444434 16697
rect 444378 16623 444434 16632
rect 445496 9178 445524 331894
rect 445484 9172 445536 9178
rect 445484 9114 445536 9120
rect 445392 7132 445444 7138
rect 445392 7074 445444 7080
rect 444288 5024 444340 5030
rect 444288 4966 444340 4972
rect 444196 4956 444248 4962
rect 444196 4898 444248 4904
rect 442908 3596 442960 3602
rect 442908 3538 442960 3544
rect 442264 2916 442316 2922
rect 442264 2858 442316 2864
rect 443000 2848 443052 2854
rect 443000 2790 443052 2796
rect 443012 480 443040 2790
rect 444208 480 444236 4898
rect 445404 480 445432 7074
rect 445588 4962 445616 337350
rect 445576 4956 445628 4962
rect 445576 4898 445628 4904
rect 445680 2854 445708 340054
rect 445956 337686 445984 340068
rect 446338 340054 446628 340082
rect 446798 340054 447088 340082
rect 445944 337680 445996 337686
rect 445944 337622 445996 337628
rect 446600 335594 446628 340054
rect 447060 337906 447088 340054
rect 447060 337878 447180 337906
rect 447048 337680 447100 337686
rect 447048 337622 447100 337628
rect 446600 335566 446996 335594
rect 446968 9110 446996 335566
rect 446956 9104 447008 9110
rect 446956 9046 447008 9052
rect 447060 4894 447088 337622
rect 447152 337498 447180 337878
rect 447244 337686 447272 340068
rect 447232 337680 447284 337686
rect 448072 337668 448100 340190
rect 448164 337793 448192 340068
rect 448150 337784 448206 337793
rect 448150 337719 448206 337728
rect 448624 337686 448652 340068
rect 449098 340054 449388 340082
rect 449162 337784 449218 337793
rect 449162 337719 449218 337728
rect 448428 337680 448480 337686
rect 448072 337640 448376 337668
rect 447232 337622 447284 337628
rect 447324 337612 447376 337618
rect 447324 337554 447376 337560
rect 447336 337498 447364 337554
rect 447152 337470 447364 337498
rect 447230 134328 447286 134337
rect 447230 134263 447286 134272
rect 447138 134056 447194 134065
rect 447244 134042 447272 134263
rect 447194 134014 447272 134042
rect 447138 133991 447194 134000
rect 447230 64016 447286 64025
rect 447230 63951 447286 63960
rect 447138 63744 447194 63753
rect 447244 63730 447272 63951
rect 447194 63702 447272 63730
rect 447138 63679 447194 63688
rect 447230 40488 447286 40497
rect 447230 40423 447286 40432
rect 447138 40216 447194 40225
rect 447244 40202 447272 40423
rect 447194 40174 447272 40202
rect 447138 40151 447194 40160
rect 447230 16960 447286 16969
rect 447230 16895 447286 16904
rect 447244 16726 447272 16895
rect 447232 16720 447284 16726
rect 447232 16662 447284 16668
rect 448348 9042 448376 337640
rect 448428 337622 448480 337628
rect 448612 337680 448664 337686
rect 448612 337622 448664 337628
rect 448336 9036 448388 9042
rect 448336 8978 448388 8984
rect 447048 4888 447100 4894
rect 447048 4830 447100 4836
rect 448440 4826 448468 337622
rect 448980 8968 449032 8974
rect 448980 8910 449032 8916
rect 447784 4820 447836 4826
rect 447784 4762 447836 4768
rect 448428 4820 448480 4826
rect 448428 4762 448480 4768
rect 446588 2984 446640 2990
rect 446588 2926 446640 2932
rect 445668 2848 445720 2854
rect 445668 2790 445720 2796
rect 446600 480 446628 2926
rect 447796 480 447824 4762
rect 448992 480 449020 8910
rect 449176 3534 449204 337719
rect 449360 337226 449388 340054
rect 449544 337385 449572 340068
rect 502984 338088 503036 338094
rect 502984 338030 503036 338036
rect 500224 338020 500276 338026
rect 500224 337962 500276 337968
rect 449808 337680 449860 337686
rect 449808 337622 449860 337628
rect 449530 337376 449586 337385
rect 449530 337311 449586 337320
rect 449360 337198 449756 337226
rect 449254 87272 449310 87281
rect 449254 87207 449310 87216
rect 449268 87038 449296 87207
rect 449256 87032 449308 87038
rect 449256 86974 449308 86980
rect 449254 29336 449310 29345
rect 449254 29271 449310 29280
rect 449268 29102 449296 29271
rect 449256 29096 449308 29102
rect 449256 29038 449308 29044
rect 449728 8974 449756 337198
rect 449716 8968 449768 8974
rect 449716 8910 449768 8916
rect 449820 4865 449848 337622
rect 496084 337340 496136 337346
rect 496084 337282 496136 337288
rect 492680 337272 492732 337278
rect 492680 337214 492732 337220
rect 485780 337204 485832 337210
rect 485780 337146 485832 337152
rect 477500 337136 477552 337142
rect 477500 337078 477552 337084
rect 470600 337000 470652 337006
rect 470600 336942 470652 336948
rect 463700 336932 463752 336938
rect 463700 336874 463752 336880
rect 456800 336864 456852 336870
rect 456800 336806 456852 336812
rect 449900 336728 449952 336734
rect 449900 336670 449952 336676
rect 449806 4856 449862 4865
rect 449806 4791 449862 4800
rect 449164 3528 449216 3534
rect 449164 3470 449216 3476
rect 449912 626 449940 336670
rect 454406 180976 454462 180985
rect 454406 180911 454408 180920
rect 454460 180911 454462 180920
rect 454408 180882 454460 180888
rect 456064 8832 456116 8838
rect 456064 8774 456116 8780
rect 452476 8764 452528 8770
rect 452476 8706 452528 8712
rect 451280 4208 451332 4214
rect 451280 4150 451332 4156
rect 449912 598 450216 626
rect 450188 480 450216 598
rect 451292 480 451320 4150
rect 452488 480 452516 8706
rect 454868 5636 454920 5642
rect 454868 5578 454920 5584
rect 453672 3460 453724 3466
rect 453672 3402 453724 3408
rect 453684 480 453712 3402
rect 454880 480 454908 5578
rect 456076 480 456104 8774
rect 456812 3346 456840 336806
rect 458362 180976 458418 180985
rect 458362 180911 458364 180920
rect 458416 180911 458418 180920
rect 458364 180882 458416 180888
rect 460846 134600 460902 134609
rect 460846 134535 460902 134544
rect 460860 134201 460888 134535
rect 460846 134192 460902 134201
rect 460846 134127 460902 134136
rect 463606 87544 463662 87553
rect 463606 87479 463662 87488
rect 463620 87145 463648 87479
rect 463606 87136 463662 87145
rect 463606 87071 463662 87080
rect 460846 64288 460902 64297
rect 460846 64223 460902 64232
rect 460860 63889 460888 64223
rect 460846 63880 460902 63889
rect 460846 63815 460902 63824
rect 460846 40760 460902 40769
rect 460846 40695 460902 40704
rect 460860 40361 460888 40695
rect 460846 40352 460902 40361
rect 460846 40287 460902 40296
rect 463240 9648 463292 9654
rect 463240 9590 463292 9596
rect 459652 8900 459704 8906
rect 459652 8842 459704 8848
rect 458456 5704 458508 5710
rect 458456 5646 458508 5652
rect 456812 3318 457300 3346
rect 457272 480 457300 3318
rect 458468 480 458496 5646
rect 459664 480 459692 8842
rect 462044 5772 462096 5778
rect 462044 5714 462096 5720
rect 460848 3120 460900 3126
rect 460848 3062 460900 3068
rect 460860 480 460888 3062
rect 462056 480 462084 5714
rect 463252 480 463280 9590
rect 463712 3482 463740 336874
rect 463792 87032 463844 87038
rect 463790 87000 463792 87009
rect 466552 87032 466604 87038
rect 463844 87000 463846 87009
rect 463790 86935 463846 86944
rect 466550 87000 466552 87009
rect 466604 87000 466606 87009
rect 466550 86935 466606 86944
rect 466828 9580 466880 9586
rect 466828 9522 466880 9528
rect 465632 5840 465684 5846
rect 465632 5782 465684 5788
rect 463712 3454 464476 3482
rect 464448 480 464476 3454
rect 465644 480 465672 5782
rect 466840 480 466868 9522
rect 470324 9512 470376 9518
rect 470324 9454 470376 9460
rect 469128 5908 469180 5914
rect 469128 5850 469180 5856
rect 467932 3188 467984 3194
rect 467932 3130 467984 3136
rect 467944 480 467972 3130
rect 469140 480 469168 5850
rect 470336 480 470364 9454
rect 470612 3346 470640 336942
rect 471886 29472 471942 29481
rect 471886 29407 471942 29416
rect 471900 29073 471928 29407
rect 476028 29232 476080 29238
rect 476026 29200 476028 29209
rect 476080 29200 476082 29209
rect 476026 29135 476082 29144
rect 471886 29064 471942 29073
rect 471886 28999 471942 29008
rect 471886 17096 471942 17105
rect 471886 17031 471942 17040
rect 471900 16697 471928 17031
rect 476028 16856 476080 16862
rect 476026 16824 476028 16833
rect 476080 16824 476082 16833
rect 476026 16759 476082 16768
rect 471886 16688 471942 16697
rect 471886 16623 471942 16632
rect 476304 6044 476356 6050
rect 476304 5986 476356 5992
rect 472716 5976 472768 5982
rect 472716 5918 472768 5924
rect 470612 3318 471560 3346
rect 471532 480 471560 3318
rect 472728 480 472756 5918
rect 475108 3324 475160 3330
rect 475108 3266 475160 3272
rect 473912 2848 473964 2854
rect 473912 2790 473964 2796
rect 473924 480 473952 2790
rect 475120 480 475148 3266
rect 476316 480 476344 5986
rect 477512 4214 477540 337078
rect 477592 337068 477644 337074
rect 477592 337010 477644 337016
rect 477500 4208 477552 4214
rect 477500 4150 477552 4156
rect 477604 3482 477632 337010
rect 482926 29336 482982 29345
rect 482926 29271 482982 29280
rect 482940 29238 482968 29271
rect 482928 29232 482980 29238
rect 482928 29174 482980 29180
rect 482926 16960 482982 16969
rect 482926 16895 482982 16904
rect 482940 16862 482968 16895
rect 482928 16856 482980 16862
rect 482928 16798 482980 16804
rect 483480 7200 483532 7206
rect 483480 7142 483532 7148
rect 479892 6112 479944 6118
rect 479892 6054 479944 6060
rect 478696 4208 478748 4214
rect 478696 4150 478748 4156
rect 477512 3454 477632 3482
rect 477512 480 477540 3454
rect 478708 480 478736 4150
rect 479904 480 479932 6054
rect 481088 3052 481140 3058
rect 481088 2994 481140 3000
rect 481100 480 481128 2994
rect 482284 2984 482336 2990
rect 482284 2926 482336 2932
rect 482296 480 482324 2926
rect 483492 480 483520 7142
rect 484584 6860 484636 6866
rect 484584 6802 484636 6808
rect 484596 480 484624 6802
rect 485792 480 485820 337146
rect 490564 7336 490616 7342
rect 490564 7278 490616 7284
rect 486976 7268 487028 7274
rect 486976 7210 487028 7216
rect 486988 480 487016 7210
rect 488172 6792 488224 6798
rect 488172 6734 488224 6740
rect 488184 480 488212 6734
rect 489368 3256 489420 3262
rect 489368 3198 489420 3204
rect 489380 480 489408 3198
rect 490576 480 490604 7278
rect 491760 6724 491812 6730
rect 491760 6666 491812 6672
rect 491772 480 491800 6666
rect 492692 610 492720 337214
rect 494152 7404 494204 7410
rect 494152 7346 494204 7352
rect 492680 604 492732 610
rect 492680 546 492732 552
rect 492956 604 493008 610
rect 492956 546 493008 552
rect 492968 480 492996 546
rect 494164 480 494192 7346
rect 495348 6656 495400 6662
rect 495348 6598 495400 6604
rect 495360 480 495388 6598
rect 496096 3194 496124 337282
rect 497740 7472 497792 7478
rect 497740 7414 497792 7420
rect 496544 3392 496596 3398
rect 496544 3334 496596 3340
rect 496084 3188 496136 3194
rect 496084 3130 496136 3136
rect 496556 480 496584 3334
rect 497752 480 497780 7414
rect 498936 6588 498988 6594
rect 498936 6530 498988 6536
rect 498948 480 498976 6530
rect 500236 3398 500264 337962
rect 501236 7540 501288 7546
rect 501236 7482 501288 7488
rect 500224 3392 500276 3398
rect 500224 3334 500276 3340
rect 500132 3188 500184 3194
rect 500132 3130 500184 3136
rect 500144 480 500172 3130
rect 501248 480 501276 7482
rect 502432 6520 502484 6526
rect 502432 6462 502484 6468
rect 502444 480 502472 6462
rect 502996 3262 503024 338030
rect 507124 337952 507176 337958
rect 507124 337894 507176 337900
rect 504824 8288 504876 8294
rect 504824 8230 504876 8236
rect 503628 4140 503680 4146
rect 503628 4082 503680 4088
rect 502984 3256 503036 3262
rect 502984 3198 503036 3204
rect 503640 480 503668 4082
rect 504836 480 504864 8230
rect 506020 6452 506072 6458
rect 506020 6394 506072 6400
rect 506032 480 506060 6394
rect 507136 4146 507164 337894
rect 514024 337884 514076 337890
rect 514024 337826 514076 337832
rect 511264 337816 511316 337822
rect 511264 337758 511316 337764
rect 508412 8220 508464 8226
rect 508412 8162 508464 8168
rect 507124 4140 507176 4146
rect 507124 4082 507176 4088
rect 507216 3392 507268 3398
rect 507216 3334 507268 3340
rect 507228 480 507256 3334
rect 508424 480 508452 8162
rect 509608 6384 509660 6390
rect 509608 6326 509660 6332
rect 509620 480 509648 6326
rect 510804 4072 510856 4078
rect 510804 4014 510856 4020
rect 510816 480 510844 4014
rect 511276 3126 511304 337758
rect 513196 6316 513248 6322
rect 513196 6258 513248 6264
rect 512000 4276 512052 4282
rect 512000 4218 512052 4224
rect 511264 3120 511316 3126
rect 511264 3062 511316 3068
rect 512012 480 512040 4218
rect 513208 480 513236 6258
rect 514036 3194 514064 337826
rect 518164 337748 518216 337754
rect 518164 337690 518216 337696
rect 516784 6248 516836 6254
rect 516784 6190 516836 6196
rect 515588 4344 515640 4350
rect 515588 4286 515640 4292
rect 514392 3392 514444 3398
rect 514392 3334 514444 3340
rect 514024 3188 514076 3194
rect 514024 3130 514076 3136
rect 514404 480 514432 3334
rect 515600 480 515628 4286
rect 516796 480 516824 6190
rect 517888 4004 517940 4010
rect 517888 3946 517940 3952
rect 517900 480 517928 3946
rect 518176 3262 518204 337690
rect 529204 337680 529256 337686
rect 529204 337622 529256 337628
rect 527824 337612 527876 337618
rect 527824 337554 527876 337560
rect 525064 337544 525116 337550
rect 525064 337486 525116 337492
rect 520924 337476 520976 337482
rect 520924 337418 520976 337424
rect 520280 6180 520332 6186
rect 520280 6122 520332 6128
rect 519084 4412 519136 4418
rect 519084 4354 519136 4360
rect 518164 3256 518216 3262
rect 518164 3198 518216 3204
rect 519096 480 519124 4354
rect 520292 480 520320 6122
rect 520936 3330 520964 337418
rect 523684 337408 523736 337414
rect 523684 337350 523736 337356
rect 522672 4480 522724 4486
rect 522672 4422 522724 4428
rect 521476 4140 521528 4146
rect 521476 4082 521528 4088
rect 520924 3324 520976 3330
rect 520924 3266 520976 3272
rect 521488 480 521516 4082
rect 522684 480 522712 4422
rect 523696 3398 523724 337350
rect 523868 8152 523920 8158
rect 523868 8094 523920 8100
rect 523684 3392 523736 3398
rect 523684 3334 523736 3340
rect 523880 480 523908 8094
rect 525076 4146 525104 337486
rect 527456 8084 527508 8090
rect 527456 8026 527508 8032
rect 526260 4548 526312 4554
rect 526260 4490 526312 4496
rect 525064 4140 525116 4146
rect 525064 4082 525116 4088
rect 525064 3936 525116 3942
rect 525064 3878 525116 3884
rect 525076 480 525104 3878
rect 526272 480 526300 4490
rect 527468 480 527496 8026
rect 527836 4078 527864 337554
rect 527824 4072 527876 4078
rect 527824 4014 527876 4020
rect 529216 4010 529244 337622
rect 530582 337376 530638 337385
rect 530582 337311 530638 337320
rect 529848 4616 529900 4622
rect 529848 4558 529900 4564
rect 529204 4004 529256 4010
rect 529204 3946 529256 3952
rect 528652 3120 528704 3126
rect 528652 3062 528704 3068
rect 528664 480 528692 3062
rect 529860 480 529888 4558
rect 530596 3942 530624 337311
rect 577516 299470 577544 559846
rect 577608 322930 577636 559914
rect 579712 557524 579764 557530
rect 579712 557466 579764 557472
rect 579724 557297 579752 557466
rect 579710 557288 579766 557297
rect 579710 557223 579766 557232
rect 579816 552702 579844 560186
rect 580080 560176 580132 560182
rect 580080 560118 580132 560124
rect 579896 560108 579948 560114
rect 579896 560050 579948 560056
rect 579804 552696 579856 552702
rect 579804 552638 579856 552644
rect 579804 546440 579856 546446
rect 579804 546382 579856 546388
rect 579816 545601 579844 546382
rect 579802 545592 579858 545601
rect 579802 545527 579858 545536
rect 579804 534064 579856 534070
rect 579804 534006 579856 534012
rect 579816 533905 579844 534006
rect 579802 533896 579858 533905
rect 579802 533831 579858 533840
rect 579804 510604 579856 510610
rect 579804 510546 579856 510552
rect 579816 510377 579844 510546
rect 579802 510368 579858 510377
rect 579802 510303 579858 510312
rect 579804 499520 579856 499526
rect 579804 499462 579856 499468
rect 579816 498681 579844 499462
rect 579802 498672 579858 498681
rect 579802 498607 579858 498616
rect 579804 463684 579856 463690
rect 579804 463626 579856 463632
rect 579816 463457 579844 463626
rect 579802 463448 579858 463457
rect 579802 463383 579858 463392
rect 579804 452600 579856 452606
rect 579804 452542 579856 452548
rect 579816 451761 579844 452542
rect 579802 451752 579858 451761
rect 579802 451687 579858 451696
rect 579804 440224 579856 440230
rect 579804 440166 579856 440172
rect 579816 439929 579844 440166
rect 579802 439920 579858 439929
rect 579802 439855 579858 439864
rect 579804 416764 579856 416770
rect 579804 416706 579856 416712
rect 579816 416537 579844 416706
rect 579802 416528 579858 416537
rect 579802 416463 579858 416472
rect 579804 405680 579856 405686
rect 579804 405622 579856 405628
rect 579816 404841 579844 405622
rect 579802 404832 579858 404841
rect 579802 404767 579858 404776
rect 579804 393304 579856 393310
rect 579804 393246 579856 393252
rect 579816 393009 579844 393246
rect 579802 393000 579858 393009
rect 579802 392935 579858 392944
rect 579804 369844 579856 369850
rect 579804 369786 579856 369792
rect 579816 369617 579844 369786
rect 579802 369608 579858 369617
rect 579802 369543 579858 369552
rect 579908 357921 579936 560050
rect 579988 560040 580040 560046
rect 579988 559982 580040 559988
rect 579894 357912 579950 357921
rect 579894 357847 579950 357856
rect 579896 346384 579948 346390
rect 579896 346326 579948 346332
rect 579908 346089 579936 346326
rect 579894 346080 579950 346089
rect 579894 346015 579950 346024
rect 577596 322924 577648 322930
rect 577596 322866 577648 322872
rect 579896 322924 579948 322930
rect 579896 322866 579948 322872
rect 579908 322697 579936 322866
rect 579894 322688 579950 322697
rect 579894 322623 579950 322632
rect 580000 310865 580028 559982
rect 579986 310856 580042 310865
rect 579986 310791 580042 310800
rect 577504 299464 577556 299470
rect 577504 299406 577556 299412
rect 579896 299464 579948 299470
rect 579896 299406 579948 299412
rect 579908 299169 579936 299406
rect 579894 299160 579950 299169
rect 579894 299095 579950 299104
rect 580092 275777 580120 560118
rect 580172 559836 580224 559842
rect 580172 559778 580224 559784
rect 580078 275768 580134 275777
rect 580078 275703 580134 275712
rect 580184 263945 580212 559778
rect 580264 559496 580316 559502
rect 580264 559438 580316 559444
rect 580170 263936 580226 263945
rect 580170 263871 580226 263880
rect 580276 76265 580304 559438
rect 580368 111489 580396 562391
rect 580448 559564 580500 559570
rect 580448 559506 580500 559512
rect 580460 123185 580488 559506
rect 580552 158409 580580 562527
rect 580908 562488 580960 562494
rect 580908 562430 580960 562436
rect 580724 559700 580776 559706
rect 580724 559642 580776 559648
rect 580632 559632 580684 559638
rect 580632 559574 580684 559580
rect 580644 170105 580672 559574
rect 580736 217025 580764 559642
rect 580816 552696 580868 552702
rect 580816 552638 580868 552644
rect 580828 228857 580856 552638
rect 580920 252249 580948 562430
rect 580906 252240 580962 252249
rect 580906 252175 580962 252184
rect 580814 228848 580870 228857
rect 580814 228783 580870 228792
rect 580722 217016 580778 217025
rect 580722 216951 580778 216960
rect 580630 170096 580686 170105
rect 580630 170031 580686 170040
rect 580538 158400 580594 158409
rect 580538 158335 580594 158344
rect 580446 123176 580502 123185
rect 580446 123111 580502 123120
rect 580354 111480 580410 111489
rect 580354 111415 580410 111424
rect 580262 76256 580318 76265
rect 580262 76191 580318 76200
rect 555976 9444 556028 9450
rect 555976 9386 556028 9392
rect 531044 8016 531096 8022
rect 531044 7958 531096 7964
rect 530584 3936 530636 3942
rect 530584 3878 530636 3884
rect 531056 480 531084 7958
rect 534540 7948 534592 7954
rect 534540 7890 534592 7896
rect 533436 4684 533488 4690
rect 533436 4626 533488 4632
rect 532240 3868 532292 3874
rect 532240 3810 532292 3816
rect 532252 480 532280 3810
rect 533448 480 533476 4626
rect 534552 480 534580 7890
rect 538128 7880 538180 7886
rect 538128 7822 538180 7828
rect 536932 4752 536984 4758
rect 536932 4694 536984 4700
rect 535736 3188 535788 3194
rect 535736 3130 535788 3136
rect 535748 480 535776 3130
rect 536944 480 536972 4694
rect 538140 480 538168 7822
rect 541716 7812 541768 7818
rect 541716 7754 541768 7760
rect 540520 5500 540572 5506
rect 540520 5442 540572 5448
rect 539324 3800 539376 3806
rect 539324 3742 539376 3748
rect 539336 480 539364 3742
rect 540532 480 540560 5442
rect 541728 480 541756 7754
rect 545304 7744 545356 7750
rect 545304 7686 545356 7692
rect 544108 5432 544160 5438
rect 544108 5374 544160 5380
rect 542912 3256 542964 3262
rect 542912 3198 542964 3204
rect 542924 480 542952 3198
rect 544120 480 544148 5374
rect 545316 480 545344 7686
rect 548892 7676 548944 7682
rect 548892 7618 548944 7624
rect 547696 5364 547748 5370
rect 547696 5306 547748 5312
rect 546500 3732 546552 3738
rect 546500 3674 546552 3680
rect 546512 480 546540 3674
rect 547708 480 547736 5306
rect 548904 480 548932 7618
rect 552388 7608 552440 7614
rect 552388 7550 552440 7556
rect 551192 5296 551244 5302
rect 551192 5238 551244 5244
rect 550088 3324 550140 3330
rect 550088 3266 550140 3272
rect 550100 480 550128 3266
rect 551204 480 551232 5238
rect 552400 480 552428 7550
rect 554780 5228 554832 5234
rect 554780 5170 554832 5176
rect 553584 3392 553636 3398
rect 553584 3334 553636 3340
rect 553596 480 553624 3334
rect 554792 480 554820 5170
rect 555988 480 556016 9386
rect 559564 9376 559616 9382
rect 559564 9318 559616 9324
rect 558368 5160 558420 5166
rect 558368 5102 558420 5108
rect 557172 3664 557224 3670
rect 557172 3606 557224 3612
rect 557184 480 557212 3606
rect 558380 480 558408 5102
rect 559576 480 559604 9318
rect 563152 9308 563204 9314
rect 563152 9250 563204 9256
rect 561956 5092 562008 5098
rect 561956 5034 562008 5040
rect 560760 4140 560812 4146
rect 560760 4082 560812 4088
rect 560772 480 560800 4082
rect 561968 480 561996 5034
rect 563164 480 563192 9250
rect 566740 9240 566792 9246
rect 566740 9182 566792 9188
rect 565544 5024 565596 5030
rect 565544 4966 565596 4972
rect 564348 3596 564400 3602
rect 564348 3538 564400 3544
rect 564360 480 564388 3538
rect 565556 480 565584 4966
rect 566752 480 566780 9182
rect 570236 9172 570288 9178
rect 570236 9114 570288 9120
rect 569040 4956 569092 4962
rect 569040 4898 569092 4904
rect 567844 4072 567896 4078
rect 567844 4014 567896 4020
rect 567856 480 567884 4014
rect 569052 480 569080 4898
rect 570248 480 570276 9114
rect 573824 9104 573876 9110
rect 573824 9046 573876 9052
rect 572628 4888 572680 4894
rect 572628 4830 572680 4836
rect 571432 3528 571484 3534
rect 571432 3470 571484 3476
rect 571444 480 571472 3470
rect 572640 480 572668 4830
rect 573836 480 573864 9046
rect 577412 9036 577464 9042
rect 577412 8978 577464 8984
rect 576216 4820 576268 4826
rect 576216 4762 576268 4768
rect 575020 4004 575072 4010
rect 575020 3946 575072 3952
rect 575032 480 575060 3946
rect 576228 480 576256 4762
rect 577424 480 577452 8978
rect 581000 8968 581052 8974
rect 581000 8910 581052 8916
rect 579802 4856 579858 4865
rect 579802 4791 579858 4800
rect 578608 3460 578660 3466
rect 578608 3402 578660 3408
rect 578620 480 578648 3402
rect 579816 480 579844 4791
rect 581012 480 581040 8910
rect 582196 3936 582248 3942
rect 582196 3878 582248 3884
rect 582208 480 582236 3878
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 8114 700304 8170 700360
rect 3514 682216 3570 682272
rect 3422 667956 3478 667992
rect 3422 667936 3424 667956
rect 3424 667936 3476 667956
rect 3476 667936 3478 667956
rect 3054 653520 3110 653576
rect 3422 624824 3478 624880
rect 3422 610408 3478 610464
rect 3238 595992 3294 596048
rect 3422 567296 3478 567352
rect 249982 562944 250038 563000
rect 288622 562944 288678 563000
rect 4158 562672 4214 562728
rect 3974 562536 4030 562592
rect 2962 558184 3018 558240
rect 2778 553052 2780 553072
rect 2780 553052 2832 553072
rect 2832 553052 2834 553072
rect 2778 553016 2834 553052
rect 2962 538600 3018 538656
rect 3790 562264 3846 562320
rect 3054 509904 3110 509960
rect 3054 495524 3056 495544
rect 3056 495524 3108 495544
rect 3108 495524 3110 495544
rect 3054 495488 3110 495524
rect 3054 481108 3056 481128
rect 3056 481108 3108 481128
rect 3108 481108 3110 481128
rect 3054 481072 3110 481108
rect 3146 452376 3202 452432
rect 3146 437960 3202 438016
rect 2778 423680 2834 423736
rect 3238 394984 3294 395040
rect 3146 380604 3148 380624
rect 3148 380604 3200 380624
rect 3200 380604 3202 380624
rect 3146 380568 3202 380604
rect 2778 366152 2834 366208
rect 3606 561720 3662 561776
rect 3422 559000 3478 559056
rect 3330 323040 3386 323096
rect 2778 294344 2834 294400
rect 3146 280100 3148 280120
rect 3148 280100 3200 280120
rect 3200 280100 3202 280120
rect 3146 280064 3202 280100
rect 3146 252456 3202 252512
rect 3146 251232 3202 251288
rect 2778 208156 2780 208176
rect 2780 208156 2832 208176
rect 2832 208156 2834 208176
rect 2778 208120 2834 208156
rect 2778 179424 2834 179480
rect 2778 165008 2834 165064
rect 2778 136348 2780 136368
rect 2780 136348 2832 136368
rect 2832 136348 2834 136368
rect 2778 136312 2834 136348
rect 2778 122068 2780 122088
rect 2780 122068 2832 122088
rect 2832 122068 2834 122088
rect 2778 122032 2834 122068
rect 2778 78920 2834 78976
rect 4066 265648 4122 265704
rect 3974 236952 4030 237008
rect 3882 222536 3938 222592
rect 3790 193840 3846 193896
rect 3698 150728 3754 150784
rect 3606 107616 3662 107672
rect 3514 93200 3570 93256
rect 3422 64504 3478 64560
rect 4066 50088 4122 50144
rect 242254 562536 242310 562592
rect 248050 562536 248106 562592
rect 5354 562264 5410 562320
rect 5078 562128 5134 562184
rect 4894 561856 4950 561912
rect 5354 561992 5410 562048
rect 243818 562400 243874 562456
rect 253846 560360 253902 560416
rect 325698 560904 325754 560960
rect 325698 560632 325754 560688
rect 345018 560768 345074 560824
rect 344926 560632 344982 560688
rect 357346 560768 357402 560824
rect 357346 560496 357402 560552
rect 365718 700304 365774 700360
rect 367006 560768 367062 560824
rect 367006 560496 367062 560552
rect 580170 697992 580226 698048
rect 494886 686024 494942 686080
rect 494242 685888 494298 685944
rect 580170 686296 580226 686352
rect 580170 674600 580226 674656
rect 372250 560088 372306 560144
rect 580170 651072 580226 651128
rect 580170 639376 580226 639432
rect 580170 627680 580226 627736
rect 580170 604152 580226 604208
rect 580170 592456 580226 592512
rect 580170 580760 580226 580816
rect 404358 562808 404414 562864
rect 386234 560904 386290 560960
rect 386234 560496 386290 560552
rect 386418 560496 386474 560552
rect 386510 560360 386566 560416
rect 385130 559952 385186 560008
rect 389086 560088 389142 560144
rect 291566 559816 291622 559872
rect 296626 559816 296682 559872
rect 304262 559816 304318 559872
rect 240138 559444 240140 559464
rect 240140 559444 240192 559464
rect 240192 559444 240194 559464
rect 240138 559408 240194 559444
rect 252650 559544 252706 559600
rect 277306 559544 277362 559600
rect 231030 559272 231086 559328
rect 232870 559272 232926 559328
rect 234618 559272 234674 559328
rect 236734 559272 236790 559328
rect 238206 559272 238262 559328
rect 248786 559272 248842 559328
rect 252558 559272 252614 559328
rect 296626 559544 296682 559600
rect 369858 559544 369914 559600
rect 304262 559408 304318 559464
rect 395802 560360 395858 560416
rect 395986 560360 396042 560416
rect 400218 560788 400274 560824
rect 400218 560768 400220 560788
rect 400220 560768 400272 560788
rect 400272 560768 400274 560788
rect 398930 560496 398986 560552
rect 398746 560360 398802 560416
rect 400218 560380 400274 560416
rect 400218 560360 400220 560380
rect 400220 560360 400272 560380
rect 400272 560360 400274 560380
rect 400218 560244 400274 560280
rect 400218 560224 400220 560244
rect 400220 560224 400272 560244
rect 400272 560224 400274 560244
rect 400218 560108 400274 560144
rect 400218 560088 400220 560108
rect 400220 560088 400272 560108
rect 400272 560088 400274 560108
rect 400218 559972 400274 560008
rect 400586 560788 400642 560824
rect 400586 560768 400588 560788
rect 400588 560768 400640 560788
rect 400640 560768 400642 560788
rect 400586 560380 400642 560416
rect 400586 560360 400588 560380
rect 400588 560360 400640 560380
rect 400640 560360 400642 560380
rect 400586 560244 400642 560280
rect 400586 560224 400588 560244
rect 400588 560224 400640 560244
rect 400640 560224 400642 560244
rect 400586 560108 400642 560144
rect 400586 560088 400588 560108
rect 400588 560088 400640 560108
rect 400640 560088 400642 560108
rect 400218 559952 400220 559972
rect 400220 559952 400272 559972
rect 400272 559952 400274 559972
rect 400586 559972 400642 560008
rect 405738 560496 405794 560552
rect 405830 560360 405886 560416
rect 411258 560360 411314 560416
rect 415950 562672 416006 562728
rect 441066 562672 441122 562728
rect 419814 562264 419870 562320
rect 423678 562128 423734 562184
rect 425610 561992 425666 562048
rect 424322 560768 424378 560824
rect 429474 561856 429530 561912
rect 437202 561720 437258 561776
rect 431866 560768 431922 560824
rect 431866 560496 431922 560552
rect 400586 559952 400588 559972
rect 400588 559952 400640 559972
rect 400640 559952 400642 559972
rect 400310 559852 400312 559872
rect 400312 559852 400364 559872
rect 400364 559852 400366 559872
rect 400310 559816 400366 559852
rect 400678 559852 400680 559872
rect 400680 559852 400732 559872
rect 400732 559852 400734 559872
rect 400678 559816 400734 559852
rect 409878 559852 409880 559872
rect 409880 559852 409932 559872
rect 409932 559852 409934 559872
rect 409878 559816 409934 559852
rect 419354 559852 419356 559872
rect 419356 559852 419408 559872
rect 419408 559852 419410 559872
rect 419354 559816 419410 559852
rect 394054 559544 394110 559600
rect 405922 559544 405978 559600
rect 277306 559272 277362 559328
rect 291566 559272 291622 559328
rect 361302 559272 361358 559328
rect 361486 559272 361542 559328
rect 383198 559272 383254 559328
rect 434626 559408 434682 559464
rect 394054 559272 394110 559328
rect 442814 559408 442870 559464
rect 434626 559272 434682 559328
rect 444562 559272 444618 559328
rect 446586 559272 446642 559328
rect 448518 559272 448574 559328
rect 580538 562536 580594 562592
rect 580354 562400 580410 562456
rect 10322 337320 10378 337376
rect 4066 8200 4122 8256
rect 3974 7520 4030 7576
rect 4066 7112 4122 7168
rect 6458 3304 6514 3360
rect 55218 6160 55274 6216
rect 138018 337184 138074 337240
rect 147586 337184 147642 337240
rect 157338 337184 157394 337240
rect 166906 337184 166962 337240
rect 176658 337184 176714 337240
rect 186226 337184 186282 337240
rect 195978 337184 196034 337240
rect 205546 337184 205602 337240
rect 215298 337184 215354 337240
rect 224866 337184 224922 337240
rect 132590 8880 132646 8936
rect 205086 4800 205142 4856
rect 229374 298016 229430 298072
rect 229558 298016 229614 298072
rect 229282 240080 229338 240136
rect 229558 240080 229614 240136
rect 229282 202852 229284 202872
rect 229284 202852 229336 202872
rect 229336 202852 229338 202872
rect 229282 202816 229338 202852
rect 229558 202816 229614 202872
rect 229282 183504 229338 183560
rect 229558 183504 229614 183560
rect 229282 144880 229338 144936
rect 229558 144880 229614 144936
rect 229282 125568 229338 125624
rect 229558 125568 229614 125624
rect 229374 22208 229430 22264
rect 229374 17992 229430 18048
rect 231766 337320 231822 337376
rect 230570 7520 230626 7576
rect 232134 3304 232190 3360
rect 234618 277344 234674 277400
rect 234802 277344 234858 277400
rect 235078 240080 235134 240136
rect 235262 240080 235318 240136
rect 234894 220768 234950 220824
rect 235170 220768 235226 220824
rect 234894 211112 234950 211168
rect 235170 211112 235226 211168
rect 234894 162832 234950 162888
rect 235078 162832 235134 162888
rect 235078 143656 235134 143712
rect 235170 143520 235226 143576
rect 234802 85720 234858 85776
rect 234802 85584 234858 85640
rect 239034 296656 239090 296712
rect 239310 296656 239366 296712
rect 240230 278704 240286 278760
rect 240414 278704 240470 278760
rect 240230 259392 240286 259448
rect 240414 259392 240470 259448
rect 239126 240116 239128 240136
rect 239128 240116 239180 240136
rect 239180 240116 239182 240136
rect 239126 240080 239182 240116
rect 240230 240080 240286 240136
rect 240414 240080 240470 240136
rect 239218 239944 239274 240000
rect 239126 220804 239128 220824
rect 239128 220804 239180 220824
rect 239180 220804 239182 220824
rect 239126 220768 239182 220804
rect 240230 220768 240286 220824
rect 240414 220768 240470 220824
rect 239034 220632 239090 220688
rect 240230 211112 240286 211168
rect 240414 211112 240470 211168
rect 240414 173884 240416 173904
rect 240416 173884 240468 173904
rect 240468 173884 240470 173904
rect 240414 173848 240470 173884
rect 240598 173848 240654 173904
rect 239126 164192 239182 164248
rect 239310 164192 239366 164248
rect 238666 32544 238722 32600
rect 238666 29144 238722 29200
rect 240046 91160 240102 91216
rect 240046 87080 240102 87136
rect 240414 18128 240470 18184
rect 240322 17992 240378 18048
rect 241610 106256 241666 106312
rect 241610 17992 241666 18048
rect 241886 278704 241942 278760
rect 242070 278704 242126 278760
rect 241886 259392 241942 259448
rect 242070 259392 242126 259448
rect 241886 240080 241942 240136
rect 242070 240080 242126 240136
rect 241886 220768 241942 220824
rect 242070 220768 242126 220824
rect 241886 211112 241942 211168
rect 242070 211112 242126 211168
rect 241794 106256 241850 106312
rect 241794 18128 241850 18184
rect 244094 202816 244150 202872
rect 244278 202816 244334 202872
rect 244094 135224 244150 135280
rect 244278 135224 244334 135280
rect 245750 231784 245806 231840
rect 245934 231784 245990 231840
rect 245750 144880 245806 144936
rect 245934 144880 245990 144936
rect 245750 125568 245806 125624
rect 245934 125568 245990 125624
rect 249706 29280 249762 29336
rect 249706 28872 249762 28928
rect 250166 335280 250222 335336
rect 250258 335144 250314 335200
rect 249982 325624 250038 325680
rect 250258 325624 250314 325680
rect 249982 6160 250038 6216
rect 251178 288360 251234 288416
rect 251178 219408 251234 219464
rect 251178 143520 251234 143576
rect 251178 133900 251180 133920
rect 251180 133900 251232 133920
rect 251232 133900 251234 133920
rect 251178 133864 251234 133900
rect 251178 85584 251234 85640
rect 251362 288360 251418 288416
rect 251362 219408 251418 219464
rect 251546 200096 251602 200152
rect 251730 200096 251786 200152
rect 251454 182280 251510 182336
rect 251638 182008 251694 182064
rect 251454 172508 251510 172544
rect 251454 172488 251456 172508
rect 251456 172488 251508 172508
rect 251508 172488 251510 172508
rect 251638 172488 251694 172544
rect 251362 143540 251418 143576
rect 251362 143520 251364 143540
rect 251364 143520 251416 143540
rect 251416 143520 251418 143540
rect 251362 105032 251418 105088
rect 251454 104896 251510 104952
rect 251362 85584 251418 85640
rect 251454 56752 251510 56808
rect 251454 56480 251510 56536
rect 251362 8336 251418 8392
rect 251546 8336 251602 8392
rect 253938 306312 253994 306368
rect 253754 87080 253810 87136
rect 253938 87080 253994 87136
rect 254122 306312 254178 306368
rect 254214 241440 254270 241496
rect 254398 241440 254454 241496
rect 254214 222128 254270 222184
rect 254398 222128 254454 222184
rect 254214 191800 254270 191856
rect 254398 191800 254454 191856
rect 254214 154536 254270 154592
rect 254398 154536 254454 154592
rect 254214 135224 254270 135280
rect 254398 135224 254454 135280
rect 255318 143520 255374 143576
rect 255594 251096 255650 251152
rect 255778 251096 255834 251152
rect 255686 191936 255742 191992
rect 255594 191820 255650 191856
rect 255594 191800 255596 191820
rect 255596 191800 255648 191820
rect 255648 191800 255650 191820
rect 255502 143520 255558 143576
rect 260746 134136 260802 134192
rect 261206 211112 261262 211168
rect 261390 211112 261446 211168
rect 261390 125704 261446 125760
rect 261298 125568 261354 125624
rect 262494 144880 262550 144936
rect 262678 144880 262734 144936
rect 267278 270680 267334 270736
rect 267002 270544 267058 270600
rect 267002 269048 267058 269104
rect 267186 269048 267242 269104
rect 267002 164192 267058 164248
rect 267278 164056 267334 164112
rect 267002 154536 267058 154592
rect 267278 154536 267334 154592
rect 267002 19216 267058 19272
rect 267278 19080 267334 19136
rect 269118 134156 269174 134192
rect 269118 134136 269120 134156
rect 269120 134136 269172 134156
rect 269172 134136 269174 134156
rect 270498 180820 270500 180840
rect 270500 180820 270552 180840
rect 270552 180820 270554 180840
rect 270498 180784 270554 180820
rect 270498 40332 270500 40352
rect 270500 40332 270552 40352
rect 270552 40332 270554 40352
rect 270498 40296 270554 40332
rect 270498 29180 270500 29200
rect 270500 29180 270552 29200
rect 270552 29180 270554 29200
rect 270498 29144 270554 29180
rect 272982 63824 273038 63880
rect 273166 63824 273222 63880
rect 273902 337320 273958 337376
rect 273994 29280 274050 29336
rect 275374 181056 275430 181112
rect 275374 134000 275430 134056
rect 278962 8880 279018 8936
rect 280526 40332 280528 40352
rect 280528 40332 280580 40352
rect 280580 40332 280582 40352
rect 280526 40296 280582 40332
rect 282734 134000 282790 134056
rect 282918 134000 282974 134056
rect 282826 87236 282882 87272
rect 282826 87216 282828 87236
rect 282828 87216 282880 87236
rect 282880 87216 282882 87236
rect 284942 29280 284998 29336
rect 284942 29008 284998 29064
rect 287334 222128 287390 222184
rect 287518 222128 287574 222184
rect 287334 202816 287390 202872
rect 287518 202816 287574 202872
rect 287242 124208 287298 124264
rect 287518 124208 287574 124264
rect 287334 67632 287390 67688
rect 287426 67496 287482 67552
rect 287242 28872 287298 28928
rect 287334 28736 287390 28792
rect 288806 299376 288862 299432
rect 288990 299376 289046 299432
rect 290186 135360 290242 135416
rect 290094 135224 290150 135280
rect 291474 278704 291530 278760
rect 291658 278704 291714 278760
rect 291566 230460 291568 230480
rect 291568 230460 291620 230480
rect 291620 230460 291622 230480
rect 291566 230424 291622 230460
rect 291750 230424 291806 230480
rect 291382 183504 291438 183560
rect 291566 183504 291622 183560
rect 291474 173884 291476 173904
rect 291476 173884 291528 173904
rect 291528 173884 291530 173904
rect 291474 173848 291530 173884
rect 291750 173848 291806 173904
rect 291566 164192 291622 164248
rect 291750 164192 291806 164248
rect 291566 154672 291622 154728
rect 291658 154400 291714 154456
rect 291566 135360 291622 135416
rect 291566 135088 291622 135144
rect 291566 102040 291622 102096
rect 291474 101904 291530 101960
rect 291842 29552 291898 29608
rect 291842 29008 291898 29064
rect 292762 87236 292818 87272
rect 292762 87216 292764 87236
rect 292764 87216 292816 87236
rect 292816 87216 292818 87236
rect 297546 40296 297602 40352
rect 297546 40024 297602 40080
rect 299754 35944 299810 36000
rect 299938 35944 299994 36000
rect 304998 113192 305054 113248
rect 305274 278704 305330 278760
rect 305550 278704 305606 278760
rect 305274 113192 305330 113248
rect 306286 29416 306342 29472
rect 306286 29144 306342 29200
rect 305182 15136 305238 15192
rect 305366 15136 305422 15192
rect 306378 4800 306434 4856
rect 308034 212508 308036 212528
rect 308036 212508 308088 212528
rect 308088 212508 308090 212528
rect 308034 212472 308090 212508
rect 308218 212472 308274 212528
rect 308034 193196 308036 193216
rect 308036 193196 308088 193216
rect 308088 193196 308090 193216
rect 308034 193160 308090 193196
rect 308310 193160 308366 193216
rect 309046 181076 309102 181112
rect 309046 181056 309048 181076
rect 309048 181056 309100 181076
rect 309100 181056 309102 181076
rect 309046 134000 309102 134056
rect 309046 133728 309102 133784
rect 307942 86944 307998 87000
rect 308126 86944 308182 87000
rect 307942 44104 307998 44160
rect 308218 44104 308274 44160
rect 310150 328480 310206 328536
rect 309414 328344 309470 328400
rect 309322 201476 309378 201512
rect 309322 201456 309324 201476
rect 309324 201456 309376 201476
rect 309376 201456 309378 201476
rect 309506 201456 309562 201512
rect 310426 180784 310482 180840
rect 310794 315968 310850 316024
rect 310886 315832 310942 315888
rect 310702 229064 310758 229120
rect 310978 229064 311034 229120
rect 310794 180784 310850 180840
rect 311070 93880 311126 93936
rect 310978 93744 311034 93800
rect 312082 181076 312138 181112
rect 312082 181056 312084 181076
rect 312084 181056 312136 181076
rect 312136 181056 312138 181076
rect 314014 328480 314070 328536
rect 313738 328344 313794 328400
rect 313462 315968 313518 316024
rect 313646 315968 313702 316024
rect 315946 29144 316002 29200
rect 315946 29008 316002 29064
rect 316314 201456 316370 201512
rect 316498 201456 316554 201512
rect 317510 134020 317566 134056
rect 317510 134000 317512 134020
rect 317512 134000 317564 134020
rect 317564 134000 317566 134020
rect 325146 338272 325202 338328
rect 324594 338136 324650 338192
rect 324594 251096 324650 251152
rect 324778 251096 324834 251152
rect 324594 231820 324596 231840
rect 324596 231820 324648 231840
rect 324648 231820 324650 231840
rect 324594 231784 324650 231820
rect 324870 231820 324872 231840
rect 324872 231820 324924 231840
rect 324924 231820 324926 231840
rect 324870 231784 324926 231820
rect 324502 172488 324558 172544
rect 324686 172488 324742 172544
rect 324594 144880 324650 144936
rect 324778 144880 324834 144936
rect 324778 135360 324834 135416
rect 324594 135224 324650 135280
rect 324686 115912 324742 115968
rect 324870 115912 324926 115968
rect 325606 29552 325662 29608
rect 325606 29280 325662 29336
rect 326986 181328 327042 181384
rect 326986 181056 327042 181112
rect 326986 133864 327042 133920
rect 326986 87216 327042 87272
rect 326986 86944 327042 87000
rect 326802 63724 326804 63744
rect 326804 63724 326856 63744
rect 326856 63724 326858 63744
rect 326802 63688 326858 63724
rect 327354 278704 327410 278760
rect 327630 278704 327686 278760
rect 327354 230424 327410 230480
rect 327538 230424 327594 230480
rect 327354 201456 327410 201512
rect 327538 201456 327594 201512
rect 327446 138216 327502 138272
rect 327354 135244 327410 135280
rect 327354 135224 327356 135244
rect 327356 135224 327408 135244
rect 327408 135224 327410 135244
rect 327262 133900 327264 133920
rect 327264 133900 327316 133920
rect 327316 133900 327318 133920
rect 327262 133864 327318 133900
rect 327538 106392 327594 106448
rect 327446 106256 327502 106312
rect 328458 125588 328514 125624
rect 328458 125568 328460 125588
rect 328460 125568 328512 125588
rect 328512 125568 328514 125588
rect 328366 40568 328422 40624
rect 328366 40160 328422 40216
rect 328734 125568 328790 125624
rect 332322 337320 332378 337376
rect 335266 63824 335322 63880
rect 336646 134136 336702 134192
rect 336646 87216 336702 87272
rect 336646 86944 336702 87000
rect 336922 48184 336978 48240
rect 337014 48048 337070 48104
rect 337934 40568 337990 40624
rect 337934 40024 337990 40080
rect 342350 241440 342406 241496
rect 342534 241440 342590 241496
rect 342350 222128 342406 222184
rect 342534 222128 342590 222184
rect 342350 193160 342406 193216
rect 342534 193160 342590 193216
rect 343914 172488 343970 172544
rect 344098 172488 344154 172544
rect 342534 164328 342590 164384
rect 343914 164328 343970 164384
rect 342534 164192 342590 164248
rect 343914 164192 343970 164248
rect 342534 114552 342590 114608
rect 342718 114552 342774 114608
rect 345294 251368 345350 251424
rect 345202 251232 345258 251288
rect 345018 172488 345074 172544
rect 345294 172488 345350 172544
rect 347778 280200 347834 280256
rect 347962 280200 348018 280256
rect 347962 231784 348018 231840
rect 348146 231784 348202 231840
rect 347962 212472 348018 212528
rect 348146 212472 348202 212528
rect 347962 193160 348018 193216
rect 348146 193160 348202 193216
rect 347962 173848 348018 173904
rect 348146 173848 348202 173904
rect 347962 164192 348018 164248
rect 348146 164192 348202 164248
rect 347962 144880 348018 144936
rect 348146 144880 348202 144936
rect 347962 125588 348018 125624
rect 347962 125568 347964 125588
rect 347964 125568 348016 125588
rect 348016 125568 348018 125588
rect 348146 125568 348202 125624
rect 347962 106276 348018 106312
rect 347962 106256 347964 106276
rect 347964 106256 348016 106276
rect 348016 106256 348018 106276
rect 348146 106256 348202 106312
rect 348330 63960 348386 64016
rect 348330 63688 348386 63744
rect 347962 45464 348018 45520
rect 348054 45328 348110 45384
rect 348054 26152 348110 26208
rect 348238 26152 348294 26208
rect 348054 24792 348110 24848
rect 348238 24792 348294 24848
rect 356058 87116 356060 87136
rect 356060 87116 356112 87136
rect 356112 87116 356114 87136
rect 356058 87080 356114 87116
rect 356058 40160 356114 40216
rect 357438 134036 357440 134056
rect 357440 134036 357492 134056
rect 357492 134036 357494 134056
rect 357438 134000 357494 134036
rect 359554 63708 359610 63744
rect 359554 63688 359556 63708
rect 359556 63688 359608 63708
rect 359608 63688 359610 63708
rect 360014 16788 360070 16824
rect 360014 16768 360016 16788
rect 360016 16768 360068 16788
rect 360068 16768 360070 16788
rect 361118 134036 361120 134056
rect 361120 134036 361172 134056
rect 361172 134036 361174 134056
rect 361118 134000 361174 134036
rect 361118 16788 361174 16824
rect 361118 16768 361120 16788
rect 361120 16768 361172 16788
rect 361172 16768 361174 16788
rect 362130 181464 362186 181520
rect 362130 180784 362186 180840
rect 362958 241440 363014 241496
rect 363142 241440 363198 241496
rect 362958 222128 363014 222184
rect 363142 222128 363198 222184
rect 362958 202816 363014 202872
rect 363142 202816 363198 202872
rect 362958 183504 363014 183560
rect 363142 183504 363198 183560
rect 362958 154536 363014 154592
rect 363234 154536 363290 154592
rect 362958 135224 363014 135280
rect 363234 135224 363290 135280
rect 362958 115912 363014 115968
rect 363234 115912 363290 115968
rect 362958 96600 363014 96656
rect 363234 96600 363290 96656
rect 365626 87352 365682 87408
rect 365626 63552 365682 63608
rect 365626 40060 365628 40080
rect 365628 40060 365680 40080
rect 365680 40060 365682 40080
rect 365626 40024 365682 40060
rect 398470 180956 398472 180976
rect 398472 180956 398524 180976
rect 398524 180956 398526 180976
rect 398470 180920 398526 180956
rect 398470 134036 398472 134056
rect 398472 134036 398524 134056
rect 398524 134036 398526 134056
rect 398470 134000 398526 134036
rect 398470 87100 398526 87136
rect 398470 87080 398472 87100
rect 398472 87080 398524 87100
rect 398524 87080 398526 87100
rect 398470 63724 398472 63744
rect 398472 63724 398524 63744
rect 398524 63724 398526 63744
rect 398470 63688 398526 63724
rect 398470 40196 398472 40216
rect 398472 40196 398524 40216
rect 398524 40196 398526 40216
rect 398470 40160 398526 40196
rect 398470 29180 398472 29200
rect 398472 29180 398524 29200
rect 398524 29180 398526 29200
rect 398470 29144 398526 29180
rect 398470 16804 398472 16824
rect 398472 16804 398524 16824
rect 398524 16804 398526 16824
rect 398470 16768 398526 16804
rect 399022 180956 399024 180976
rect 399024 180956 399076 180976
rect 399076 180956 399078 180976
rect 399022 180920 399078 180956
rect 399022 134036 399024 134056
rect 399024 134036 399076 134056
rect 399076 134036 399078 134056
rect 399022 134000 399078 134036
rect 398838 87100 398894 87136
rect 398838 87080 398840 87100
rect 398840 87080 398892 87100
rect 398892 87080 398894 87100
rect 399022 63724 399024 63744
rect 399024 63724 399076 63744
rect 399076 63724 399078 63744
rect 399022 63688 399078 63724
rect 399022 40196 399024 40216
rect 399024 40196 399076 40216
rect 399076 40196 399078 40216
rect 399022 40160 399078 40196
rect 399022 29180 399024 29200
rect 399024 29180 399076 29200
rect 399076 29180 399078 29200
rect 399022 29144 399078 29180
rect 399022 16804 399024 16824
rect 399024 16804 399076 16824
rect 399076 16804 399078 16824
rect 399022 16768 399078 16804
rect 417882 180956 417884 180976
rect 417884 180956 417936 180976
rect 417936 180956 417938 180976
rect 417882 180920 417938 180956
rect 417882 134036 417884 134056
rect 417884 134036 417936 134056
rect 417936 134036 417938 134056
rect 417882 134000 417938 134036
rect 417882 87116 417884 87136
rect 417884 87116 417936 87136
rect 417936 87116 417938 87136
rect 417882 87080 417938 87116
rect 417882 63708 417938 63744
rect 417882 63688 417884 63708
rect 417884 63688 417936 63708
rect 417936 63688 417938 63708
rect 417882 40196 417884 40216
rect 417884 40196 417936 40216
rect 417936 40196 417938 40216
rect 417882 40160 417938 40196
rect 417882 29164 417938 29200
rect 417882 29144 417884 29164
rect 417884 29144 417936 29164
rect 417936 29144 417938 29164
rect 417882 16768 417938 16824
rect 417882 16360 417938 16416
rect 418342 180956 418344 180976
rect 418344 180956 418396 180976
rect 418396 180956 418398 180976
rect 418342 180920 418398 180956
rect 418342 134036 418344 134056
rect 418344 134036 418396 134056
rect 418396 134036 418398 134056
rect 418342 134000 418398 134036
rect 418342 87116 418344 87136
rect 418344 87116 418396 87136
rect 418396 87116 418398 87136
rect 418342 87080 418398 87116
rect 418342 40196 418344 40216
rect 418344 40196 418396 40216
rect 418396 40196 418398 40216
rect 418342 40160 418398 40196
rect 418158 29164 418214 29200
rect 418158 29144 418160 29164
rect 418160 29144 418212 29164
rect 418212 29144 418214 29164
rect 419630 63708 419686 63744
rect 419630 63688 419632 63708
rect 419632 63688 419684 63708
rect 419684 63688 419686 63708
rect 425150 87216 425206 87272
rect 425058 86944 425114 87000
rect 425058 16668 425060 16688
rect 425060 16668 425112 16688
rect 425112 16668 425114 16688
rect 425058 16632 425114 16668
rect 434994 337864 435050 337920
rect 434350 299376 434406 299432
rect 434350 289856 434406 289912
rect 434350 280064 434406 280120
rect 434350 270544 434406 270600
rect 434350 260752 434406 260808
rect 434350 251232 434406 251288
rect 434350 173848 434406 173904
rect 434442 164192 434498 164248
rect 434534 143520 434590 143576
rect 435178 212472 435234 212528
rect 435362 212472 435418 212528
rect 435178 202816 435234 202872
rect 435362 202816 435418 202872
rect 434718 143520 434774 143576
rect 434258 48184 434314 48240
rect 434442 41248 434498 41304
rect 435178 87080 435234 87136
rect 435178 86944 435234 87000
rect 434626 16904 434682 16960
rect 438214 337864 438270 337920
rect 443918 183504 443974 183560
rect 444102 183504 444158 183560
rect 444378 86980 444380 87000
rect 444380 86980 444432 87000
rect 444432 86980 444434 87000
rect 444378 86944 444434 86980
rect 444378 29044 444380 29064
rect 444380 29044 444432 29064
rect 444432 29044 444434 29064
rect 444378 29008 444434 29044
rect 444378 16668 444380 16688
rect 444380 16668 444432 16688
rect 444432 16668 444434 16688
rect 444378 16632 444434 16668
rect 448150 337728 448206 337784
rect 449162 337728 449218 337784
rect 447230 134272 447286 134328
rect 447138 134000 447194 134056
rect 447230 63960 447286 64016
rect 447138 63688 447194 63744
rect 447230 40432 447286 40488
rect 447138 40160 447194 40216
rect 447230 16904 447286 16960
rect 449530 337320 449586 337376
rect 449254 87216 449310 87272
rect 449254 29280 449310 29336
rect 449806 4800 449862 4856
rect 454406 180940 454462 180976
rect 454406 180920 454408 180940
rect 454408 180920 454460 180940
rect 454460 180920 454462 180940
rect 458362 180940 458418 180976
rect 458362 180920 458364 180940
rect 458364 180920 458416 180940
rect 458416 180920 458418 180940
rect 460846 134544 460902 134600
rect 460846 134136 460902 134192
rect 463606 87488 463662 87544
rect 463606 87080 463662 87136
rect 460846 64232 460902 64288
rect 460846 63824 460902 63880
rect 460846 40704 460902 40760
rect 460846 40296 460902 40352
rect 463790 86980 463792 87000
rect 463792 86980 463844 87000
rect 463844 86980 463846 87000
rect 463790 86944 463846 86980
rect 466550 86980 466552 87000
rect 466552 86980 466604 87000
rect 466604 86980 466606 87000
rect 466550 86944 466606 86980
rect 471886 29416 471942 29472
rect 476026 29180 476028 29200
rect 476028 29180 476080 29200
rect 476080 29180 476082 29200
rect 476026 29144 476082 29180
rect 471886 29008 471942 29064
rect 471886 17040 471942 17096
rect 476026 16804 476028 16824
rect 476028 16804 476080 16824
rect 476080 16804 476082 16824
rect 476026 16768 476082 16804
rect 471886 16632 471942 16688
rect 482926 29280 482982 29336
rect 482926 16904 482982 16960
rect 530582 337320 530638 337376
rect 579710 557232 579766 557288
rect 579802 545536 579858 545592
rect 579802 533840 579858 533896
rect 579802 510312 579858 510368
rect 579802 498616 579858 498672
rect 579802 463392 579858 463448
rect 579802 451696 579858 451752
rect 579802 439864 579858 439920
rect 579802 416472 579858 416528
rect 579802 404776 579858 404832
rect 579802 392944 579858 393000
rect 579802 369552 579858 369608
rect 579894 357856 579950 357912
rect 579894 346024 579950 346080
rect 579894 322632 579950 322688
rect 579986 310800 580042 310856
rect 579894 299104 579950 299160
rect 580078 275712 580134 275768
rect 580170 263880 580226 263936
rect 580906 252184 580962 252240
rect 580814 228792 580870 228848
rect 580722 216960 580778 217016
rect 580630 170040 580686 170096
rect 580538 158344 580594 158400
rect 580446 123120 580502 123176
rect 580354 111424 580410 111480
rect 580262 76200 580318 76256
rect 579802 4800 579858 4856
<< metal3 >>
rect 8109 700362 8175 700365
rect 365713 700362 365779 700365
rect 8109 700360 365779 700362
rect 8109 700304 8114 700360
rect 8170 700304 365718 700360
rect 365774 700304 365779 700360
rect 8109 700302 365779 700304
rect 8109 700299 8175 700302
rect 365713 700299 365779 700302
rect 580165 698050 580231 698053
rect 583520 698050 584960 698140
rect 580165 698048 584960 698050
rect 580165 697992 580170 698048
rect 580226 697992 584960 698048
rect 580165 697990 584960 697992
rect 580165 697987 580231 697990
rect 583520 697900 584960 697990
rect -960 696540 480 696780
rect 580165 686354 580231 686357
rect 583520 686354 584960 686444
rect 580165 686352 584960 686354
rect 580165 686296 580170 686352
rect 580226 686296 584960 686352
rect 580165 686294 584960 686296
rect 580165 686291 580231 686294
rect 583520 686204 584960 686294
rect 494881 686082 494947 686085
rect 494102 686080 494947 686082
rect 494102 686024 494886 686080
rect 494942 686024 494947 686080
rect 494102 686022 494947 686024
rect 494102 685946 494162 686022
rect 494881 686019 494947 686022
rect 494237 685946 494303 685949
rect 494102 685944 494303 685946
rect 494102 685888 494242 685944
rect 494298 685888 494303 685944
rect 494102 685886 494303 685888
rect 494237 685883 494303 685886
rect -960 682274 480 682364
rect 3509 682274 3575 682277
rect -960 682272 3575 682274
rect -960 682216 3514 682272
rect 3570 682216 3575 682272
rect -960 682214 3575 682216
rect -960 682124 480 682214
rect 3509 682211 3575 682214
rect 580165 674658 580231 674661
rect 583520 674658 584960 674748
rect 580165 674656 584960 674658
rect 580165 674600 580170 674656
rect 580226 674600 584960 674656
rect 580165 674598 584960 674600
rect 580165 674595 580231 674598
rect 583520 674508 584960 674598
rect -960 667994 480 668084
rect 3417 667994 3483 667997
rect -960 667992 3483 667994
rect -960 667936 3422 667992
rect 3478 667936 3483 667992
rect -960 667934 3483 667936
rect -960 667844 480 667934
rect 3417 667931 3483 667934
rect 583520 662676 584960 662916
rect -960 653578 480 653668
rect 3049 653578 3115 653581
rect -960 653576 3115 653578
rect -960 653520 3054 653576
rect 3110 653520 3115 653576
rect -960 653518 3115 653520
rect -960 653428 480 653518
rect 3049 653515 3115 653518
rect 580165 651130 580231 651133
rect 583520 651130 584960 651220
rect 580165 651128 584960 651130
rect 580165 651072 580170 651128
rect 580226 651072 584960 651128
rect 580165 651070 584960 651072
rect 580165 651067 580231 651070
rect 583520 650980 584960 651070
rect 580165 639434 580231 639437
rect 583520 639434 584960 639524
rect 580165 639432 584960 639434
rect 580165 639376 580170 639432
rect 580226 639376 584960 639432
rect 580165 639374 584960 639376
rect 580165 639371 580231 639374
rect 583520 639284 584960 639374
rect -960 639012 480 639252
rect 580165 627738 580231 627741
rect 583520 627738 584960 627828
rect 580165 627736 584960 627738
rect 580165 627680 580170 627736
rect 580226 627680 584960 627736
rect 580165 627678 584960 627680
rect 580165 627675 580231 627678
rect 583520 627588 584960 627678
rect -960 624882 480 624972
rect 3417 624882 3483 624885
rect -960 624880 3483 624882
rect -960 624824 3422 624880
rect 3478 624824 3483 624880
rect -960 624822 3483 624824
rect -960 624732 480 624822
rect 3417 624819 3483 624822
rect 583520 615756 584960 615996
rect -960 610466 480 610556
rect 3417 610466 3483 610469
rect -960 610464 3483 610466
rect -960 610408 3422 610464
rect 3478 610408 3483 610464
rect -960 610406 3483 610408
rect -960 610316 480 610406
rect 3417 610403 3483 610406
rect 580165 604210 580231 604213
rect 583520 604210 584960 604300
rect 580165 604208 584960 604210
rect 580165 604152 580170 604208
rect 580226 604152 584960 604208
rect 580165 604150 584960 604152
rect 580165 604147 580231 604150
rect 583520 604060 584960 604150
rect -960 596050 480 596140
rect 3233 596050 3299 596053
rect -960 596048 3299 596050
rect -960 595992 3238 596048
rect 3294 595992 3299 596048
rect -960 595990 3299 595992
rect -960 595900 480 595990
rect 3233 595987 3299 595990
rect 580165 592514 580231 592517
rect 583520 592514 584960 592604
rect 580165 592512 584960 592514
rect 580165 592456 580170 592512
rect 580226 592456 584960 592512
rect 580165 592454 584960 592456
rect 580165 592451 580231 592454
rect 583520 592364 584960 592454
rect -960 581620 480 581860
rect 580165 580818 580231 580821
rect 583520 580818 584960 580908
rect 580165 580816 584960 580818
rect 580165 580760 580170 580816
rect 580226 580760 584960 580816
rect 580165 580758 584960 580760
rect 580165 580755 580231 580758
rect 583520 580668 584960 580758
rect 583520 568836 584960 569076
rect -960 567354 480 567444
rect 3417 567354 3483 567357
rect -960 567352 3483 567354
rect -960 567296 3422 567352
rect 3478 567296 3483 567352
rect -960 567294 3483 567296
rect -960 567204 480 567294
rect 3417 567291 3483 567294
rect 357382 563076 357388 563140
rect 357452 563138 357458 563140
rect 366950 563138 366956 563140
rect 357452 563078 366956 563138
rect 357452 563076 357458 563078
rect 366950 563076 366956 563078
rect 367020 563076 367026 563140
rect 237782 562940 237788 563004
rect 237852 563002 237858 563004
rect 249977 563002 250043 563005
rect 237852 563000 250043 563002
rect 237852 562944 249982 563000
rect 250038 562944 250043 563000
rect 237852 562942 250043 562944
rect 237852 562940 237858 562942
rect 249977 562939 250043 562942
rect 252502 562940 252508 563004
rect 252572 563002 252578 563004
rect 253606 563002 253612 563004
rect 252572 562942 253612 563002
rect 252572 562940 252578 562942
rect 253606 562940 253612 562942
rect 253676 562940 253682 563004
rect 266302 562940 266308 563004
rect 266372 563002 266378 563004
rect 275870 563002 275876 563004
rect 266372 562942 275876 563002
rect 266372 562940 266378 562942
rect 275870 562940 275876 562942
rect 275940 562940 275946 563004
rect 288617 563002 288683 563005
rect 446254 563002 446260 563004
rect 288617 563000 446260 563002
rect 288617 562944 288622 563000
rect 288678 562944 446260 563000
rect 288617 562942 446260 562944
rect 288617 562939 288683 562942
rect 446254 562940 446260 562942
rect 446324 562940 446330 563004
rect 236862 562804 236868 562868
rect 236932 562866 236938 562868
rect 404353 562866 404419 562869
rect 236932 562864 404419 562866
rect 236932 562808 404358 562864
rect 404414 562808 404419 562864
rect 236932 562806 404419 562808
rect 236932 562804 236938 562806
rect 404353 562803 404419 562806
rect 4153 562730 4219 562733
rect 5206 562730 5212 562732
rect 4153 562728 5212 562730
rect 4153 562672 4158 562728
rect 4214 562672 5212 562728
rect 4153 562670 5212 562672
rect 4153 562667 4219 562670
rect 5206 562668 5212 562670
rect 5276 562668 5282 562732
rect 125542 562668 125548 562732
rect 125612 562730 125618 562732
rect 135110 562730 135116 562732
rect 125612 562670 135116 562730
rect 125612 562668 125618 562670
rect 135110 562668 135116 562670
rect 135180 562668 135186 562732
rect 164182 562668 164188 562732
rect 164252 562730 164258 562732
rect 167310 562730 167316 562732
rect 164252 562670 167316 562730
rect 164252 562668 164258 562670
rect 167310 562668 167316 562670
rect 167380 562668 167386 562732
rect 183502 562668 183508 562732
rect 183572 562730 183578 562732
rect 193070 562730 193076 562732
rect 183572 562670 193076 562730
rect 183572 562668 183578 562670
rect 193070 562668 193076 562670
rect 193140 562668 193146 562732
rect 205030 562668 205036 562732
rect 205100 562730 205106 562732
rect 207606 562730 207612 562732
rect 205100 562670 207612 562730
rect 205100 562668 205106 562670
rect 207606 562668 207612 562670
rect 207676 562668 207682 562732
rect 236494 562668 236500 562732
rect 236564 562730 236570 562732
rect 415945 562730 416011 562733
rect 236564 562728 416011 562730
rect 236564 562672 415950 562728
rect 416006 562672 416011 562728
rect 236564 562670 416011 562672
rect 236564 562668 236570 562670
rect 415945 562667 416011 562670
rect 424358 562668 424364 562732
rect 424428 562730 424434 562732
rect 428406 562730 428412 562732
rect 424428 562670 428412 562730
rect 424428 562668 424434 562670
rect 428406 562668 428412 562670
rect 428476 562668 428482 562732
rect 436134 562668 436140 562732
rect 436204 562730 436210 562732
rect 441061 562730 441127 562733
rect 436204 562728 441127 562730
rect 436204 562672 441066 562728
rect 441122 562672 441127 562728
rect 436204 562670 441127 562672
rect 436204 562668 436210 562670
rect 441061 562667 441127 562670
rect 3969 562594 4035 562597
rect 242249 562594 242315 562597
rect 248045 562594 248111 562597
rect 580533 562594 580599 562597
rect 3969 562592 5642 562594
rect 3969 562536 3974 562592
rect 4030 562536 5642 562592
rect 3969 562534 5642 562536
rect 3969 562531 4035 562534
rect 3785 562322 3851 562325
rect 5349 562322 5415 562325
rect 3785 562320 5415 562322
rect 3785 562264 3790 562320
rect 3846 562264 5354 562320
rect 5410 562264 5415 562320
rect 3785 562262 5415 562264
rect 5582 562322 5642 562534
rect 242249 562592 244106 562594
rect 242249 562536 242254 562592
rect 242310 562536 244106 562592
rect 242249 562534 244106 562536
rect 242249 562531 242315 562534
rect 237966 562396 237972 562460
rect 238036 562458 238042 562460
rect 243813 562458 243879 562461
rect 238036 562456 243879 562458
rect 238036 562400 243818 562456
rect 243874 562400 243879 562456
rect 238036 562398 243879 562400
rect 244046 562458 244106 562534
rect 248045 562592 580599 562594
rect 248045 562536 248050 562592
rect 248106 562536 580538 562592
rect 580594 562536 580599 562592
rect 248045 562534 580599 562536
rect 248045 562531 248111 562534
rect 580533 562531 580599 562534
rect 580349 562458 580415 562461
rect 244046 562456 580415 562458
rect 244046 562400 580354 562456
rect 580410 562400 580415 562456
rect 244046 562398 580415 562400
rect 238036 562396 238042 562398
rect 243813 562395 243879 562398
rect 580349 562395 580415 562398
rect 419809 562322 419875 562325
rect 5582 562320 419875 562322
rect 5582 562264 419814 562320
rect 419870 562264 419875 562320
rect 5582 562262 419875 562264
rect 3785 562259 3851 562262
rect 5349 562259 5415 562262
rect 419809 562259 419875 562262
rect 5073 562186 5139 562189
rect 423673 562186 423739 562189
rect 5073 562184 423739 562186
rect 5073 562128 5078 562184
rect 5134 562128 423678 562184
rect 423734 562128 423739 562184
rect 5073 562126 423739 562128
rect 5073 562123 5139 562126
rect 423673 562123 423739 562126
rect 5349 562050 5415 562053
rect 425605 562050 425671 562053
rect 5349 562048 425671 562050
rect 5349 561992 5354 562048
rect 5410 561992 425610 562048
rect 425666 561992 425671 562048
rect 5349 561990 425671 561992
rect 5349 561987 5415 561990
rect 425605 561987 425671 561990
rect 4889 561914 4955 561917
rect 429469 561914 429535 561917
rect 4889 561912 429535 561914
rect 4889 561856 4894 561912
rect 4950 561856 429474 561912
rect 429530 561856 429535 561912
rect 4889 561854 429535 561856
rect 4889 561851 4955 561854
rect 429469 561851 429535 561854
rect 3601 561778 3667 561781
rect 437197 561778 437263 561781
rect 3601 561776 437263 561778
rect 3601 561720 3606 561776
rect 3662 561720 437202 561776
rect 437258 561720 437263 561776
rect 3601 561718 437263 561720
rect 3601 561715 3667 561718
rect 437197 561715 437263 561718
rect 288382 561580 288388 561644
rect 288452 561642 288458 561644
rect 293166 561642 293172 561644
rect 288452 561582 293172 561642
rect 288452 561580 288458 561582
rect 293166 561580 293172 561582
rect 293236 561580 293242 561644
rect 50470 561308 50476 561372
rect 50540 561370 50546 561372
rect 51574 561370 51580 561372
rect 50540 561310 51580 561370
rect 50540 561308 50546 561310
rect 51574 561308 51580 561310
rect 51644 561308 51650 561372
rect 85614 561308 85620 561372
rect 85684 561370 85690 561372
rect 90214 561370 90220 561372
rect 85684 561310 90220 561370
rect 85684 561308 85690 561310
rect 90214 561308 90220 561310
rect 90284 561308 90290 561372
rect 108430 561308 108436 561372
rect 108500 561370 108506 561372
rect 109718 561370 109724 561372
rect 108500 561310 109724 561370
rect 108500 561308 108506 561310
rect 109718 561308 109724 561310
rect 109788 561308 109794 561372
rect 117630 561308 117636 561372
rect 117700 561370 117706 561372
rect 120758 561370 120764 561372
rect 117700 561310 120764 561370
rect 117700 561308 117706 561310
rect 120758 561308 120764 561310
rect 120828 561308 120834 561372
rect 135662 561308 135668 561372
rect 135732 561370 135738 561372
rect 140078 561370 140084 561372
rect 135732 561310 140084 561370
rect 135732 561308 135738 561310
rect 140078 561308 140084 561310
rect 140148 561308 140154 561372
rect 147438 561308 147444 561372
rect 147508 561370 147514 561372
rect 154430 561370 154436 561372
rect 147508 561310 154436 561370
rect 147508 561308 147514 561310
rect 154430 561308 154436 561310
rect 154500 561308 154506 561372
rect 154982 561308 154988 561372
rect 155052 561370 155058 561372
rect 159398 561370 159404 561372
rect 155052 561310 159404 561370
rect 155052 561308 155058 561310
rect 159398 561308 159404 561310
rect 159468 561308 159474 561372
rect 176142 561308 176148 561372
rect 176212 561370 176218 561372
rect 178718 561370 178724 561372
rect 176212 561310 178724 561370
rect 176212 561308 176218 561310
rect 178718 561308 178724 561310
rect 178788 561308 178794 561372
rect 193622 561308 193628 561372
rect 193692 561370 193698 561372
rect 196750 561370 196756 561372
rect 193692 561310 196756 561370
rect 193692 561308 193698 561310
rect 196750 561308 196756 561310
rect 196820 561308 196826 561372
rect 223614 561308 223620 561372
rect 223684 561370 223690 561372
rect 225454 561370 225460 561372
rect 223684 561310 225460 561370
rect 223684 561308 223690 561310
rect 225454 561308 225460 561310
rect 225524 561308 225530 561372
rect 325734 561308 325740 561372
rect 325804 561370 325810 561372
rect 335118 561370 335124 561372
rect 325804 561310 335124 561370
rect 325804 561308 325810 561310
rect 335118 561308 335124 561310
rect 335188 561308 335194 561372
rect 393262 561308 393268 561372
rect 393332 561370 393338 561372
rect 406326 561370 406332 561372
rect 393332 561310 406332 561370
rect 393332 561308 393338 561310
rect 406326 561308 406332 561310
rect 406396 561308 406402 561372
rect 325693 560962 325759 560965
rect 335118 560962 335124 560964
rect 325693 560960 335124 560962
rect 325693 560904 325698 560960
rect 325754 560904 335124 560960
rect 325693 560902 335124 560904
rect 325693 560899 325759 560902
rect 335118 560900 335124 560902
rect 335188 560900 335194 560964
rect 376702 560900 376708 560964
rect 376772 560962 376778 560964
rect 386229 560962 386295 560965
rect 376772 560960 386295 560962
rect 376772 560904 386234 560960
rect 386290 560904 386295 560960
rect 376772 560902 386295 560904
rect 376772 560900 376778 560902
rect 386229 560899 386295 560902
rect 280102 560764 280108 560828
rect 280172 560826 280178 560828
rect 345013 560826 345079 560829
rect 357341 560828 357407 560829
rect 357341 560826 357388 560828
rect 280172 560766 293234 560826
rect 280172 560764 280178 560766
rect 280102 560554 280108 560556
rect 264286 560494 280108 560554
rect 253841 560418 253907 560421
rect 264286 560418 264346 560494
rect 280102 560492 280108 560494
rect 280172 560492 280178 560556
rect 293174 560554 293234 560766
rect 299430 560766 309058 560826
rect 299430 560554 299490 560766
rect 308998 560556 309058 560766
rect 345013 560824 357388 560826
rect 357452 560826 357458 560828
rect 367001 560826 367067 560829
rect 357452 560824 367067 560826
rect 345013 560768 345018 560824
rect 345074 560768 357346 560824
rect 357452 560768 367006 560824
rect 367062 560768 367067 560824
rect 345013 560766 357388 560768
rect 345013 560763 345079 560766
rect 357341 560764 357388 560766
rect 357452 560766 367067 560768
rect 357452 560764 357458 560766
rect 357341 560763 357407 560764
rect 367001 560763 367067 560766
rect 400213 560826 400279 560829
rect 400581 560826 400647 560829
rect 400213 560824 400647 560826
rect 400213 560768 400218 560824
rect 400274 560768 400586 560824
rect 400642 560768 400647 560824
rect 400213 560766 400647 560768
rect 400213 560763 400279 560766
rect 400581 560763 400647 560766
rect 424317 560826 424383 560829
rect 431861 560826 431927 560829
rect 424317 560824 431927 560826
rect 424317 560768 424322 560824
rect 424378 560768 431866 560824
rect 431922 560768 431927 560824
rect 424317 560766 431927 560768
rect 424317 560763 424383 560766
rect 431861 560763 431927 560766
rect 325693 560690 325759 560693
rect 318750 560688 325759 560690
rect 318750 560632 325698 560688
rect 325754 560632 325759 560688
rect 318750 560630 325759 560632
rect 293174 560494 299490 560554
rect 308990 560492 308996 560556
rect 309060 560492 309066 560556
rect 253841 560416 264346 560418
rect 253841 560360 253846 560416
rect 253902 560360 264346 560416
rect 253841 560358 264346 560360
rect 253841 560355 253907 560358
rect 308990 560356 308996 560420
rect 309060 560418 309066 560420
rect 318750 560418 318810 560630
rect 325693 560627 325759 560630
rect 335302 560628 335308 560692
rect 335372 560690 335378 560692
rect 344921 560690 344987 560693
rect 335372 560688 344987 560690
rect 335372 560632 344926 560688
rect 344982 560632 344987 560688
rect 335372 560630 344987 560632
rect 335372 560628 335378 560630
rect 344921 560627 344987 560630
rect 357341 560556 357407 560557
rect 357341 560552 357388 560556
rect 357452 560554 357458 560556
rect 367001 560554 367067 560557
rect 376702 560554 376708 560556
rect 357341 560496 357346 560552
rect 357341 560492 357388 560496
rect 357452 560494 357534 560554
rect 367001 560552 376708 560554
rect 367001 560496 367006 560552
rect 367062 560496 376708 560552
rect 367001 560494 376708 560496
rect 357452 560492 357458 560494
rect 357341 560491 357407 560492
rect 367001 560491 367067 560494
rect 376702 560492 376708 560494
rect 376772 560492 376778 560556
rect 386229 560554 386295 560557
rect 386413 560554 386479 560557
rect 386229 560552 386479 560554
rect 386229 560496 386234 560552
rect 386290 560496 386418 560552
rect 386474 560496 386479 560552
rect 386229 560494 386479 560496
rect 386229 560491 386295 560494
rect 386413 560491 386479 560494
rect 398925 560554 398991 560557
rect 405733 560554 405799 560557
rect 398925 560552 405799 560554
rect 398925 560496 398930 560552
rect 398986 560496 405738 560552
rect 405794 560496 405799 560552
rect 398925 560494 405799 560496
rect 398925 560491 398991 560494
rect 405733 560491 405799 560494
rect 431861 560554 431927 560557
rect 431861 560552 441722 560554
rect 431861 560496 431866 560552
rect 431922 560496 441722 560552
rect 431861 560494 441722 560496
rect 431861 560491 431927 560494
rect 309060 560358 318810 560418
rect 386505 560418 386571 560421
rect 395797 560418 395863 560421
rect 386505 560416 395863 560418
rect 386505 560360 386510 560416
rect 386566 560360 395802 560416
rect 395858 560360 395863 560416
rect 386505 560358 395863 560360
rect 309060 560356 309066 560358
rect 386505 560355 386571 560358
rect 395797 560355 395863 560358
rect 395981 560418 396047 560421
rect 398741 560418 398807 560421
rect 395981 560416 398807 560418
rect 395981 560360 395986 560416
rect 396042 560360 398746 560416
rect 398802 560360 398807 560416
rect 395981 560358 398807 560360
rect 395981 560355 396047 560358
rect 398741 560355 398807 560358
rect 400213 560418 400279 560421
rect 400581 560418 400647 560421
rect 400213 560416 400647 560418
rect 400213 560360 400218 560416
rect 400274 560360 400586 560416
rect 400642 560360 400647 560416
rect 400213 560358 400647 560360
rect 400213 560355 400279 560358
rect 400581 560355 400647 560358
rect 405825 560418 405891 560421
rect 411253 560418 411319 560421
rect 405825 560416 411319 560418
rect 405825 560360 405830 560416
rect 405886 560360 411258 560416
rect 411314 560360 411319 560416
rect 405825 560358 411319 560360
rect 405825 560355 405891 560358
rect 411253 560355 411319 560358
rect 400213 560282 400279 560285
rect 400581 560282 400647 560285
rect 400213 560280 400647 560282
rect 400213 560224 400218 560280
rect 400274 560224 400586 560280
rect 400642 560224 400647 560280
rect 400213 560222 400647 560224
rect 441662 560282 441722 560494
rect 447726 560282 447732 560284
rect 441662 560222 447732 560282
rect 400213 560219 400279 560222
rect 400581 560219 400647 560222
rect 447726 560220 447732 560222
rect 447796 560220 447802 560284
rect 372245 560146 372311 560149
rect 389081 560146 389147 560149
rect 372245 560144 389147 560146
rect 372245 560088 372250 560144
rect 372306 560088 389086 560144
rect 389142 560088 389147 560144
rect 372245 560086 389147 560088
rect 372245 560083 372311 560086
rect 389081 560083 389147 560086
rect 400213 560146 400279 560149
rect 400581 560146 400647 560149
rect 400213 560144 400647 560146
rect 400213 560088 400218 560144
rect 400274 560088 400586 560144
rect 400642 560088 400647 560144
rect 400213 560086 400647 560088
rect 400213 560083 400279 560086
rect 400581 560083 400647 560086
rect 385125 560010 385191 560013
rect 378734 560008 385191 560010
rect 378734 559952 385130 560008
rect 385186 559952 385191 560008
rect 378734 559950 385191 559952
rect 291561 559874 291627 559877
rect 296621 559874 296687 559877
rect 291561 559872 296687 559874
rect 291561 559816 291566 559872
rect 291622 559816 296626 559872
rect 296682 559816 296687 559872
rect 291561 559814 296687 559816
rect 291561 559811 291627 559814
rect 296621 559811 296687 559814
rect 299422 559812 299428 559876
rect 299492 559874 299498 559876
rect 304257 559874 304323 559877
rect 299492 559872 304323 559874
rect 299492 559816 304262 559872
rect 304318 559816 304323 559872
rect 299492 559814 304323 559816
rect 299492 559812 299498 559814
rect 304257 559811 304323 559814
rect 252645 559602 252711 559605
rect 277301 559602 277367 559605
rect 252645 559600 277367 559602
rect 252645 559544 252650 559600
rect 252706 559544 277306 559600
rect 277362 559544 277367 559600
rect 252645 559542 277367 559544
rect 252645 559539 252711 559542
rect 277301 559539 277367 559542
rect 296621 559602 296687 559605
rect 299422 559602 299428 559604
rect 296621 559600 299428 559602
rect 296621 559544 296626 559600
rect 296682 559544 299428 559600
rect 296621 559542 299428 559544
rect 296621 559539 296687 559542
rect 299422 559540 299428 559542
rect 299492 559540 299498 559604
rect 369853 559602 369919 559605
rect 378734 559602 378794 559950
rect 385125 559947 385191 559950
rect 400213 560010 400279 560013
rect 400581 560010 400647 560013
rect 400213 560008 400647 560010
rect 400213 559952 400218 560008
rect 400274 559952 400586 560008
rect 400642 559952 400647 560008
rect 400213 559950 400647 559952
rect 400213 559947 400279 559950
rect 400581 559947 400647 559950
rect 400305 559874 400371 559877
rect 400673 559874 400739 559877
rect 400305 559872 400739 559874
rect 400305 559816 400310 559872
rect 400366 559816 400678 559872
rect 400734 559816 400739 559872
rect 400305 559814 400739 559816
rect 400305 559811 400371 559814
rect 400673 559811 400739 559814
rect 409873 559874 409939 559877
rect 419349 559874 419415 559877
rect 409873 559872 419415 559874
rect 409873 559816 409878 559872
rect 409934 559816 419354 559872
rect 419410 559816 419415 559872
rect 409873 559814 419415 559816
rect 409873 559811 409939 559814
rect 419349 559811 419415 559814
rect 369853 559600 378794 559602
rect 369853 559544 369858 559600
rect 369914 559544 378794 559600
rect 369853 559542 378794 559544
rect 394049 559602 394115 559605
rect 405917 559602 405983 559605
rect 394049 559600 405983 559602
rect 394049 559544 394054 559600
rect 394110 559544 405922 559600
rect 405978 559544 405983 559600
rect 394049 559542 405983 559544
rect 369853 559539 369919 559542
rect 394049 559539 394115 559542
rect 405917 559539 405983 559542
rect 222142 559404 222148 559468
rect 222212 559466 222218 559468
rect 222212 559406 236562 559466
rect 222212 559404 222218 559406
rect 231025 559330 231091 559333
rect 231710 559330 231716 559332
rect 231025 559328 231716 559330
rect 231025 559272 231030 559328
rect 231086 559272 231716 559328
rect 231025 559270 231716 559272
rect 231025 559267 231091 559270
rect 231710 559268 231716 559270
rect 231780 559268 231786 559332
rect 232865 559330 232931 559333
rect 232998 559330 233004 559332
rect 232865 559328 233004 559330
rect 232865 559272 232870 559328
rect 232926 559272 233004 559328
rect 232865 559270 233004 559272
rect 232865 559267 232931 559270
rect 232998 559268 233004 559270
rect 233068 559268 233074 559332
rect 234286 559268 234292 559332
rect 234356 559330 234362 559332
rect 234613 559330 234679 559333
rect 234356 559328 234679 559330
rect 234356 559272 234618 559328
rect 234674 559272 234679 559328
rect 234356 559270 234679 559272
rect 234356 559268 234362 559270
rect 234613 559267 234679 559270
rect 222142 559194 222148 559196
rect 215342 559134 222148 559194
rect 3417 559058 3483 559061
rect 215342 559058 215402 559134
rect 222142 559132 222148 559134
rect 222212 559132 222218 559196
rect 3417 559056 215402 559058
rect 3417 559000 3422 559056
rect 3478 559000 215402 559056
rect 3417 558998 215402 559000
rect 236502 559058 236562 559406
rect 236678 559404 236684 559468
rect 236748 559466 236754 559468
rect 240133 559466 240199 559469
rect 304257 559466 304323 559469
rect 307702 559466 307708 559468
rect 236748 559464 240199 559466
rect 236748 559408 240138 559464
rect 240194 559408 240199 559464
rect 236748 559406 240199 559408
rect 236748 559404 236754 559406
rect 240133 559403 240199 559406
rect 252694 559406 291762 559466
rect 236729 559330 236795 559333
rect 238201 559332 238267 559333
rect 237230 559330 237236 559332
rect 236729 559328 237236 559330
rect 236729 559272 236734 559328
rect 236790 559272 237236 559328
rect 236729 559270 237236 559272
rect 236729 559267 236795 559270
rect 237230 559268 237236 559270
rect 237300 559268 237306 559332
rect 238150 559330 238156 559332
rect 238110 559270 238156 559330
rect 238220 559328 238267 559332
rect 238262 559272 238267 559328
rect 238150 559268 238156 559270
rect 238220 559268 238267 559272
rect 238201 559267 238267 559268
rect 248781 559330 248847 559333
rect 252553 559330 252619 559333
rect 248781 559328 252619 559330
rect 248781 559272 248786 559328
rect 248842 559272 252558 559328
rect 252614 559272 252619 559328
rect 248781 559270 252619 559272
rect 248781 559267 248847 559270
rect 252553 559267 252619 559270
rect 252502 559132 252508 559196
rect 252572 559194 252578 559196
rect 252694 559194 252754 559406
rect 277301 559330 277367 559333
rect 291561 559330 291627 559333
rect 277301 559328 291627 559330
rect 277301 559272 277306 559328
rect 277362 559272 291566 559328
rect 291622 559272 291627 559328
rect 277301 559270 291627 559272
rect 291702 559330 291762 559406
rect 304257 559464 307708 559466
rect 304257 559408 304262 559464
rect 304318 559408 307708 559464
rect 304257 559406 307708 559408
rect 304257 559403 304323 559406
rect 307702 559404 307708 559406
rect 307772 559404 307778 559468
rect 321694 559406 336106 559466
rect 299422 559330 299428 559332
rect 291702 559270 299428 559330
rect 277301 559267 277367 559270
rect 291561 559267 291627 559270
rect 299422 559268 299428 559270
rect 299492 559268 299498 559332
rect 307886 559268 307892 559332
rect 307956 559330 307962 559332
rect 321694 559330 321754 559406
rect 307956 559270 321754 559330
rect 336046 559330 336106 559406
rect 370086 559406 383394 559466
rect 361297 559330 361363 559333
rect 336046 559328 361363 559330
rect 336046 559272 361302 559328
rect 361358 559272 361363 559328
rect 336046 559270 361363 559272
rect 307956 559268 307962 559270
rect 361297 559267 361363 559270
rect 361481 559330 361547 559333
rect 370086 559330 370146 559406
rect 383193 559332 383259 559333
rect 383142 559330 383148 559332
rect 361481 559328 370146 559330
rect 361481 559272 361486 559328
rect 361542 559272 370146 559328
rect 361481 559270 370146 559272
rect 383102 559270 383148 559330
rect 383212 559328 383259 559332
rect 383254 559272 383259 559328
rect 361481 559267 361547 559270
rect 383142 559268 383148 559270
rect 383212 559268 383259 559272
rect 383334 559330 383394 559406
rect 384062 559404 384068 559468
rect 384132 559466 384138 559468
rect 384132 559406 394434 559466
rect 384132 559404 384138 559406
rect 394049 559330 394115 559333
rect 383334 559270 384314 559330
rect 383193 559267 383259 559268
rect 252572 559134 252754 559194
rect 252572 559132 252578 559134
rect 311934 559132 311940 559196
rect 312004 559194 312010 559196
rect 312004 559134 318810 559194
rect 312004 559132 312010 559134
rect 318750 559060 318810 559134
rect 331262 559134 336842 559194
rect 244038 559058 244044 559060
rect 236502 558998 244044 559058
rect 3417 558995 3483 558998
rect 244038 558996 244044 558998
rect 244108 558996 244114 559060
rect 299422 558996 299428 559060
rect 299492 559058 299498 559060
rect 311750 559058 311756 559060
rect 299492 558998 311756 559058
rect 299492 558996 299498 558998
rect 311750 558996 311756 558998
rect 311820 558996 311826 559060
rect 318742 558996 318748 559060
rect 318812 558996 318818 559060
rect 244038 558724 244044 558788
rect 244108 558786 244114 558788
rect 252502 558786 252508 558788
rect 244108 558726 252508 558786
rect 244108 558724 244114 558726
rect 252502 558724 252508 558726
rect 252572 558724 252578 558788
rect 318742 558724 318748 558788
rect 318812 558786 318818 558788
rect 331262 558786 331322 559134
rect 336782 559058 336842 559134
rect 352046 559132 352052 559196
rect 352116 559194 352122 559196
rect 384062 559194 384068 559196
rect 352116 559134 361498 559194
rect 352116 559132 352122 559134
rect 338062 559058 338068 559060
rect 336782 558998 338068 559058
rect 338062 558996 338068 558998
rect 338132 558996 338138 559060
rect 351862 559058 351868 559060
rect 351686 558998 351868 559058
rect 318812 558726 331322 558786
rect 318812 558724 318818 558726
rect 338062 558724 338068 558788
rect 338132 558786 338138 558788
rect 351686 558786 351746 558998
rect 351862 558996 351868 558998
rect 351932 558996 351938 559060
rect 361438 559058 361498 559134
rect 375974 559134 384068 559194
rect 375974 559058 376034 559134
rect 384062 559132 384068 559134
rect 384132 559132 384138 559196
rect 384254 559194 384314 559270
rect 394006 559328 394115 559330
rect 394006 559272 394054 559328
rect 394110 559272 394115 559328
rect 394006 559267 394115 559272
rect 394006 559194 394066 559267
rect 384254 559134 394066 559194
rect 361438 558998 376034 559058
rect 394374 559058 394434 559406
rect 409086 559404 409092 559468
rect 409156 559466 409162 559468
rect 434621 559466 434687 559469
rect 442809 559466 442875 559469
rect 409156 559406 415364 559466
rect 409156 559404 409162 559406
rect 396022 559268 396028 559332
rect 396092 559330 396098 559332
rect 396092 559270 404370 559330
rect 396092 559268 396098 559270
rect 396022 559058 396028 559060
rect 394374 558998 396028 559058
rect 396022 558996 396028 558998
rect 396092 558996 396098 559060
rect 404310 559058 404370 559270
rect 415304 559194 415364 559406
rect 434621 559464 442875 559466
rect 434621 559408 434626 559464
rect 434682 559408 442814 559464
rect 442870 559408 442875 559464
rect 434621 559406 442875 559408
rect 434621 559403 434687 559406
rect 442809 559403 442875 559406
rect 427678 559330 428106 559364
rect 434621 559330 434687 559333
rect 427678 559328 434687 559330
rect 427678 559304 434626 559328
rect 427678 559194 427738 559304
rect 428046 559272 434626 559304
rect 434682 559272 434687 559328
rect 428046 559270 434687 559272
rect 434621 559267 434687 559270
rect 444414 559268 444420 559332
rect 444484 559330 444490 559332
rect 444557 559330 444623 559333
rect 444484 559328 444623 559330
rect 444484 559272 444562 559328
rect 444618 559272 444623 559328
rect 444484 559270 444623 559272
rect 444484 559268 444490 559270
rect 444557 559267 444623 559270
rect 445702 559268 445708 559332
rect 445772 559330 445778 559332
rect 446581 559330 446647 559333
rect 448513 559332 448579 559333
rect 448462 559330 448468 559332
rect 445772 559328 446647 559330
rect 445772 559272 446586 559328
rect 446642 559272 446647 559328
rect 445772 559270 446647 559272
rect 448422 559270 448468 559330
rect 448532 559328 448579 559332
rect 448574 559272 448579 559328
rect 445772 559268 445778 559270
rect 446581 559267 446647 559270
rect 448462 559268 448468 559270
rect 448532 559268 448579 559272
rect 448513 559267 448579 559268
rect 415304 559134 427738 559194
rect 409086 559058 409092 559060
rect 404310 558998 409092 559058
rect 409086 558996 409092 558998
rect 409156 558996 409162 559060
rect 338132 558726 351746 558786
rect 338132 558724 338138 558726
rect 2957 558242 3023 558245
rect 383142 558242 383148 558244
rect 2957 558240 383148 558242
rect 2957 558184 2962 558240
rect 3018 558184 383148 558240
rect 2957 558182 383148 558184
rect 2957 558179 3023 558182
rect 383142 558180 383148 558182
rect 383212 558180 383218 558244
rect 579705 557290 579771 557293
rect 583520 557290 584960 557380
rect 579705 557288 584960 557290
rect 579705 557232 579710 557288
rect 579766 557232 584960 557288
rect 579705 557230 584960 557232
rect 579705 557227 579771 557230
rect 583520 557140 584960 557230
rect -960 553074 480 553164
rect 2773 553074 2839 553077
rect -960 553072 2839 553074
rect -960 553016 2778 553072
rect 2834 553016 2839 553072
rect -960 553014 2839 553016
rect -960 552924 480 553014
rect 2773 553011 2839 553014
rect 579797 545594 579863 545597
rect 583520 545594 584960 545684
rect 579797 545592 584960 545594
rect 579797 545536 579802 545592
rect 579858 545536 584960 545592
rect 579797 545534 584960 545536
rect 579797 545531 579863 545534
rect 583520 545444 584960 545534
rect -960 538658 480 538748
rect 2957 538658 3023 538661
rect -960 538656 3023 538658
rect -960 538600 2962 538656
rect 3018 538600 3023 538656
rect -960 538598 3023 538600
rect -960 538508 480 538598
rect 2957 538595 3023 538598
rect 579797 533898 579863 533901
rect 583520 533898 584960 533988
rect 579797 533896 584960 533898
rect 579797 533840 579802 533896
rect 579858 533840 584960 533896
rect 579797 533838 584960 533840
rect 579797 533835 579863 533838
rect 583520 533748 584960 533838
rect -960 524092 480 524332
rect 583520 521916 584960 522156
rect 579797 510370 579863 510373
rect 583520 510370 584960 510460
rect 579797 510368 584960 510370
rect 579797 510312 579802 510368
rect 579858 510312 584960 510368
rect 579797 510310 584960 510312
rect 579797 510307 579863 510310
rect 583520 510220 584960 510310
rect -960 509962 480 510052
rect 3049 509962 3115 509965
rect -960 509960 3115 509962
rect -960 509904 3054 509960
rect 3110 509904 3115 509960
rect -960 509902 3115 509904
rect -960 509812 480 509902
rect 3049 509899 3115 509902
rect 579797 498674 579863 498677
rect 583520 498674 584960 498764
rect 579797 498672 584960 498674
rect 579797 498616 579802 498672
rect 579858 498616 584960 498672
rect 579797 498614 584960 498616
rect 579797 498611 579863 498614
rect 583520 498524 584960 498614
rect -960 495546 480 495636
rect 3049 495546 3115 495549
rect -960 495544 3115 495546
rect -960 495488 3054 495544
rect 3110 495488 3115 495544
rect -960 495486 3115 495488
rect -960 495396 480 495486
rect 3049 495483 3115 495486
rect 583520 486842 584960 486932
rect 583342 486782 584960 486842
rect 446254 486100 446260 486164
rect 446324 486162 446330 486164
rect 446324 486102 451290 486162
rect 446324 486100 446330 486102
rect 451230 486026 451290 486102
rect 460982 486102 470610 486162
rect 451230 485966 460858 486026
rect 460798 485890 460858 485966
rect 460982 485890 461042 486102
rect 470550 486026 470610 486102
rect 480302 486102 489930 486162
rect 470550 485966 480178 486026
rect 460798 485830 461042 485890
rect 480118 485890 480178 485966
rect 480302 485890 480362 486102
rect 489870 486026 489930 486102
rect 499622 486102 509250 486162
rect 489870 485966 499498 486026
rect 480118 485830 480362 485890
rect 499438 485890 499498 485966
rect 499622 485890 499682 486102
rect 509190 486026 509250 486102
rect 518942 486102 528570 486162
rect 509190 485966 518818 486026
rect 499438 485830 499682 485890
rect 518758 485890 518818 485966
rect 518942 485890 519002 486102
rect 528510 486026 528570 486102
rect 538262 486102 547890 486162
rect 528510 485966 538138 486026
rect 518758 485830 519002 485890
rect 538078 485890 538138 485966
rect 538262 485890 538322 486102
rect 547830 486026 547890 486102
rect 557582 486102 567210 486162
rect 547830 485966 557458 486026
rect 538078 485830 538322 485890
rect 557398 485890 557458 485966
rect 557582 485890 557642 486102
rect 567150 486026 567210 486102
rect 583342 486026 583402 486782
rect 583520 486692 584960 486782
rect 567150 485966 576778 486026
rect 557398 485830 557642 485890
rect 576718 485890 576778 485966
rect 576902 485966 583402 486026
rect 576902 485890 576962 485966
rect 576718 485830 576962 485890
rect -960 481130 480 481220
rect 3049 481130 3115 481133
rect -960 481128 3115 481130
rect -960 481072 3054 481128
rect 3110 481072 3115 481128
rect -960 481070 3115 481072
rect -960 480980 480 481070
rect 3049 481067 3115 481070
rect 583520 474996 584960 475236
rect -960 466700 480 466940
rect 579797 463450 579863 463453
rect 583520 463450 584960 463540
rect 579797 463448 584960 463450
rect 579797 463392 579802 463448
rect 579858 463392 584960 463448
rect 579797 463390 584960 463392
rect 579797 463387 579863 463390
rect 583520 463300 584960 463390
rect -960 452434 480 452524
rect 3141 452434 3207 452437
rect -960 452432 3207 452434
rect -960 452376 3146 452432
rect 3202 452376 3207 452432
rect -960 452374 3207 452376
rect -960 452284 480 452374
rect 3141 452371 3207 452374
rect 579797 451754 579863 451757
rect 583520 451754 584960 451844
rect 579797 451752 584960 451754
rect 579797 451696 579802 451752
rect 579858 451696 584960 451752
rect 579797 451694 584960 451696
rect 579797 451691 579863 451694
rect 583520 451604 584960 451694
rect 579797 439922 579863 439925
rect 583520 439922 584960 440012
rect 579797 439920 584960 439922
rect 579797 439864 579802 439920
rect 579858 439864 584960 439920
rect 579797 439862 584960 439864
rect 579797 439859 579863 439862
rect 583520 439772 584960 439862
rect -960 438018 480 438108
rect 3141 438018 3207 438021
rect -960 438016 3207 438018
rect -960 437960 3146 438016
rect 3202 437960 3207 438016
rect -960 437958 3207 437960
rect -960 437868 480 437958
rect 3141 437955 3207 437958
rect 583520 428076 584960 428316
rect -960 423738 480 423828
rect 2773 423738 2839 423741
rect -960 423736 2839 423738
rect -960 423680 2778 423736
rect 2834 423680 2839 423736
rect -960 423678 2839 423680
rect -960 423588 480 423678
rect 2773 423675 2839 423678
rect 579797 416530 579863 416533
rect 583520 416530 584960 416620
rect 579797 416528 584960 416530
rect 579797 416472 579802 416528
rect 579858 416472 584960 416528
rect 579797 416470 584960 416472
rect 579797 416467 579863 416470
rect 583520 416380 584960 416470
rect -960 409172 480 409412
rect 579797 404834 579863 404837
rect 583520 404834 584960 404924
rect 579797 404832 584960 404834
rect 579797 404776 579802 404832
rect 579858 404776 584960 404832
rect 579797 404774 584960 404776
rect 579797 404771 579863 404774
rect 583520 404684 584960 404774
rect -960 395042 480 395132
rect 3233 395042 3299 395045
rect -960 395040 3299 395042
rect -960 394984 3238 395040
rect 3294 394984 3299 395040
rect -960 394982 3299 394984
rect -960 394892 480 394982
rect 3233 394979 3299 394982
rect 579797 393002 579863 393005
rect 583520 393002 584960 393092
rect 579797 393000 584960 393002
rect 579797 392944 579802 393000
rect 579858 392944 584960 393000
rect 579797 392942 584960 392944
rect 579797 392939 579863 392942
rect 583520 392852 584960 392942
rect 583520 381156 584960 381396
rect -960 380626 480 380716
rect 3141 380626 3207 380629
rect -960 380624 3207 380626
rect -960 380568 3146 380624
rect 3202 380568 3207 380624
rect -960 380566 3207 380568
rect -960 380476 480 380566
rect 3141 380563 3207 380566
rect 579797 369610 579863 369613
rect 583520 369610 584960 369700
rect 579797 369608 584960 369610
rect 579797 369552 579802 369608
rect 579858 369552 584960 369608
rect 579797 369550 584960 369552
rect 579797 369547 579863 369550
rect 583520 369460 584960 369550
rect -960 366210 480 366300
rect 2773 366210 2839 366213
rect -960 366208 2839 366210
rect -960 366152 2778 366208
rect 2834 366152 2839 366208
rect -960 366150 2839 366152
rect -960 366060 480 366150
rect 2773 366147 2839 366150
rect 579889 357914 579955 357917
rect 583520 357914 584960 358004
rect 579889 357912 584960 357914
rect 579889 357856 579894 357912
rect 579950 357856 584960 357912
rect 579889 357854 584960 357856
rect 579889 357851 579955 357854
rect 583520 357764 584960 357854
rect -960 351780 480 352020
rect 579889 346082 579955 346085
rect 583520 346082 584960 346172
rect 579889 346080 584960 346082
rect 579889 346024 579894 346080
rect 579950 346024 584960 346080
rect 579889 346022 584960 346024
rect 579889 346019 579955 346022
rect 583520 345932 584960 346022
rect 325141 338330 325207 338333
rect 324454 338328 325207 338330
rect 324454 338272 325146 338328
rect 325202 338272 325207 338328
rect 324454 338270 325207 338272
rect 324454 338194 324514 338270
rect 325141 338267 325207 338270
rect 324589 338194 324655 338197
rect 324454 338192 324655 338194
rect 324454 338136 324594 338192
rect 324650 338136 324655 338192
rect 324454 338134 324655 338136
rect 324589 338131 324655 338134
rect 236862 338058 236868 338060
rect 614 337998 236868 338058
rect -960 337514 480 337604
rect 614 337514 674 337998
rect 236862 337996 236868 337998
rect 236932 337996 236938 338060
rect 434989 337922 435055 337925
rect 438209 337922 438275 337925
rect 434989 337920 438275 337922
rect 434989 337864 434994 337920
rect 435050 337864 438214 337920
rect 438270 337864 438275 337920
rect 434989 337862 438275 337864
rect 434989 337859 435055 337862
rect 438209 337859 438275 337862
rect 448145 337786 448211 337789
rect 449157 337786 449223 337789
rect 448145 337784 449223 337786
rect 448145 337728 448150 337784
rect 448206 337728 449162 337784
rect 449218 337728 449223 337784
rect 448145 337726 449223 337728
rect 448145 337723 448211 337726
rect 449157 337723 449223 337726
rect -960 337454 674 337514
rect -960 337364 480 337454
rect 10317 337378 10383 337381
rect 231761 337378 231827 337381
rect 10317 337376 231827 337378
rect 10317 337320 10322 337376
rect 10378 337320 231766 337376
rect 231822 337320 231827 337376
rect 10317 337318 231827 337320
rect 10317 337315 10383 337318
rect 231761 337315 231827 337318
rect 273897 337378 273963 337381
rect 332317 337378 332383 337381
rect 273897 337376 332383 337378
rect 273897 337320 273902 337376
rect 273958 337320 332322 337376
rect 332378 337320 332383 337376
rect 273897 337318 332383 337320
rect 273897 337315 273963 337318
rect 332317 337315 332383 337318
rect 449525 337378 449591 337381
rect 530577 337378 530643 337381
rect 449525 337376 530643 337378
rect 449525 337320 449530 337376
rect 449586 337320 530582 337376
rect 530638 337320 530643 337376
rect 449525 337318 530643 337320
rect 449525 337315 449591 337318
rect 530577 337315 530643 337318
rect 138013 337242 138079 337245
rect 147581 337242 147647 337245
rect 138013 337240 147647 337242
rect 138013 337184 138018 337240
rect 138074 337184 147586 337240
rect 147642 337184 147647 337240
rect 138013 337182 147647 337184
rect 138013 337179 138079 337182
rect 147581 337179 147647 337182
rect 157333 337242 157399 337245
rect 166901 337242 166967 337245
rect 157333 337240 166967 337242
rect 157333 337184 157338 337240
rect 157394 337184 166906 337240
rect 166962 337184 166967 337240
rect 157333 337182 166967 337184
rect 157333 337179 157399 337182
rect 166901 337179 166967 337182
rect 176653 337242 176719 337245
rect 186221 337242 186287 337245
rect 176653 337240 186287 337242
rect 176653 337184 176658 337240
rect 176714 337184 186226 337240
rect 186282 337184 186287 337240
rect 176653 337182 186287 337184
rect 176653 337179 176719 337182
rect 186221 337179 186287 337182
rect 195973 337242 196039 337245
rect 205541 337242 205607 337245
rect 195973 337240 205607 337242
rect 195973 337184 195978 337240
rect 196034 337184 205546 337240
rect 205602 337184 205607 337240
rect 195973 337182 205607 337184
rect 195973 337179 196039 337182
rect 205541 337179 205607 337182
rect 215293 337242 215359 337245
rect 224861 337242 224927 337245
rect 215293 337240 224927 337242
rect 215293 337184 215298 337240
rect 215354 337184 224866 337240
rect 224922 337184 224927 337240
rect 215293 337182 224927 337184
rect 215293 337179 215359 337182
rect 224861 337179 224927 337182
rect 250161 335338 250227 335341
rect 250118 335336 250227 335338
rect 250118 335280 250166 335336
rect 250222 335280 250227 335336
rect 250118 335275 250227 335280
rect 250118 335202 250178 335275
rect 250253 335202 250319 335205
rect 250118 335200 250319 335202
rect 250118 335144 250258 335200
rect 250314 335144 250319 335200
rect 250118 335142 250319 335144
rect 250253 335139 250319 335142
rect 583520 334236 584960 334476
rect 310145 328538 310211 328541
rect 314009 328538 314075 328541
rect 309366 328536 310211 328538
rect 309366 328480 310150 328536
rect 310206 328480 310211 328536
rect 309366 328478 310211 328480
rect 309366 328405 309426 328478
rect 310145 328475 310211 328478
rect 313598 328536 314075 328538
rect 313598 328480 314014 328536
rect 314070 328480 314075 328536
rect 313598 328478 314075 328480
rect 309366 328400 309475 328405
rect 309366 328344 309414 328400
rect 309470 328344 309475 328400
rect 309366 328342 309475 328344
rect 313598 328402 313658 328478
rect 314009 328475 314075 328478
rect 313733 328402 313799 328405
rect 313598 328400 313799 328402
rect 313598 328344 313738 328400
rect 313794 328344 313799 328400
rect 313598 328342 313799 328344
rect 309409 328339 309475 328342
rect 313733 328339 313799 328342
rect 249977 325682 250043 325685
rect 250253 325682 250319 325685
rect 249977 325680 250319 325682
rect 249977 325624 249982 325680
rect 250038 325624 250258 325680
rect 250314 325624 250319 325680
rect 249977 325622 250319 325624
rect 249977 325619 250043 325622
rect 250253 325619 250319 325622
rect -960 323098 480 323188
rect 3325 323098 3391 323101
rect -960 323096 3391 323098
rect -960 323040 3330 323096
rect 3386 323040 3391 323096
rect -960 323038 3391 323040
rect -960 322948 480 323038
rect 3325 323035 3391 323038
rect 579889 322690 579955 322693
rect 583520 322690 584960 322780
rect 579889 322688 584960 322690
rect 579889 322632 579894 322688
rect 579950 322632 584960 322688
rect 579889 322630 584960 322632
rect 579889 322627 579955 322630
rect 583520 322540 584960 322630
rect 310789 316026 310855 316029
rect 310654 316024 310855 316026
rect 310654 315968 310794 316024
rect 310850 315968 310855 316024
rect 310654 315966 310855 315968
rect 310654 315890 310714 315966
rect 310789 315963 310855 315966
rect 313457 316026 313523 316029
rect 313641 316026 313707 316029
rect 313457 316024 313707 316026
rect 313457 315968 313462 316024
rect 313518 315968 313646 316024
rect 313702 315968 313707 316024
rect 313457 315966 313707 315968
rect 313457 315963 313523 315966
rect 313641 315963 313707 315966
rect 310881 315890 310947 315893
rect 310654 315888 310947 315890
rect 310654 315832 310886 315888
rect 310942 315832 310947 315888
rect 310654 315830 310947 315832
rect 310881 315827 310947 315830
rect 579981 310858 580047 310861
rect 583520 310858 584960 310948
rect 579981 310856 584960 310858
rect 579981 310800 579986 310856
rect 580042 310800 584960 310856
rect 579981 310798 584960 310800
rect 579981 310795 580047 310798
rect 583520 310708 584960 310798
rect 236678 309090 236684 309092
rect 614 309030 236684 309090
rect -960 308818 480 308908
rect 614 308818 674 309030
rect 236678 309028 236684 309030
rect 236748 309028 236754 309092
rect -960 308758 674 308818
rect -960 308668 480 308758
rect 253933 306370 253999 306373
rect 254117 306370 254183 306373
rect 253933 306368 254183 306370
rect 253933 306312 253938 306368
rect 253994 306312 254122 306368
rect 254178 306312 254183 306368
rect 253933 306310 254183 306312
rect 253933 306307 253999 306310
rect 254117 306307 254183 306310
rect 288801 299434 288867 299437
rect 288985 299434 289051 299437
rect 288801 299432 289051 299434
rect 288801 299376 288806 299432
rect 288862 299376 288990 299432
rect 289046 299376 289051 299432
rect 288801 299374 289051 299376
rect 288801 299371 288867 299374
rect 288985 299371 289051 299374
rect 434345 299434 434411 299437
rect 434478 299434 434484 299436
rect 434345 299432 434484 299434
rect 434345 299376 434350 299432
rect 434406 299376 434484 299432
rect 434345 299374 434484 299376
rect 434345 299371 434411 299374
rect 434478 299372 434484 299374
rect 434548 299372 434554 299436
rect 579889 299162 579955 299165
rect 583520 299162 584960 299252
rect 579889 299160 584960 299162
rect 579889 299104 579894 299160
rect 579950 299104 584960 299160
rect 579889 299102 584960 299104
rect 579889 299099 579955 299102
rect 583520 299012 584960 299102
rect 229369 298074 229435 298077
rect 229553 298074 229619 298077
rect 229369 298072 229619 298074
rect 229369 298016 229374 298072
rect 229430 298016 229558 298072
rect 229614 298016 229619 298072
rect 229369 298014 229619 298016
rect 229369 298011 229435 298014
rect 229553 298011 229619 298014
rect 239029 296714 239095 296717
rect 239305 296714 239371 296717
rect 239029 296712 239371 296714
rect 239029 296656 239034 296712
rect 239090 296656 239310 296712
rect 239366 296656 239371 296712
rect 239029 296654 239371 296656
rect 239029 296651 239095 296654
rect 239305 296651 239371 296654
rect -960 294402 480 294492
rect 2773 294402 2839 294405
rect -960 294400 2839 294402
rect -960 294344 2778 294400
rect 2834 294344 2839 294400
rect -960 294342 2839 294344
rect -960 294252 480 294342
rect 2773 294339 2839 294342
rect 434345 289914 434411 289917
rect 434478 289914 434484 289916
rect 434345 289912 434484 289914
rect 434345 289856 434350 289912
rect 434406 289856 434484 289912
rect 434345 289854 434484 289856
rect 434345 289851 434411 289854
rect 434478 289852 434484 289854
rect 434548 289852 434554 289916
rect 251173 288418 251239 288421
rect 251357 288418 251423 288421
rect 251173 288416 251423 288418
rect 251173 288360 251178 288416
rect 251234 288360 251362 288416
rect 251418 288360 251423 288416
rect 251173 288358 251423 288360
rect 251173 288355 251239 288358
rect 251357 288355 251423 288358
rect 583520 287316 584960 287556
rect 347773 280258 347839 280261
rect 347957 280258 348023 280261
rect 347773 280256 348023 280258
rect -960 280122 480 280212
rect 347773 280200 347778 280256
rect 347834 280200 347962 280256
rect 348018 280200 348023 280256
rect 347773 280198 348023 280200
rect 347773 280195 347839 280198
rect 347957 280195 348023 280198
rect 3141 280122 3207 280125
rect -960 280120 3207 280122
rect -960 280064 3146 280120
rect 3202 280064 3207 280120
rect -960 280062 3207 280064
rect -960 279972 480 280062
rect 3141 280059 3207 280062
rect 434345 280122 434411 280125
rect 434478 280122 434484 280124
rect 434345 280120 434484 280122
rect 434345 280064 434350 280120
rect 434406 280064 434484 280120
rect 434345 280062 434484 280064
rect 434345 280059 434411 280062
rect 434478 280060 434484 280062
rect 434548 280060 434554 280124
rect 240225 278762 240291 278765
rect 240409 278762 240475 278765
rect 240225 278760 240475 278762
rect 240225 278704 240230 278760
rect 240286 278704 240414 278760
rect 240470 278704 240475 278760
rect 240225 278702 240475 278704
rect 240225 278699 240291 278702
rect 240409 278699 240475 278702
rect 241881 278762 241947 278765
rect 242065 278762 242131 278765
rect 241881 278760 242131 278762
rect 241881 278704 241886 278760
rect 241942 278704 242070 278760
rect 242126 278704 242131 278760
rect 241881 278702 242131 278704
rect 241881 278699 241947 278702
rect 242065 278699 242131 278702
rect 291469 278762 291535 278765
rect 291653 278762 291719 278765
rect 291469 278760 291719 278762
rect 291469 278704 291474 278760
rect 291530 278704 291658 278760
rect 291714 278704 291719 278760
rect 291469 278702 291719 278704
rect 291469 278699 291535 278702
rect 291653 278699 291719 278702
rect 305269 278762 305335 278765
rect 305545 278762 305611 278765
rect 305269 278760 305611 278762
rect 305269 278704 305274 278760
rect 305330 278704 305550 278760
rect 305606 278704 305611 278760
rect 305269 278702 305611 278704
rect 305269 278699 305335 278702
rect 305545 278699 305611 278702
rect 327349 278762 327415 278765
rect 327625 278762 327691 278765
rect 327349 278760 327691 278762
rect 327349 278704 327354 278760
rect 327410 278704 327630 278760
rect 327686 278704 327691 278760
rect 327349 278702 327691 278704
rect 327349 278699 327415 278702
rect 327625 278699 327691 278702
rect 234613 277402 234679 277405
rect 234797 277402 234863 277405
rect 234613 277400 234863 277402
rect 234613 277344 234618 277400
rect 234674 277344 234802 277400
rect 234858 277344 234863 277400
rect 234613 277342 234863 277344
rect 234613 277339 234679 277342
rect 234797 277339 234863 277342
rect 580073 275770 580139 275773
rect 583520 275770 584960 275860
rect 580073 275768 584960 275770
rect 580073 275712 580078 275768
rect 580134 275712 584960 275768
rect 580073 275710 584960 275712
rect 580073 275707 580139 275710
rect 583520 275620 584960 275710
rect 267273 270738 267339 270741
rect 266862 270736 267339 270738
rect 266862 270680 267278 270736
rect 267334 270680 267339 270736
rect 266862 270678 267339 270680
rect 266862 270602 266922 270678
rect 267273 270675 267339 270678
rect 266997 270602 267063 270605
rect 266862 270600 267063 270602
rect 266862 270544 267002 270600
rect 267058 270544 267063 270600
rect 266862 270542 267063 270544
rect 266997 270539 267063 270542
rect 434345 270602 434411 270605
rect 434478 270602 434484 270604
rect 434345 270600 434484 270602
rect 434345 270544 434350 270600
rect 434406 270544 434484 270600
rect 434345 270542 434484 270544
rect 434345 270539 434411 270542
rect 434478 270540 434484 270542
rect 434548 270540 434554 270604
rect 266997 269106 267063 269109
rect 267181 269106 267247 269109
rect 266997 269104 267247 269106
rect 266997 269048 267002 269104
rect 267058 269048 267186 269104
rect 267242 269048 267247 269104
rect 266997 269046 267247 269048
rect 266997 269043 267063 269046
rect 267181 269043 267247 269046
rect -960 265706 480 265796
rect 4061 265706 4127 265709
rect -960 265704 4127 265706
rect -960 265648 4066 265704
rect 4122 265648 4127 265704
rect -960 265646 4127 265648
rect -960 265556 480 265646
rect 4061 265643 4127 265646
rect 580165 263938 580231 263941
rect 583520 263938 584960 264028
rect 580165 263936 584960 263938
rect 580165 263880 580170 263936
rect 580226 263880 584960 263936
rect 580165 263878 584960 263880
rect 580165 263875 580231 263878
rect 583520 263788 584960 263878
rect 434345 260810 434411 260813
rect 434478 260810 434484 260812
rect 434345 260808 434484 260810
rect 434345 260752 434350 260808
rect 434406 260752 434484 260808
rect 434345 260750 434484 260752
rect 434345 260747 434411 260750
rect 434478 260748 434484 260750
rect 434548 260748 434554 260812
rect 240225 259450 240291 259453
rect 240409 259450 240475 259453
rect 240225 259448 240475 259450
rect 240225 259392 240230 259448
rect 240286 259392 240414 259448
rect 240470 259392 240475 259448
rect 240225 259390 240475 259392
rect 240225 259387 240291 259390
rect 240409 259387 240475 259390
rect 241881 259450 241947 259453
rect 242065 259450 242131 259453
rect 241881 259448 242131 259450
rect 241881 259392 241886 259448
rect 241942 259392 242070 259448
rect 242126 259392 242131 259448
rect 241881 259390 242131 259392
rect 241881 259387 241947 259390
rect 242065 259387 242131 259390
rect 3141 252514 3207 252517
rect 236494 252514 236500 252516
rect 3141 252512 236500 252514
rect 3141 252456 3146 252512
rect 3202 252456 236500 252512
rect 3141 252454 236500 252456
rect 3141 252451 3207 252454
rect 236494 252452 236500 252454
rect 236564 252452 236570 252516
rect 580901 252242 580967 252245
rect 583520 252242 584960 252332
rect 580901 252240 584960 252242
rect 580901 252184 580906 252240
rect 580962 252184 584960 252240
rect 580901 252182 584960 252184
rect 580901 252179 580967 252182
rect 583520 252092 584960 252182
rect 345289 251426 345355 251429
rect 345062 251424 345355 251426
rect -960 251290 480 251380
rect 345062 251368 345294 251424
rect 345350 251368 345355 251424
rect 345062 251366 345355 251368
rect 3141 251290 3207 251293
rect -960 251288 3207 251290
rect -960 251232 3146 251288
rect 3202 251232 3207 251288
rect -960 251230 3207 251232
rect 345062 251290 345122 251366
rect 345289 251363 345355 251366
rect 345197 251290 345263 251293
rect 345062 251288 345263 251290
rect 345062 251232 345202 251288
rect 345258 251232 345263 251288
rect 345062 251230 345263 251232
rect -960 251140 480 251230
rect 3141 251227 3207 251230
rect 345197 251227 345263 251230
rect 434345 251290 434411 251293
rect 434478 251290 434484 251292
rect 434345 251288 434484 251290
rect 434345 251232 434350 251288
rect 434406 251232 434484 251288
rect 434345 251230 434484 251232
rect 434345 251227 434411 251230
rect 434478 251228 434484 251230
rect 434548 251228 434554 251292
rect 255589 251154 255655 251157
rect 255773 251154 255839 251157
rect 255589 251152 255839 251154
rect 255589 251096 255594 251152
rect 255650 251096 255778 251152
rect 255834 251096 255839 251152
rect 255589 251094 255839 251096
rect 255589 251091 255655 251094
rect 255773 251091 255839 251094
rect 324589 251154 324655 251157
rect 324773 251154 324839 251157
rect 324589 251152 324839 251154
rect 324589 251096 324594 251152
rect 324650 251096 324778 251152
rect 324834 251096 324839 251152
rect 324589 251094 324839 251096
rect 324589 251091 324655 251094
rect 324773 251091 324839 251094
rect 254209 241498 254275 241501
rect 254393 241498 254459 241501
rect 254209 241496 254459 241498
rect 254209 241440 254214 241496
rect 254270 241440 254398 241496
rect 254454 241440 254459 241496
rect 254209 241438 254459 241440
rect 254209 241435 254275 241438
rect 254393 241435 254459 241438
rect 342345 241498 342411 241501
rect 342529 241498 342595 241501
rect 342345 241496 342595 241498
rect 342345 241440 342350 241496
rect 342406 241440 342534 241496
rect 342590 241440 342595 241496
rect 342345 241438 342595 241440
rect 342345 241435 342411 241438
rect 342529 241435 342595 241438
rect 362953 241498 363019 241501
rect 363137 241498 363203 241501
rect 362953 241496 363203 241498
rect 362953 241440 362958 241496
rect 363014 241440 363142 241496
rect 363198 241440 363203 241496
rect 362953 241438 363203 241440
rect 362953 241435 363019 241438
rect 363137 241435 363203 241438
rect 583520 240396 584960 240636
rect 229277 240138 229343 240141
rect 229553 240138 229619 240141
rect 229277 240136 229619 240138
rect 229277 240080 229282 240136
rect 229338 240080 229558 240136
rect 229614 240080 229619 240136
rect 229277 240078 229619 240080
rect 229277 240075 229343 240078
rect 229553 240075 229619 240078
rect 235073 240138 235139 240141
rect 235257 240138 235323 240141
rect 239121 240138 239187 240141
rect 235073 240136 235323 240138
rect 235073 240080 235078 240136
rect 235134 240080 235262 240136
rect 235318 240080 235323 240136
rect 235073 240078 235323 240080
rect 235073 240075 235139 240078
rect 235257 240075 235323 240078
rect 239078 240136 239187 240138
rect 239078 240080 239126 240136
rect 239182 240080 239187 240136
rect 239078 240075 239187 240080
rect 240225 240138 240291 240141
rect 240409 240138 240475 240141
rect 240225 240136 240475 240138
rect 240225 240080 240230 240136
rect 240286 240080 240414 240136
rect 240470 240080 240475 240136
rect 240225 240078 240475 240080
rect 240225 240075 240291 240078
rect 240409 240075 240475 240078
rect 241881 240138 241947 240141
rect 242065 240138 242131 240141
rect 241881 240136 242131 240138
rect 241881 240080 241886 240136
rect 241942 240080 242070 240136
rect 242126 240080 242131 240136
rect 241881 240078 242131 240080
rect 241881 240075 241947 240078
rect 242065 240075 242131 240078
rect 239078 240002 239138 240075
rect 239213 240002 239279 240005
rect 239078 240000 239279 240002
rect 239078 239944 239218 240000
rect 239274 239944 239279 240000
rect 239078 239942 239279 239944
rect 239213 239939 239279 239942
rect -960 237010 480 237100
rect 3969 237010 4035 237013
rect -960 237008 4035 237010
rect -960 236952 3974 237008
rect 4030 236952 4035 237008
rect -960 236950 4035 236952
rect -960 236860 480 236950
rect 3969 236947 4035 236950
rect 245745 231842 245811 231845
rect 245929 231842 245995 231845
rect 245745 231840 245995 231842
rect 245745 231784 245750 231840
rect 245806 231784 245934 231840
rect 245990 231784 245995 231840
rect 245745 231782 245995 231784
rect 245745 231779 245811 231782
rect 245929 231779 245995 231782
rect 324589 231842 324655 231845
rect 324865 231842 324931 231845
rect 324589 231840 324931 231842
rect 324589 231784 324594 231840
rect 324650 231784 324870 231840
rect 324926 231784 324931 231840
rect 324589 231782 324931 231784
rect 324589 231779 324655 231782
rect 324865 231779 324931 231782
rect 347957 231842 348023 231845
rect 348141 231842 348207 231845
rect 347957 231840 348207 231842
rect 347957 231784 347962 231840
rect 348018 231784 348146 231840
rect 348202 231784 348207 231840
rect 347957 231782 348207 231784
rect 347957 231779 348023 231782
rect 348141 231779 348207 231782
rect 291561 230482 291627 230485
rect 291745 230482 291811 230485
rect 291561 230480 291811 230482
rect 291561 230424 291566 230480
rect 291622 230424 291750 230480
rect 291806 230424 291811 230480
rect 291561 230422 291811 230424
rect 291561 230419 291627 230422
rect 291745 230419 291811 230422
rect 327349 230482 327415 230485
rect 327533 230482 327599 230485
rect 327349 230480 327599 230482
rect 327349 230424 327354 230480
rect 327410 230424 327538 230480
rect 327594 230424 327599 230480
rect 327349 230422 327599 230424
rect 327349 230419 327415 230422
rect 327533 230419 327599 230422
rect 310697 229122 310763 229125
rect 310973 229122 311039 229125
rect 310697 229120 311039 229122
rect 310697 229064 310702 229120
rect 310758 229064 310978 229120
rect 311034 229064 311039 229120
rect 310697 229062 311039 229064
rect 310697 229059 310763 229062
rect 310973 229059 311039 229062
rect 580809 228850 580875 228853
rect 583520 228850 584960 228940
rect 580809 228848 584960 228850
rect 580809 228792 580814 228848
rect 580870 228792 584960 228848
rect 580809 228790 584960 228792
rect 580809 228787 580875 228790
rect 583520 228700 584960 228790
rect -960 222594 480 222684
rect 3877 222594 3943 222597
rect -960 222592 3943 222594
rect -960 222536 3882 222592
rect 3938 222536 3943 222592
rect -960 222534 3943 222536
rect -960 222444 480 222534
rect 3877 222531 3943 222534
rect 254209 222186 254275 222189
rect 254393 222186 254459 222189
rect 254209 222184 254459 222186
rect 254209 222128 254214 222184
rect 254270 222128 254398 222184
rect 254454 222128 254459 222184
rect 254209 222126 254459 222128
rect 254209 222123 254275 222126
rect 254393 222123 254459 222126
rect 287329 222186 287395 222189
rect 287513 222186 287579 222189
rect 287329 222184 287579 222186
rect 287329 222128 287334 222184
rect 287390 222128 287518 222184
rect 287574 222128 287579 222184
rect 287329 222126 287579 222128
rect 287329 222123 287395 222126
rect 287513 222123 287579 222126
rect 342345 222186 342411 222189
rect 342529 222186 342595 222189
rect 342345 222184 342595 222186
rect 342345 222128 342350 222184
rect 342406 222128 342534 222184
rect 342590 222128 342595 222184
rect 342345 222126 342595 222128
rect 342345 222123 342411 222126
rect 342529 222123 342595 222126
rect 362953 222186 363019 222189
rect 363137 222186 363203 222189
rect 362953 222184 363203 222186
rect 362953 222128 362958 222184
rect 363014 222128 363142 222184
rect 363198 222128 363203 222184
rect 362953 222126 363203 222128
rect 362953 222123 363019 222126
rect 363137 222123 363203 222126
rect 234889 220826 234955 220829
rect 235165 220826 235231 220829
rect 239121 220826 239187 220829
rect 234889 220824 235231 220826
rect 234889 220768 234894 220824
rect 234950 220768 235170 220824
rect 235226 220768 235231 220824
rect 234889 220766 235231 220768
rect 234889 220763 234955 220766
rect 235165 220763 235231 220766
rect 239078 220824 239187 220826
rect 239078 220768 239126 220824
rect 239182 220768 239187 220824
rect 239078 220763 239187 220768
rect 240225 220826 240291 220829
rect 240409 220826 240475 220829
rect 240225 220824 240475 220826
rect 240225 220768 240230 220824
rect 240286 220768 240414 220824
rect 240470 220768 240475 220824
rect 240225 220766 240475 220768
rect 240225 220763 240291 220766
rect 240409 220763 240475 220766
rect 241881 220826 241947 220829
rect 242065 220826 242131 220829
rect 241881 220824 242131 220826
rect 241881 220768 241886 220824
rect 241942 220768 242070 220824
rect 242126 220768 242131 220824
rect 241881 220766 242131 220768
rect 241881 220763 241947 220766
rect 242065 220763 242131 220766
rect 239078 220693 239138 220763
rect 239029 220688 239138 220693
rect 239029 220632 239034 220688
rect 239090 220632 239138 220688
rect 239029 220630 239138 220632
rect 239029 220627 239095 220630
rect 251173 219466 251239 219469
rect 251357 219466 251423 219469
rect 251173 219464 251423 219466
rect 251173 219408 251178 219464
rect 251234 219408 251362 219464
rect 251418 219408 251423 219464
rect 251173 219406 251423 219408
rect 251173 219403 251239 219406
rect 251357 219403 251423 219406
rect 580717 217018 580783 217021
rect 583520 217018 584960 217108
rect 580717 217016 584960 217018
rect 580717 216960 580722 217016
rect 580778 216960 584960 217016
rect 580717 216958 584960 216960
rect 580717 216955 580783 216958
rect 583520 216868 584960 216958
rect 308029 212530 308095 212533
rect 308213 212530 308279 212533
rect 308029 212528 308279 212530
rect 308029 212472 308034 212528
rect 308090 212472 308218 212528
rect 308274 212472 308279 212528
rect 308029 212470 308279 212472
rect 308029 212467 308095 212470
rect 308213 212467 308279 212470
rect 347957 212530 348023 212533
rect 348141 212530 348207 212533
rect 347957 212528 348207 212530
rect 347957 212472 347962 212528
rect 348018 212472 348146 212528
rect 348202 212472 348207 212528
rect 347957 212470 348207 212472
rect 347957 212467 348023 212470
rect 348141 212467 348207 212470
rect 435173 212530 435239 212533
rect 435357 212530 435423 212533
rect 435173 212528 435423 212530
rect 435173 212472 435178 212528
rect 435234 212472 435362 212528
rect 435418 212472 435423 212528
rect 435173 212470 435423 212472
rect 435173 212467 435239 212470
rect 435357 212467 435423 212470
rect 234889 211170 234955 211173
rect 235165 211170 235231 211173
rect 234889 211168 235231 211170
rect 234889 211112 234894 211168
rect 234950 211112 235170 211168
rect 235226 211112 235231 211168
rect 234889 211110 235231 211112
rect 234889 211107 234955 211110
rect 235165 211107 235231 211110
rect 240225 211170 240291 211173
rect 240409 211170 240475 211173
rect 240225 211168 240475 211170
rect 240225 211112 240230 211168
rect 240286 211112 240414 211168
rect 240470 211112 240475 211168
rect 240225 211110 240475 211112
rect 240225 211107 240291 211110
rect 240409 211107 240475 211110
rect 241881 211170 241947 211173
rect 242065 211170 242131 211173
rect 241881 211168 242131 211170
rect 241881 211112 241886 211168
rect 241942 211112 242070 211168
rect 242126 211112 242131 211168
rect 241881 211110 242131 211112
rect 241881 211107 241947 211110
rect 242065 211107 242131 211110
rect 261201 211170 261267 211173
rect 261385 211170 261451 211173
rect 261201 211168 261451 211170
rect 261201 211112 261206 211168
rect 261262 211112 261390 211168
rect 261446 211112 261451 211168
rect 261201 211110 261451 211112
rect 261201 211107 261267 211110
rect 261385 211107 261451 211110
rect -960 208178 480 208268
rect 2773 208178 2839 208181
rect -960 208176 2839 208178
rect -960 208120 2778 208176
rect 2834 208120 2839 208176
rect -960 208118 2839 208120
rect -960 208028 480 208118
rect 2773 208115 2839 208118
rect 583520 205322 584960 205412
rect 583342 205262 584960 205322
rect 447726 204580 447732 204644
rect 447796 204642 447802 204644
rect 447796 204582 451290 204642
rect 447796 204580 447802 204582
rect 451230 204506 451290 204582
rect 460982 204582 470610 204642
rect 451230 204446 460858 204506
rect 460798 204370 460858 204446
rect 460982 204370 461042 204582
rect 470550 204506 470610 204582
rect 480302 204582 489930 204642
rect 470550 204446 480178 204506
rect 460798 204310 461042 204370
rect 480118 204370 480178 204446
rect 480302 204370 480362 204582
rect 489870 204506 489930 204582
rect 499622 204582 509250 204642
rect 489870 204446 499498 204506
rect 480118 204310 480362 204370
rect 499438 204370 499498 204446
rect 499622 204370 499682 204582
rect 509190 204506 509250 204582
rect 518942 204582 528570 204642
rect 509190 204446 518818 204506
rect 499438 204310 499682 204370
rect 518758 204370 518818 204446
rect 518942 204370 519002 204582
rect 528510 204506 528570 204582
rect 538262 204582 547890 204642
rect 528510 204446 538138 204506
rect 518758 204310 519002 204370
rect 538078 204370 538138 204446
rect 538262 204370 538322 204582
rect 547830 204506 547890 204582
rect 557582 204582 567210 204642
rect 547830 204446 557458 204506
rect 538078 204310 538322 204370
rect 557398 204370 557458 204446
rect 557582 204370 557642 204582
rect 567150 204506 567210 204582
rect 583342 204506 583402 205262
rect 583520 205172 584960 205262
rect 567150 204446 576778 204506
rect 557398 204310 557642 204370
rect 576718 204370 576778 204446
rect 576902 204446 583402 204506
rect 576902 204370 576962 204446
rect 576718 204310 576962 204370
rect 229277 202874 229343 202877
rect 229553 202874 229619 202877
rect 229277 202872 229619 202874
rect 229277 202816 229282 202872
rect 229338 202816 229558 202872
rect 229614 202816 229619 202872
rect 229277 202814 229619 202816
rect 229277 202811 229343 202814
rect 229553 202811 229619 202814
rect 244089 202874 244155 202877
rect 244273 202874 244339 202877
rect 244089 202872 244339 202874
rect 244089 202816 244094 202872
rect 244150 202816 244278 202872
rect 244334 202816 244339 202872
rect 244089 202814 244339 202816
rect 244089 202811 244155 202814
rect 244273 202811 244339 202814
rect 287329 202874 287395 202877
rect 287513 202874 287579 202877
rect 287329 202872 287579 202874
rect 287329 202816 287334 202872
rect 287390 202816 287518 202872
rect 287574 202816 287579 202872
rect 287329 202814 287579 202816
rect 287329 202811 287395 202814
rect 287513 202811 287579 202814
rect 362953 202874 363019 202877
rect 363137 202874 363203 202877
rect 362953 202872 363203 202874
rect 362953 202816 362958 202872
rect 363014 202816 363142 202872
rect 363198 202816 363203 202872
rect 362953 202814 363203 202816
rect 362953 202811 363019 202814
rect 363137 202811 363203 202814
rect 435173 202874 435239 202877
rect 435357 202874 435423 202877
rect 435173 202872 435423 202874
rect 435173 202816 435178 202872
rect 435234 202816 435362 202872
rect 435418 202816 435423 202872
rect 435173 202814 435423 202816
rect 435173 202811 435239 202814
rect 435357 202811 435423 202814
rect 309317 201514 309383 201517
rect 309501 201514 309567 201517
rect 309317 201512 309567 201514
rect 309317 201456 309322 201512
rect 309378 201456 309506 201512
rect 309562 201456 309567 201512
rect 309317 201454 309567 201456
rect 309317 201451 309383 201454
rect 309501 201451 309567 201454
rect 316309 201514 316375 201517
rect 316493 201514 316559 201517
rect 316309 201512 316559 201514
rect 316309 201456 316314 201512
rect 316370 201456 316498 201512
rect 316554 201456 316559 201512
rect 316309 201454 316559 201456
rect 316309 201451 316375 201454
rect 316493 201451 316559 201454
rect 327349 201514 327415 201517
rect 327533 201514 327599 201517
rect 327349 201512 327599 201514
rect 327349 201456 327354 201512
rect 327410 201456 327538 201512
rect 327594 201456 327599 201512
rect 327349 201454 327599 201456
rect 327349 201451 327415 201454
rect 327533 201451 327599 201454
rect 251541 200154 251607 200157
rect 251725 200154 251791 200157
rect 251541 200152 251791 200154
rect 251541 200096 251546 200152
rect 251602 200096 251730 200152
rect 251786 200096 251791 200152
rect 251541 200094 251791 200096
rect 251541 200091 251607 200094
rect 251725 200091 251791 200094
rect -960 193898 480 193988
rect 3785 193898 3851 193901
rect -960 193896 3851 193898
rect -960 193840 3790 193896
rect 3846 193840 3851 193896
rect -960 193838 3851 193840
rect -960 193748 480 193838
rect 3785 193835 3851 193838
rect 583520 193476 584960 193716
rect 308029 193218 308095 193221
rect 308305 193218 308371 193221
rect 308029 193216 308371 193218
rect 308029 193160 308034 193216
rect 308090 193160 308310 193216
rect 308366 193160 308371 193216
rect 308029 193158 308371 193160
rect 308029 193155 308095 193158
rect 308305 193155 308371 193158
rect 342345 193218 342411 193221
rect 342529 193218 342595 193221
rect 342345 193216 342595 193218
rect 342345 193160 342350 193216
rect 342406 193160 342534 193216
rect 342590 193160 342595 193216
rect 342345 193158 342595 193160
rect 342345 193155 342411 193158
rect 342529 193155 342595 193158
rect 347957 193218 348023 193221
rect 348141 193218 348207 193221
rect 347957 193216 348207 193218
rect 347957 193160 347962 193216
rect 348018 193160 348146 193216
rect 348202 193160 348207 193216
rect 347957 193158 348207 193160
rect 347957 193155 348023 193158
rect 348141 193155 348207 193158
rect 255681 191994 255747 191997
rect 255454 191992 255747 191994
rect 255454 191936 255686 191992
rect 255742 191936 255747 191992
rect 255454 191934 255747 191936
rect 254209 191858 254275 191861
rect 254393 191858 254459 191861
rect 254209 191856 254459 191858
rect 254209 191800 254214 191856
rect 254270 191800 254398 191856
rect 254454 191800 254459 191856
rect 254209 191798 254459 191800
rect 255454 191858 255514 191934
rect 255681 191931 255747 191934
rect 255589 191858 255655 191861
rect 255454 191856 255655 191858
rect 255454 191800 255594 191856
rect 255650 191800 255655 191856
rect 255454 191798 255655 191800
rect 254209 191795 254275 191798
rect 254393 191795 254459 191798
rect 255589 191795 255655 191798
rect 229277 183562 229343 183565
rect 229553 183562 229619 183565
rect 229277 183560 229619 183562
rect 229277 183504 229282 183560
rect 229338 183504 229558 183560
rect 229614 183504 229619 183560
rect 229277 183502 229619 183504
rect 229277 183499 229343 183502
rect 229553 183499 229619 183502
rect 291377 183562 291443 183565
rect 291561 183562 291627 183565
rect 291377 183560 291627 183562
rect 291377 183504 291382 183560
rect 291438 183504 291566 183560
rect 291622 183504 291627 183560
rect 291377 183502 291627 183504
rect 291377 183499 291443 183502
rect 291561 183499 291627 183502
rect 362953 183562 363019 183565
rect 363137 183562 363203 183565
rect 362953 183560 363203 183562
rect 362953 183504 362958 183560
rect 363014 183504 363142 183560
rect 363198 183504 363203 183560
rect 362953 183502 363203 183504
rect 362953 183499 363019 183502
rect 363137 183499 363203 183502
rect 443913 183562 443979 183565
rect 444097 183562 444163 183565
rect 443913 183560 444163 183562
rect 443913 183504 443918 183560
rect 443974 183504 444102 183560
rect 444158 183504 444163 183560
rect 443913 183502 444163 183504
rect 443913 183499 443979 183502
rect 444097 183499 444163 183502
rect 251449 182338 251515 182341
rect 251406 182336 251515 182338
rect 251406 182280 251454 182336
rect 251510 182280 251515 182336
rect 251406 182275 251515 182280
rect 251406 182066 251466 182275
rect 251633 182066 251699 182069
rect 251406 182064 251699 182066
rect 251406 182008 251638 182064
rect 251694 182008 251699 182064
rect 251406 182006 251699 182008
rect 251633 182003 251699 182006
rect 583520 181930 584960 182020
rect 583342 181870 584960 181930
rect 357382 181460 357388 181524
rect 357452 181522 357458 181524
rect 362125 181522 362191 181525
rect 357452 181520 362191 181522
rect 357452 181464 362130 181520
rect 362186 181464 362191 181520
rect 357452 181462 362191 181464
rect 357452 181460 357458 181462
rect 362125 181459 362191 181462
rect 326981 181386 327047 181389
rect 317462 181384 327047 181386
rect 317462 181328 326986 181384
rect 327042 181328 327047 181384
rect 317462 181326 327047 181328
rect 299238 181250 299244 181252
rect 292438 181190 299244 181250
rect 237782 181052 237788 181116
rect 237852 181114 237858 181116
rect 241462 181114 241468 181116
rect 237852 181054 241468 181114
rect 237852 181052 237858 181054
rect 241462 181052 241468 181054
rect 241532 181052 241538 181116
rect 275369 181114 275435 181117
rect 254534 181054 260850 181114
rect 241462 180780 241468 180844
rect 241532 180842 241538 180844
rect 254534 180842 254594 181054
rect 260790 180978 260850 181054
rect 275369 181112 284954 181114
rect 275369 181056 275374 181112
rect 275430 181056 284954 181112
rect 275369 181054 284954 181056
rect 275369 181051 275435 181054
rect 284894 180978 284954 181054
rect 292438 180978 292498 181190
rect 299238 181188 299244 181190
rect 299308 181188 299314 181252
rect 299422 181052 299428 181116
rect 299492 181114 299498 181116
rect 309041 181114 309107 181117
rect 299492 181112 309107 181114
rect 299492 181056 309046 181112
rect 309102 181056 309107 181112
rect 299492 181054 309107 181056
rect 299492 181052 299498 181054
rect 309041 181051 309107 181054
rect 312077 181114 312143 181117
rect 317462 181114 317522 181326
rect 326981 181323 327047 181326
rect 357382 181250 357388 181252
rect 350582 181190 357388 181250
rect 312077 181112 317522 181114
rect 312077 181056 312082 181112
rect 312138 181056 317522 181112
rect 312077 181054 317522 181056
rect 326981 181114 327047 181117
rect 326981 181112 331138 181114
rect 326981 181056 326986 181112
rect 327042 181056 331138 181112
rect 326981 181054 331138 181056
rect 312077 181051 312143 181054
rect 326981 181051 327047 181054
rect 260790 180918 261034 180978
rect 284894 180918 292498 180978
rect 331078 180978 331138 181054
rect 350582 180978 350642 181190
rect 357382 181188 357388 181190
rect 357452 181188 357458 181252
rect 376710 181190 386338 181250
rect 376710 180978 376770 181190
rect 331078 180918 331506 180978
rect 241532 180782 254594 180842
rect 260974 180842 261034 180918
rect 270493 180842 270559 180845
rect 260974 180840 270559 180842
rect 260974 180784 270498 180840
rect 270554 180784 270559 180840
rect 260974 180782 270559 180784
rect 241532 180780 241538 180782
rect 270493 180779 270559 180782
rect 310421 180842 310487 180845
rect 310789 180842 310855 180845
rect 310421 180840 310855 180842
rect 310421 180784 310426 180840
rect 310482 180784 310794 180840
rect 310850 180784 310855 180840
rect 310421 180782 310855 180784
rect 331446 180842 331506 180918
rect 342854 180918 350642 180978
rect 369902 180918 376770 180978
rect 342854 180842 342914 180918
rect 331446 180808 340706 180842
rect 340830 180808 342914 180842
rect 331446 180782 342914 180808
rect 362125 180842 362191 180845
rect 369902 180842 369962 180918
rect 362125 180840 369962 180842
rect 362125 180784 362130 180840
rect 362186 180784 369962 180840
rect 362125 180782 369962 180784
rect 386278 180842 386338 181190
rect 427678 181054 437490 181114
rect 398465 180978 398531 180981
rect 389222 180976 398531 180978
rect 389222 180920 398470 180976
rect 398526 180920 398531 180976
rect 389222 180918 398531 180920
rect 389222 180842 389282 180918
rect 398465 180915 398531 180918
rect 399017 180978 399083 180981
rect 417877 180978 417943 180981
rect 399017 180976 405658 180978
rect 399017 180920 399022 180976
rect 399078 180920 405658 180976
rect 399017 180918 405658 180920
rect 399017 180915 399083 180918
rect 386278 180782 389282 180842
rect 405598 180842 405658 180918
rect 408542 180976 417943 180978
rect 408542 180920 417882 180976
rect 417938 180920 417943 180976
rect 408542 180918 417943 180920
rect 408542 180842 408602 180918
rect 417877 180915 417943 180918
rect 418337 180978 418403 180981
rect 418337 180976 424978 180978
rect 418337 180920 418342 180976
rect 418398 180920 424978 180976
rect 418337 180918 424978 180920
rect 418337 180915 418403 180918
rect 405598 180782 408602 180842
rect 424918 180842 424978 180918
rect 427678 180842 427738 181054
rect 424918 180782 427738 180842
rect 437430 180842 437490 181054
rect 476070 181054 485698 181114
rect 454401 180978 454467 180981
rect 447182 180976 454467 180978
rect 447182 180920 454406 180976
rect 454462 180920 454467 180976
rect 447182 180918 454467 180920
rect 447182 180842 447242 180918
rect 454401 180915 454467 180918
rect 458357 180978 458423 180981
rect 458357 180976 466378 180978
rect 458357 180920 458362 180976
rect 458418 180920 466378 180976
rect 458357 180918 466378 180920
rect 458357 180915 458423 180918
rect 437430 180782 447242 180842
rect 466318 180842 466378 180918
rect 476070 180842 476130 181054
rect 466318 180782 476130 180842
rect 485638 180842 485698 181054
rect 495390 181054 505018 181114
rect 495390 180842 495450 181054
rect 485638 180782 495450 180842
rect 504958 180842 505018 181054
rect 514710 181054 524338 181114
rect 514710 180842 514770 181054
rect 504958 180782 514770 180842
rect 524278 180842 524338 181054
rect 528510 181054 547890 181114
rect 528510 180842 528570 181054
rect 547830 180978 547890 181054
rect 557582 181054 567210 181114
rect 547830 180918 557458 180978
rect 524278 180782 528570 180842
rect 557398 180842 557458 180918
rect 557582 180842 557642 181054
rect 567150 180978 567210 181054
rect 583342 180978 583402 181870
rect 583520 181780 584960 181870
rect 567150 180918 583402 180978
rect 557398 180782 557642 180842
rect 310421 180779 310487 180782
rect 310789 180779 310855 180782
rect 340646 180748 340890 180782
rect 362125 180779 362191 180782
rect -960 179482 480 179572
rect 2773 179482 2839 179485
rect -960 179480 2839 179482
rect -960 179424 2778 179480
rect 2834 179424 2839 179480
rect -960 179422 2839 179424
rect -960 179332 480 179422
rect 2773 179419 2839 179422
rect 240409 173906 240475 173909
rect 240593 173906 240659 173909
rect 240409 173904 240659 173906
rect 240409 173848 240414 173904
rect 240470 173848 240598 173904
rect 240654 173848 240659 173904
rect 240409 173846 240659 173848
rect 240409 173843 240475 173846
rect 240593 173843 240659 173846
rect 291469 173906 291535 173909
rect 291745 173906 291811 173909
rect 291469 173904 291811 173906
rect 291469 173848 291474 173904
rect 291530 173848 291750 173904
rect 291806 173848 291811 173904
rect 291469 173846 291811 173848
rect 291469 173843 291535 173846
rect 291745 173843 291811 173846
rect 347957 173906 348023 173909
rect 348141 173906 348207 173909
rect 434345 173908 434411 173909
rect 347957 173904 348207 173906
rect 347957 173848 347962 173904
rect 348018 173848 348146 173904
rect 348202 173848 348207 173904
rect 347957 173846 348207 173848
rect 347957 173843 348023 173846
rect 348141 173843 348207 173846
rect 434294 173844 434300 173908
rect 434364 173906 434411 173908
rect 434364 173904 434456 173906
rect 434406 173848 434456 173904
rect 434364 173846 434456 173848
rect 434364 173844 434411 173846
rect 434345 173843 434411 173844
rect 251449 172546 251515 172549
rect 251633 172546 251699 172549
rect 251449 172544 251699 172546
rect 251449 172488 251454 172544
rect 251510 172488 251638 172544
rect 251694 172488 251699 172544
rect 251449 172486 251699 172488
rect 251449 172483 251515 172486
rect 251633 172483 251699 172486
rect 324497 172546 324563 172549
rect 324681 172546 324747 172549
rect 324497 172544 324747 172546
rect 324497 172488 324502 172544
rect 324558 172488 324686 172544
rect 324742 172488 324747 172544
rect 324497 172486 324747 172488
rect 324497 172483 324563 172486
rect 324681 172483 324747 172486
rect 343909 172546 343975 172549
rect 344093 172546 344159 172549
rect 343909 172544 344159 172546
rect 343909 172488 343914 172544
rect 343970 172488 344098 172544
rect 344154 172488 344159 172544
rect 343909 172486 344159 172488
rect 343909 172483 343975 172486
rect 344093 172483 344159 172486
rect 345013 172546 345079 172549
rect 345289 172546 345355 172549
rect 345013 172544 345355 172546
rect 345013 172488 345018 172544
rect 345074 172488 345294 172544
rect 345350 172488 345355 172544
rect 345013 172486 345355 172488
rect 345013 172483 345079 172486
rect 345289 172483 345355 172486
rect 580625 170098 580691 170101
rect 583520 170098 584960 170188
rect 580625 170096 584960 170098
rect 580625 170040 580630 170096
rect 580686 170040 584960 170096
rect 580625 170038 584960 170040
rect 580625 170035 580691 170038
rect 583520 169948 584960 170038
rect -960 165066 480 165156
rect 2773 165066 2839 165069
rect -960 165064 2839 165066
rect -960 165008 2778 165064
rect 2834 165008 2839 165064
rect -960 165006 2839 165008
rect -960 164916 480 165006
rect 2773 165003 2839 165006
rect 342529 164386 342595 164389
rect 343909 164386 343975 164389
rect 342529 164384 342730 164386
rect 342529 164328 342534 164384
rect 342590 164328 342730 164384
rect 342529 164326 342730 164328
rect 342529 164323 342595 164326
rect 239121 164250 239187 164253
rect 239305 164250 239371 164253
rect 239121 164248 239371 164250
rect 239121 164192 239126 164248
rect 239182 164192 239310 164248
rect 239366 164192 239371 164248
rect 239121 164190 239371 164192
rect 239121 164187 239187 164190
rect 239305 164187 239371 164190
rect 266997 164250 267063 164253
rect 291561 164250 291627 164253
rect 291745 164250 291811 164253
rect 266997 164248 267290 164250
rect 266997 164192 267002 164248
rect 267058 164192 267290 164248
rect 266997 164190 267290 164192
rect 266997 164187 267063 164190
rect 267230 164117 267290 164190
rect 291561 164248 291811 164250
rect 291561 164192 291566 164248
rect 291622 164192 291750 164248
rect 291806 164192 291811 164248
rect 291561 164190 291811 164192
rect 291561 164187 291627 164190
rect 291745 164187 291811 164190
rect 342529 164250 342595 164253
rect 342670 164250 342730 164326
rect 342529 164248 342730 164250
rect 342529 164192 342534 164248
rect 342590 164192 342730 164248
rect 342529 164190 342730 164192
rect 343774 164384 343975 164386
rect 343774 164328 343914 164384
rect 343970 164328 343975 164384
rect 343774 164326 343975 164328
rect 343774 164250 343834 164326
rect 343909 164323 343975 164326
rect 343909 164250 343975 164253
rect 343774 164248 343975 164250
rect 343774 164192 343914 164248
rect 343970 164192 343975 164248
rect 343774 164190 343975 164192
rect 342529 164187 342595 164190
rect 343909 164187 343975 164190
rect 347957 164250 348023 164253
rect 348141 164250 348207 164253
rect 347957 164248 348207 164250
rect 347957 164192 347962 164248
rect 348018 164192 348146 164248
rect 348202 164192 348207 164248
rect 347957 164190 348207 164192
rect 347957 164187 348023 164190
rect 348141 164187 348207 164190
rect 434294 164188 434300 164252
rect 434364 164250 434370 164252
rect 434437 164250 434503 164253
rect 434364 164248 434503 164250
rect 434364 164192 434442 164248
rect 434498 164192 434503 164248
rect 434364 164190 434503 164192
rect 434364 164188 434370 164190
rect 434437 164187 434503 164190
rect 267230 164112 267339 164117
rect 267230 164056 267278 164112
rect 267334 164056 267339 164112
rect 267230 164054 267339 164056
rect 267273 164051 267339 164054
rect 234889 162890 234955 162893
rect 235073 162890 235139 162893
rect 234889 162888 235139 162890
rect 234889 162832 234894 162888
rect 234950 162832 235078 162888
rect 235134 162832 235139 162888
rect 234889 162830 235139 162832
rect 234889 162827 234955 162830
rect 235073 162827 235139 162830
rect 580533 158402 580599 158405
rect 583520 158402 584960 158492
rect 580533 158400 584960 158402
rect 580533 158344 580538 158400
rect 580594 158344 584960 158400
rect 580533 158342 584960 158344
rect 580533 158339 580599 158342
rect 583520 158252 584960 158342
rect 291561 154730 291627 154733
rect 291518 154728 291627 154730
rect 291518 154672 291566 154728
rect 291622 154672 291627 154728
rect 291518 154667 291627 154672
rect 254209 154594 254275 154597
rect 254393 154594 254459 154597
rect 254209 154592 254459 154594
rect 254209 154536 254214 154592
rect 254270 154536 254398 154592
rect 254454 154536 254459 154592
rect 254209 154534 254459 154536
rect 254209 154531 254275 154534
rect 254393 154531 254459 154534
rect 266997 154594 267063 154597
rect 267273 154594 267339 154597
rect 266997 154592 267339 154594
rect 266997 154536 267002 154592
rect 267058 154536 267278 154592
rect 267334 154536 267339 154592
rect 266997 154534 267339 154536
rect 266997 154531 267063 154534
rect 267273 154531 267339 154534
rect 291518 154458 291578 154667
rect 362953 154594 363019 154597
rect 363229 154594 363295 154597
rect 362953 154592 363295 154594
rect 362953 154536 362958 154592
rect 363014 154536 363234 154592
rect 363290 154536 363295 154592
rect 362953 154534 363295 154536
rect 362953 154531 363019 154534
rect 363229 154531 363295 154534
rect 291653 154458 291719 154461
rect 291518 154456 291719 154458
rect 291518 154400 291658 154456
rect 291714 154400 291719 154456
rect 291518 154398 291719 154400
rect 291653 154395 291719 154398
rect -960 150786 480 150876
rect 3693 150786 3759 150789
rect -960 150784 3759 150786
rect -960 150728 3698 150784
rect 3754 150728 3759 150784
rect -960 150726 3759 150728
rect -960 150636 480 150726
rect 3693 150723 3759 150726
rect 583520 146556 584960 146796
rect 229277 144938 229343 144941
rect 229553 144938 229619 144941
rect 229277 144936 229619 144938
rect 229277 144880 229282 144936
rect 229338 144880 229558 144936
rect 229614 144880 229619 144936
rect 229277 144878 229619 144880
rect 229277 144875 229343 144878
rect 229553 144875 229619 144878
rect 245745 144938 245811 144941
rect 245929 144938 245995 144941
rect 245745 144936 245995 144938
rect 245745 144880 245750 144936
rect 245806 144880 245934 144936
rect 245990 144880 245995 144936
rect 245745 144878 245995 144880
rect 245745 144875 245811 144878
rect 245929 144875 245995 144878
rect 262489 144938 262555 144941
rect 262673 144938 262739 144941
rect 262489 144936 262739 144938
rect 262489 144880 262494 144936
rect 262550 144880 262678 144936
rect 262734 144880 262739 144936
rect 262489 144878 262739 144880
rect 262489 144875 262555 144878
rect 262673 144875 262739 144878
rect 324589 144938 324655 144941
rect 324773 144938 324839 144941
rect 324589 144936 324839 144938
rect 324589 144880 324594 144936
rect 324650 144880 324778 144936
rect 324834 144880 324839 144936
rect 324589 144878 324839 144880
rect 324589 144875 324655 144878
rect 324773 144875 324839 144878
rect 347957 144938 348023 144941
rect 348141 144938 348207 144941
rect 347957 144936 348207 144938
rect 347957 144880 347962 144936
rect 348018 144880 348146 144936
rect 348202 144880 348207 144936
rect 347957 144878 348207 144880
rect 347957 144875 348023 144878
rect 348141 144875 348207 144878
rect 235073 143714 235139 143717
rect 235030 143712 235139 143714
rect 235030 143656 235078 143712
rect 235134 143656 235139 143712
rect 235030 143651 235139 143656
rect 235030 143578 235090 143651
rect 235165 143578 235231 143581
rect 235030 143576 235231 143578
rect 235030 143520 235170 143576
rect 235226 143520 235231 143576
rect 235030 143518 235231 143520
rect 235165 143515 235231 143518
rect 251173 143578 251239 143581
rect 251357 143578 251423 143581
rect 251173 143576 251423 143578
rect 251173 143520 251178 143576
rect 251234 143520 251362 143576
rect 251418 143520 251423 143576
rect 251173 143518 251423 143520
rect 251173 143515 251239 143518
rect 251357 143515 251423 143518
rect 255313 143578 255379 143581
rect 255497 143578 255563 143581
rect 255313 143576 255563 143578
rect 255313 143520 255318 143576
rect 255374 143520 255502 143576
rect 255558 143520 255563 143576
rect 255313 143518 255563 143520
rect 255313 143515 255379 143518
rect 255497 143515 255563 143518
rect 434529 143578 434595 143581
rect 434713 143578 434779 143581
rect 434529 143576 434779 143578
rect 434529 143520 434534 143576
rect 434590 143520 434718 143576
rect 434774 143520 434779 143576
rect 434529 143518 434779 143520
rect 434529 143515 434595 143518
rect 434713 143515 434779 143518
rect 327441 138276 327507 138277
rect 327390 138274 327396 138276
rect 327350 138214 327396 138274
rect 327460 138272 327507 138276
rect 327502 138216 327507 138272
rect 327390 138212 327396 138214
rect 327460 138212 327507 138216
rect 327441 138211 327507 138212
rect -960 136370 480 136460
rect 2773 136370 2839 136373
rect -960 136368 2839 136370
rect -960 136312 2778 136368
rect 2834 136312 2839 136368
rect -960 136310 2839 136312
rect -960 136220 480 136310
rect 2773 136307 2839 136310
rect 290181 135418 290247 135421
rect 291561 135418 291627 135421
rect 324773 135418 324839 135421
rect 290046 135416 290247 135418
rect 290046 135360 290186 135416
rect 290242 135360 290247 135416
rect 290046 135358 290247 135360
rect 290046 135285 290106 135358
rect 290181 135355 290247 135358
rect 291518 135416 291627 135418
rect 291518 135360 291566 135416
rect 291622 135360 291627 135416
rect 291518 135355 291627 135360
rect 324454 135416 324839 135418
rect 324454 135360 324778 135416
rect 324834 135360 324839 135416
rect 324454 135358 324839 135360
rect 244089 135282 244155 135285
rect 244273 135282 244339 135285
rect 244089 135280 244339 135282
rect 244089 135224 244094 135280
rect 244150 135224 244278 135280
rect 244334 135224 244339 135280
rect 244089 135222 244339 135224
rect 244089 135219 244155 135222
rect 244273 135219 244339 135222
rect 254209 135282 254275 135285
rect 254393 135282 254459 135285
rect 254209 135280 254459 135282
rect 254209 135224 254214 135280
rect 254270 135224 254398 135280
rect 254454 135224 254459 135280
rect 254209 135222 254459 135224
rect 290046 135280 290155 135285
rect 290046 135224 290094 135280
rect 290150 135224 290155 135280
rect 290046 135222 290155 135224
rect 254209 135219 254275 135222
rect 254393 135219 254459 135222
rect 290089 135219 290155 135222
rect 291518 135149 291578 135355
rect 324454 135282 324514 135358
rect 324773 135355 324839 135358
rect 324589 135282 324655 135285
rect 327349 135284 327415 135285
rect 327349 135282 327396 135284
rect 324454 135280 324655 135282
rect 324454 135224 324594 135280
rect 324650 135224 324655 135280
rect 324454 135222 324655 135224
rect 327304 135280 327396 135282
rect 327304 135224 327354 135280
rect 327304 135222 327396 135224
rect 324589 135219 324655 135222
rect 327349 135220 327396 135222
rect 327460 135220 327466 135284
rect 362953 135282 363019 135285
rect 363229 135282 363295 135285
rect 362953 135280 363295 135282
rect 362953 135224 362958 135280
rect 363014 135224 363234 135280
rect 363290 135224 363295 135280
rect 362953 135222 363295 135224
rect 327349 135219 327415 135220
rect 362953 135219 363019 135222
rect 363229 135219 363295 135222
rect 291518 135144 291627 135149
rect 291518 135088 291566 135144
rect 291622 135088 291627 135144
rect 291518 135086 291627 135088
rect 291561 135083 291627 135086
rect 583520 134874 584960 134964
rect 583342 134814 584960 134874
rect 453982 134540 453988 134604
rect 454052 134602 454058 134604
rect 460841 134602 460907 134605
rect 454052 134600 460907 134602
rect 454052 134544 460846 134600
rect 460902 134544 460907 134600
rect 454052 134542 460907 134544
rect 454052 134540 454058 134542
rect 460841 134539 460907 134542
rect 447225 134330 447291 134333
rect 453982 134330 453988 134332
rect 376710 134270 386338 134330
rect 260741 134194 260807 134197
rect 269113 134194 269179 134197
rect 260741 134192 269179 134194
rect 260741 134136 260746 134192
rect 260802 134136 269118 134192
rect 269174 134136 269179 134192
rect 260741 134134 269179 134136
rect 260741 134131 260807 134134
rect 269113 134131 269179 134134
rect 336641 134194 336707 134197
rect 336641 134192 340522 134194
rect 336641 134136 336646 134192
rect 336702 134136 340522 134192
rect 336641 134134 340522 134136
rect 336641 134131 336707 134134
rect 275369 134058 275435 134061
rect 282729 134058 282795 134061
rect 275369 134056 282795 134058
rect 275369 134000 275374 134056
rect 275430 134000 282734 134056
rect 282790 134000 282795 134056
rect 275369 133998 282795 134000
rect 275369 133995 275435 133998
rect 282729 133995 282795 133998
rect 282913 134058 282979 134061
rect 309041 134058 309107 134061
rect 317505 134058 317571 134061
rect 282913 134056 283666 134058
rect 282913 134000 282918 134056
rect 282974 134000 283666 134056
rect 282913 133998 283666 134000
rect 282913 133995 282979 133998
rect 237966 133860 237972 133924
rect 238036 133922 238042 133924
rect 251173 133922 251239 133925
rect 238036 133920 251239 133922
rect 238036 133864 251178 133920
rect 251234 133864 251239 133920
rect 238036 133862 251239 133864
rect 283606 133922 283666 133998
rect 309041 134056 317571 134058
rect 309041 134000 309046 134056
rect 309102 134000 317510 134056
rect 317566 134000 317571 134056
rect 309041 133998 317571 134000
rect 309041 133995 309107 133998
rect 317505 133995 317571 133998
rect 326981 133922 327047 133925
rect 327257 133922 327323 133925
rect 283606 133862 289922 133922
rect 238036 133860 238042 133862
rect 251173 133859 251239 133862
rect 289862 133786 289922 133862
rect 326981 133920 327323 133922
rect 326981 133864 326986 133920
rect 327042 133864 327262 133920
rect 327318 133864 327323 133920
rect 326981 133862 327323 133864
rect 340462 133922 340522 134134
rect 357433 134058 357499 134061
rect 350582 134056 357499 134058
rect 350582 134000 357438 134056
rect 357494 134000 357499 134056
rect 350582 133998 357499 134000
rect 350582 133922 350642 133998
rect 357433 133995 357499 133998
rect 361113 134058 361179 134061
rect 376710 134058 376770 134270
rect 361113 134056 367018 134058
rect 361113 134000 361118 134056
rect 361174 134000 367018 134056
rect 361113 133998 367018 134000
rect 361113 133995 361179 133998
rect 340462 133862 350642 133922
rect 366958 133922 367018 133998
rect 369902 133998 376770 134058
rect 369902 133922 369962 133998
rect 366958 133862 369962 133922
rect 386278 133922 386338 134270
rect 447225 134328 453988 134330
rect 447225 134272 447230 134328
rect 447286 134272 453988 134328
rect 447225 134270 453988 134272
rect 447225 134267 447291 134270
rect 453982 134268 453988 134270
rect 454052 134268 454058 134332
rect 460841 134194 460907 134197
rect 460841 134192 470610 134194
rect 460841 134136 460846 134192
rect 460902 134136 470610 134192
rect 460841 134134 470610 134136
rect 460841 134131 460907 134134
rect 398465 134058 398531 134061
rect 389222 134056 398531 134058
rect 389222 134000 398470 134056
rect 398526 134000 398531 134056
rect 389222 133998 398531 134000
rect 389222 133922 389282 133998
rect 398465 133995 398531 133998
rect 399017 134058 399083 134061
rect 417877 134058 417943 134061
rect 399017 134056 405658 134058
rect 399017 134000 399022 134056
rect 399078 134000 405658 134056
rect 399017 133998 405658 134000
rect 399017 133995 399083 133998
rect 386278 133862 389282 133922
rect 405598 133922 405658 133998
rect 408542 134056 417943 134058
rect 408542 134000 417882 134056
rect 417938 134000 417943 134056
rect 408542 133998 417943 134000
rect 408542 133922 408602 133998
rect 417877 133995 417943 133998
rect 418337 134058 418403 134061
rect 447133 134058 447199 134061
rect 418337 134056 424978 134058
rect 418337 134000 418342 134056
rect 418398 134000 424978 134056
rect 418337 133998 424978 134000
rect 418337 133995 418403 133998
rect 405598 133862 408602 133922
rect 424918 133922 424978 133998
rect 427862 134056 447199 134058
rect 427862 134000 447138 134056
rect 447194 134000 447199 134056
rect 427862 133998 447199 134000
rect 470550 134058 470610 134134
rect 480302 134134 489930 134194
rect 470550 133998 480178 134058
rect 427862 133922 427922 133998
rect 447133 133995 447199 133998
rect 424918 133862 427922 133922
rect 480118 133922 480178 133998
rect 480302 133922 480362 134134
rect 489870 134058 489930 134134
rect 499622 134134 509250 134194
rect 489870 133998 499498 134058
rect 480118 133862 480362 133922
rect 499438 133922 499498 133998
rect 499622 133922 499682 134134
rect 509190 134058 509250 134134
rect 518942 134134 528570 134194
rect 509190 133998 518818 134058
rect 499438 133862 499682 133922
rect 518758 133922 518818 133998
rect 518942 133922 519002 134134
rect 528510 134058 528570 134134
rect 538262 134134 547890 134194
rect 528510 133998 538138 134058
rect 518758 133862 519002 133922
rect 538078 133922 538138 133998
rect 538262 133922 538322 134134
rect 547830 134058 547890 134134
rect 557582 134134 567210 134194
rect 547830 133998 557458 134058
rect 538078 133862 538322 133922
rect 557398 133922 557458 133998
rect 557582 133922 557642 134134
rect 567150 134058 567210 134134
rect 583342 134058 583402 134814
rect 583520 134724 584960 134814
rect 567150 133998 576778 134058
rect 557398 133862 557642 133922
rect 576718 133922 576778 133998
rect 576902 133998 583402 134058
rect 576902 133922 576962 133998
rect 576718 133862 576962 133922
rect 326981 133859 327047 133862
rect 327257 133859 327323 133862
rect 309041 133786 309107 133789
rect 289862 133784 309107 133786
rect 289862 133728 309046 133784
rect 309102 133728 309107 133784
rect 289862 133726 309107 133728
rect 309041 133723 309107 133726
rect 261385 125762 261451 125765
rect 261342 125760 261451 125762
rect 261342 125704 261390 125760
rect 261446 125704 261451 125760
rect 261342 125699 261451 125704
rect 261342 125629 261402 125699
rect 229277 125626 229343 125629
rect 229553 125626 229619 125629
rect 229277 125624 229619 125626
rect 229277 125568 229282 125624
rect 229338 125568 229558 125624
rect 229614 125568 229619 125624
rect 229277 125566 229619 125568
rect 229277 125563 229343 125566
rect 229553 125563 229619 125566
rect 245745 125626 245811 125629
rect 245929 125626 245995 125629
rect 245745 125624 245995 125626
rect 245745 125568 245750 125624
rect 245806 125568 245934 125624
rect 245990 125568 245995 125624
rect 245745 125566 245995 125568
rect 245745 125563 245811 125566
rect 245929 125563 245995 125566
rect 261293 125624 261402 125629
rect 261293 125568 261298 125624
rect 261354 125568 261402 125624
rect 261293 125566 261402 125568
rect 328453 125626 328519 125629
rect 328729 125626 328795 125629
rect 328453 125624 328795 125626
rect 328453 125568 328458 125624
rect 328514 125568 328734 125624
rect 328790 125568 328795 125624
rect 328453 125566 328795 125568
rect 261293 125563 261359 125566
rect 328453 125563 328519 125566
rect 328729 125563 328795 125566
rect 347957 125626 348023 125629
rect 348141 125626 348207 125629
rect 347957 125624 348207 125626
rect 347957 125568 347962 125624
rect 348018 125568 348146 125624
rect 348202 125568 348207 125624
rect 347957 125566 348207 125568
rect 347957 125563 348023 125566
rect 348141 125563 348207 125566
rect 287237 124266 287303 124269
rect 287513 124266 287579 124269
rect 287237 124264 287579 124266
rect 287237 124208 287242 124264
rect 287298 124208 287518 124264
rect 287574 124208 287579 124264
rect 287237 124206 287579 124208
rect 287237 124203 287303 124206
rect 287513 124203 287579 124206
rect 580441 123178 580507 123181
rect 583520 123178 584960 123268
rect 580441 123176 584960 123178
rect 580441 123120 580446 123176
rect 580502 123120 584960 123176
rect 580441 123118 584960 123120
rect 580441 123115 580507 123118
rect 583520 123028 584960 123118
rect -960 122090 480 122180
rect 2773 122090 2839 122093
rect -960 122088 2839 122090
rect -960 122032 2778 122088
rect 2834 122032 2839 122088
rect -960 122030 2839 122032
rect -960 121940 480 122030
rect 2773 122027 2839 122030
rect 324681 115970 324747 115973
rect 324865 115970 324931 115973
rect 324681 115968 324931 115970
rect 324681 115912 324686 115968
rect 324742 115912 324870 115968
rect 324926 115912 324931 115968
rect 324681 115910 324931 115912
rect 324681 115907 324747 115910
rect 324865 115907 324931 115910
rect 362953 115970 363019 115973
rect 363229 115970 363295 115973
rect 362953 115968 363295 115970
rect 362953 115912 362958 115968
rect 363014 115912 363234 115968
rect 363290 115912 363295 115968
rect 362953 115910 363295 115912
rect 362953 115907 363019 115910
rect 363229 115907 363295 115910
rect 342529 114610 342595 114613
rect 342713 114610 342779 114613
rect 342529 114608 342779 114610
rect 342529 114552 342534 114608
rect 342590 114552 342718 114608
rect 342774 114552 342779 114608
rect 342529 114550 342779 114552
rect 342529 114547 342595 114550
rect 342713 114547 342779 114550
rect 304993 113250 305059 113253
rect 305269 113250 305335 113253
rect 304993 113248 305335 113250
rect 304993 113192 304998 113248
rect 305054 113192 305274 113248
rect 305330 113192 305335 113248
rect 304993 113190 305335 113192
rect 304993 113187 305059 113190
rect 305269 113187 305335 113190
rect 580349 111482 580415 111485
rect 583520 111482 584960 111572
rect 580349 111480 584960 111482
rect 580349 111424 580354 111480
rect 580410 111424 584960 111480
rect 580349 111422 584960 111424
rect 580349 111419 580415 111422
rect 583520 111332 584960 111422
rect -960 107674 480 107764
rect 3601 107674 3667 107677
rect -960 107672 3667 107674
rect -960 107616 3606 107672
rect 3662 107616 3667 107672
rect -960 107614 3667 107616
rect -960 107524 480 107614
rect 3601 107611 3667 107614
rect 327533 106450 327599 106453
rect 327398 106448 327599 106450
rect 327398 106392 327538 106448
rect 327594 106392 327599 106448
rect 327398 106390 327599 106392
rect 327398 106317 327458 106390
rect 327533 106387 327599 106390
rect 241605 106314 241671 106317
rect 241789 106314 241855 106317
rect 241605 106312 241855 106314
rect 241605 106256 241610 106312
rect 241666 106256 241794 106312
rect 241850 106256 241855 106312
rect 241605 106254 241855 106256
rect 327398 106312 327507 106317
rect 327398 106256 327446 106312
rect 327502 106256 327507 106312
rect 327398 106254 327507 106256
rect 241605 106251 241671 106254
rect 241789 106251 241855 106254
rect 327441 106251 327507 106254
rect 347957 106314 348023 106317
rect 348141 106314 348207 106317
rect 347957 106312 348207 106314
rect 347957 106256 347962 106312
rect 348018 106256 348146 106312
rect 348202 106256 348207 106312
rect 347957 106254 348207 106256
rect 347957 106251 348023 106254
rect 348141 106251 348207 106254
rect 251357 105090 251423 105093
rect 251357 105088 251650 105090
rect 251357 105032 251362 105088
rect 251418 105032 251650 105088
rect 251357 105030 251650 105032
rect 251357 105027 251423 105030
rect 251449 104954 251515 104957
rect 251590 104954 251650 105030
rect 251449 104952 251650 104954
rect 251449 104896 251454 104952
rect 251510 104896 251650 104952
rect 251449 104894 251650 104896
rect 251449 104891 251515 104894
rect 291561 102098 291627 102101
rect 291561 102096 291762 102098
rect 291561 102040 291566 102096
rect 291622 102040 291762 102096
rect 291561 102038 291762 102040
rect 291561 102035 291627 102038
rect 291469 101962 291535 101965
rect 291702 101962 291762 102038
rect 291469 101960 291762 101962
rect 291469 101904 291474 101960
rect 291530 101904 291762 101960
rect 291469 101902 291762 101904
rect 291469 101899 291535 101902
rect 583520 99636 584960 99876
rect 362953 96658 363019 96661
rect 363229 96658 363295 96661
rect 362953 96656 363295 96658
rect 362953 96600 362958 96656
rect 363014 96600 363234 96656
rect 363290 96600 363295 96656
rect 362953 96598 363295 96600
rect 362953 96595 363019 96598
rect 363229 96595 363295 96598
rect 311065 93938 311131 93941
rect 311022 93936 311131 93938
rect 311022 93880 311070 93936
rect 311126 93880 311131 93936
rect 311022 93875 311131 93880
rect 311022 93805 311082 93875
rect 310973 93800 311082 93805
rect 310973 93744 310978 93800
rect 311034 93744 311082 93800
rect 310973 93742 311082 93744
rect 310973 93739 311039 93742
rect -960 93258 480 93348
rect 3509 93258 3575 93261
rect -960 93256 3575 93258
rect -960 93200 3514 93256
rect 3570 93200 3575 93256
rect -960 93198 3575 93200
rect -960 93108 480 93198
rect 3509 93195 3575 93198
rect 238150 91156 238156 91220
rect 238220 91218 238226 91220
rect 240041 91218 240107 91221
rect 238220 91216 240107 91218
rect 238220 91160 240046 91216
rect 240102 91160 240107 91216
rect 238220 91158 240107 91160
rect 238220 91156 238226 91158
rect 240041 91155 240107 91158
rect 583520 87954 584960 88044
rect 583342 87894 584960 87954
rect 299422 87484 299428 87548
rect 299492 87546 299498 87548
rect 299492 87486 312554 87546
rect 299492 87484 299498 87486
rect 254534 87214 263610 87274
rect 240041 87138 240107 87141
rect 253749 87138 253815 87141
rect 240041 87136 253815 87138
rect 240041 87080 240046 87136
rect 240102 87080 253754 87136
rect 253810 87080 253815 87136
rect 240041 87078 253815 87080
rect 240041 87075 240107 87078
rect 253749 87075 253815 87078
rect 253933 87138 253999 87141
rect 254534 87138 254594 87214
rect 253933 87136 254594 87138
rect 253933 87080 253938 87136
rect 253994 87080 254594 87136
rect 253933 87078 254594 87080
rect 253933 87075 253999 87078
rect 263550 87002 263610 87214
rect 269062 87212 269068 87276
rect 269132 87274 269138 87276
rect 282821 87274 282887 87277
rect 269132 87272 282887 87274
rect 269132 87216 282826 87272
rect 282882 87216 282887 87272
rect 269132 87214 282887 87216
rect 269132 87212 269138 87214
rect 282821 87211 282887 87214
rect 292757 87274 292823 87277
rect 299422 87274 299428 87276
rect 292757 87272 299428 87274
rect 292757 87216 292762 87272
rect 292818 87216 299428 87272
rect 292757 87214 299428 87216
rect 292757 87211 292823 87214
rect 299422 87212 299428 87214
rect 299492 87212 299498 87276
rect 312494 87274 312554 87486
rect 453982 87484 453988 87548
rect 454052 87546 454058 87548
rect 463601 87546 463667 87549
rect 454052 87544 463667 87546
rect 454052 87488 463606 87544
rect 463662 87488 463667 87544
rect 454052 87486 463667 87488
rect 454052 87484 454058 87486
rect 463601 87483 463667 87486
rect 365621 87410 365687 87413
rect 366950 87410 366956 87412
rect 365621 87408 366956 87410
rect 365621 87352 365626 87408
rect 365682 87352 366956 87408
rect 365621 87350 366956 87352
rect 365621 87347 365687 87350
rect 366950 87348 366956 87350
rect 367020 87348 367026 87412
rect 379286 87350 386338 87410
rect 317454 87274 317460 87276
rect 312494 87214 317460 87274
rect 317454 87212 317460 87214
rect 317524 87212 317530 87276
rect 326981 87274 327047 87277
rect 336641 87274 336707 87277
rect 326981 87272 336707 87274
rect 326981 87216 326986 87272
rect 327042 87216 336646 87272
rect 336702 87216 336707 87272
rect 326981 87214 336707 87216
rect 326981 87211 327047 87214
rect 336641 87211 336707 87214
rect 356053 87138 356119 87141
rect 379286 87138 379346 87350
rect 340462 87136 356119 87138
rect 340462 87080 356058 87136
rect 356114 87080 356119 87136
rect 340462 87078 356119 87080
rect 269062 87002 269068 87004
rect 263550 86942 269068 87002
rect 269062 86940 269068 86942
rect 269132 86940 269138 87004
rect 307937 87002 308003 87005
rect 308121 87002 308187 87005
rect 307937 87000 308187 87002
rect 307937 86944 307942 87000
rect 307998 86944 308126 87000
rect 308182 86944 308187 87000
rect 307937 86942 308187 86944
rect 307937 86939 308003 86942
rect 308121 86939 308187 86942
rect 317454 86940 317460 87004
rect 317524 87002 317530 87004
rect 326981 87002 327047 87005
rect 317524 87000 327047 87002
rect 317524 86944 326986 87000
rect 327042 86944 327047 87000
rect 317524 86942 327047 86944
rect 317524 86940 317530 86942
rect 326981 86939 327047 86942
rect 336641 87002 336707 87005
rect 340462 87002 340522 87078
rect 356053 87075 356119 87078
rect 369902 87078 379346 87138
rect 336641 87000 340522 87002
rect 336641 86944 336646 87000
rect 336702 86944 340522 87000
rect 336641 86942 340522 86944
rect 336641 86939 336707 86942
rect 366950 86940 366956 87004
rect 367020 87002 367026 87004
rect 369902 87002 369962 87078
rect 367020 86942 369962 87002
rect 386278 87002 386338 87350
rect 425145 87274 425211 87277
rect 449249 87274 449315 87277
rect 453982 87274 453988 87276
rect 425145 87272 437490 87274
rect 425145 87216 425150 87272
rect 425206 87216 437490 87272
rect 425145 87214 437490 87216
rect 425145 87211 425211 87214
rect 398465 87138 398531 87141
rect 389222 87136 398531 87138
rect 389222 87080 398470 87136
rect 398526 87080 398531 87136
rect 389222 87078 398531 87080
rect 389222 87002 389282 87078
rect 398465 87075 398531 87078
rect 398833 87138 398899 87141
rect 417877 87138 417943 87141
rect 398833 87136 405658 87138
rect 398833 87080 398838 87136
rect 398894 87080 405658 87136
rect 398833 87078 405658 87080
rect 398833 87075 398899 87078
rect 386278 86942 389282 87002
rect 405598 87002 405658 87078
rect 408542 87136 417943 87138
rect 408542 87080 417882 87136
rect 417938 87080 417943 87136
rect 408542 87078 417943 87080
rect 408542 87002 408602 87078
rect 417877 87075 417943 87078
rect 418337 87138 418403 87141
rect 435173 87138 435239 87141
rect 418337 87136 424978 87138
rect 418337 87080 418342 87136
rect 418398 87080 424978 87136
rect 418337 87078 424978 87080
rect 418337 87075 418403 87078
rect 405598 86942 408602 87002
rect 424918 87002 424978 87078
rect 435173 87136 435282 87138
rect 435173 87080 435178 87136
rect 435234 87080 435282 87136
rect 435173 87075 435282 87080
rect 435222 87005 435282 87075
rect 425053 87002 425119 87005
rect 424918 87000 425119 87002
rect 424918 86944 425058 87000
rect 425114 86944 425119 87000
rect 424918 86942 425119 86944
rect 367020 86940 367026 86942
rect 425053 86939 425119 86942
rect 435173 87000 435282 87005
rect 435173 86944 435178 87000
rect 435234 86944 435282 87000
rect 435173 86942 435282 86944
rect 437430 87002 437490 87214
rect 449249 87272 453988 87274
rect 449249 87216 449254 87272
rect 449310 87216 453988 87272
rect 449249 87214 453988 87216
rect 449249 87211 449315 87214
rect 453982 87212 453988 87214
rect 454052 87212 454058 87276
rect 473302 87212 473308 87276
rect 473372 87274 473378 87276
rect 473372 87214 489930 87274
rect 473372 87212 473378 87214
rect 463601 87138 463667 87141
rect 489870 87138 489930 87214
rect 499622 87214 509250 87274
rect 463601 87136 463802 87138
rect 463601 87080 463606 87136
rect 463662 87080 463802 87136
rect 463601 87078 463802 87080
rect 489870 87078 499498 87138
rect 463601 87075 463667 87078
rect 463742 87005 463802 87078
rect 444373 87002 444439 87005
rect 437430 87000 444439 87002
rect 437430 86944 444378 87000
rect 444434 86944 444439 87000
rect 437430 86942 444439 86944
rect 463742 87000 463851 87005
rect 463742 86944 463790 87000
rect 463846 86944 463851 87000
rect 463742 86942 463851 86944
rect 435173 86939 435239 86942
rect 444373 86939 444439 86942
rect 463785 86939 463851 86942
rect 466545 87002 466611 87005
rect 473302 87002 473308 87004
rect 466545 87000 473308 87002
rect 466545 86944 466550 87000
rect 466606 86944 473308 87000
rect 466545 86942 473308 86944
rect 466545 86939 466611 86942
rect 473302 86940 473308 86942
rect 473372 86940 473378 87004
rect 499438 87002 499498 87078
rect 499622 87002 499682 87214
rect 509190 87138 509250 87214
rect 518942 87214 528570 87274
rect 509190 87078 518818 87138
rect 499438 86942 499682 87002
rect 518758 87002 518818 87078
rect 518942 87002 519002 87214
rect 528510 87138 528570 87214
rect 538262 87214 547890 87274
rect 528510 87078 538138 87138
rect 518758 86942 519002 87002
rect 538078 87002 538138 87078
rect 538262 87002 538322 87214
rect 547830 87138 547890 87214
rect 557582 87214 567210 87274
rect 547830 87078 557458 87138
rect 538078 86942 538322 87002
rect 557398 87002 557458 87078
rect 557582 87002 557642 87214
rect 567150 87138 567210 87214
rect 583342 87138 583402 87894
rect 583520 87804 584960 87894
rect 567150 87078 576778 87138
rect 557398 86942 557642 87002
rect 576718 87002 576778 87078
rect 576902 87078 583402 87138
rect 576902 87002 576962 87078
rect 576718 86942 576962 87002
rect 234797 85778 234863 85781
rect 234797 85776 234906 85778
rect 234797 85720 234802 85776
rect 234858 85720 234906 85776
rect 234797 85715 234906 85720
rect 234846 85645 234906 85715
rect 234797 85640 234906 85645
rect 234797 85584 234802 85640
rect 234858 85584 234906 85640
rect 234797 85582 234906 85584
rect 251173 85642 251239 85645
rect 251357 85642 251423 85645
rect 251173 85640 251423 85642
rect 251173 85584 251178 85640
rect 251234 85584 251362 85640
rect 251418 85584 251423 85640
rect 251173 85582 251423 85584
rect 234797 85579 234863 85582
rect 251173 85579 251239 85582
rect 251357 85579 251423 85582
rect -960 78978 480 79068
rect 2773 78978 2839 78981
rect -960 78976 2839 78978
rect -960 78920 2778 78976
rect 2834 78920 2839 78976
rect -960 78918 2839 78920
rect -960 78828 480 78918
rect 2773 78915 2839 78918
rect 580257 76258 580323 76261
rect 583520 76258 584960 76348
rect 580257 76256 584960 76258
rect 580257 76200 580262 76256
rect 580318 76200 584960 76256
rect 580257 76198 584960 76200
rect 580257 76195 580323 76198
rect 583520 76108 584960 76198
rect 287329 67690 287395 67693
rect 287286 67688 287395 67690
rect 287286 67632 287334 67688
rect 287390 67632 287395 67688
rect 287286 67627 287395 67632
rect 287286 67554 287346 67627
rect 287421 67554 287487 67557
rect 287286 67552 287487 67554
rect 287286 67496 287426 67552
rect 287482 67496 287487 67552
rect 287286 67494 287487 67496
rect 287421 67491 287487 67494
rect -960 64562 480 64652
rect 3417 64562 3483 64565
rect 583520 64562 584960 64652
rect -960 64560 3483 64562
rect -960 64504 3422 64560
rect 3478 64504 3483 64560
rect -960 64502 3483 64504
rect -960 64412 480 64502
rect 3417 64499 3483 64502
rect 583342 64502 584960 64562
rect 453982 64228 453988 64292
rect 454052 64290 454058 64292
rect 460841 64290 460907 64293
rect 454052 64288 460907 64290
rect 454052 64232 460846 64288
rect 460902 64232 460907 64288
rect 454052 64230 460907 64232
rect 454052 64228 454058 64230
rect 460841 64227 460907 64230
rect 343582 63956 343588 64020
rect 343652 64018 343658 64020
rect 348325 64018 348391 64021
rect 447225 64018 447291 64021
rect 453982 64018 453988 64020
rect 343652 64016 348391 64018
rect 343652 63960 348330 64016
rect 348386 63960 348391 64016
rect 343652 63958 348391 63960
rect 343652 63956 343658 63958
rect 348325 63955 348391 63958
rect 376710 63958 386338 64018
rect 272977 63882 273043 63885
rect 253798 63880 273043 63882
rect 253798 63824 272982 63880
rect 273038 63824 273043 63880
rect 253798 63822 273043 63824
rect 237230 63548 237236 63612
rect 237300 63610 237306 63612
rect 253798 63610 253858 63822
rect 272977 63819 273043 63822
rect 273161 63882 273227 63885
rect 335261 63882 335327 63885
rect 273161 63880 274466 63882
rect 273161 63824 273166 63880
rect 273222 63824 274466 63880
rect 273161 63822 274466 63824
rect 273161 63819 273227 63822
rect 274406 63746 274466 63822
rect 289678 63822 292682 63882
rect 289678 63746 289738 63822
rect 274406 63686 289738 63746
rect 292622 63746 292682 63822
rect 335261 63880 336842 63882
rect 335261 63824 335266 63880
rect 335322 63824 336842 63880
rect 335261 63822 336842 63824
rect 335261 63819 335327 63822
rect 326797 63746 326863 63749
rect 292622 63686 317522 63746
rect 237300 63550 253858 63610
rect 317462 63610 317522 63686
rect 325742 63744 326863 63746
rect 325742 63688 326802 63744
rect 326858 63688 326863 63744
rect 325742 63686 326863 63688
rect 336782 63746 336842 63822
rect 343582 63746 343588 63748
rect 336782 63686 343588 63746
rect 325742 63610 325802 63686
rect 326797 63683 326863 63686
rect 343582 63684 343588 63686
rect 343652 63684 343658 63748
rect 348325 63746 348391 63749
rect 359549 63746 359615 63749
rect 376710 63746 376770 63958
rect 348325 63744 359615 63746
rect 348325 63688 348330 63744
rect 348386 63688 359554 63744
rect 359610 63688 359615 63744
rect 348325 63686 359615 63688
rect 348325 63683 348391 63686
rect 359549 63683 359615 63686
rect 369902 63686 376770 63746
rect 317462 63550 325802 63610
rect 365621 63610 365687 63613
rect 369902 63610 369962 63686
rect 365621 63608 369962 63610
rect 365621 63552 365626 63608
rect 365682 63552 369962 63608
rect 365621 63550 369962 63552
rect 386278 63610 386338 63958
rect 447225 64016 453988 64018
rect 447225 63960 447230 64016
rect 447286 63960 453988 64016
rect 447225 63958 453988 63960
rect 447225 63955 447291 63958
rect 453982 63956 453988 63958
rect 454052 63956 454058 64020
rect 460841 63882 460907 63885
rect 460841 63880 470610 63882
rect 460841 63824 460846 63880
rect 460902 63824 470610 63880
rect 460841 63822 470610 63824
rect 460841 63819 460907 63822
rect 398465 63746 398531 63749
rect 389222 63744 398531 63746
rect 389222 63688 398470 63744
rect 398526 63688 398531 63744
rect 389222 63686 398531 63688
rect 389222 63610 389282 63686
rect 398465 63683 398531 63686
rect 399017 63746 399083 63749
rect 417877 63746 417943 63749
rect 399017 63744 405658 63746
rect 399017 63688 399022 63744
rect 399078 63688 405658 63744
rect 399017 63686 405658 63688
rect 399017 63683 399083 63686
rect 386278 63550 389282 63610
rect 405598 63610 405658 63686
rect 408542 63744 417943 63746
rect 408542 63688 417882 63744
rect 417938 63688 417943 63744
rect 408542 63686 417943 63688
rect 408542 63610 408602 63686
rect 417877 63683 417943 63686
rect 419625 63746 419691 63749
rect 447133 63746 447199 63749
rect 419625 63744 424978 63746
rect 419625 63688 419630 63744
rect 419686 63688 424978 63744
rect 419625 63686 424978 63688
rect 419625 63683 419691 63686
rect 405598 63550 408602 63610
rect 424918 63610 424978 63686
rect 427862 63744 447199 63746
rect 427862 63688 447138 63744
rect 447194 63688 447199 63744
rect 427862 63686 447199 63688
rect 470550 63746 470610 63822
rect 480302 63822 489930 63882
rect 470550 63686 480178 63746
rect 427862 63610 427922 63686
rect 447133 63683 447199 63686
rect 424918 63550 427922 63610
rect 480118 63610 480178 63686
rect 480302 63610 480362 63822
rect 489870 63746 489930 63822
rect 499622 63822 509250 63882
rect 489870 63686 499498 63746
rect 480118 63550 480362 63610
rect 499438 63610 499498 63686
rect 499622 63610 499682 63822
rect 509190 63746 509250 63822
rect 518942 63822 528570 63882
rect 509190 63686 518818 63746
rect 499438 63550 499682 63610
rect 518758 63610 518818 63686
rect 518942 63610 519002 63822
rect 528510 63746 528570 63822
rect 538262 63822 547890 63882
rect 528510 63686 538138 63746
rect 518758 63550 519002 63610
rect 538078 63610 538138 63686
rect 538262 63610 538322 63822
rect 547830 63746 547890 63822
rect 557582 63822 567210 63882
rect 547830 63686 557458 63746
rect 538078 63550 538322 63610
rect 557398 63610 557458 63686
rect 557582 63610 557642 63822
rect 567150 63746 567210 63822
rect 583342 63746 583402 64502
rect 583520 64412 584960 64502
rect 567150 63686 576778 63746
rect 557398 63550 557642 63610
rect 576718 63610 576778 63686
rect 576902 63686 583402 63746
rect 576902 63610 576962 63686
rect 576718 63550 576962 63610
rect 237300 63548 237306 63550
rect 365621 63547 365687 63550
rect 251449 56810 251515 56813
rect 251406 56808 251515 56810
rect 251406 56752 251454 56808
rect 251510 56752 251515 56808
rect 251406 56747 251515 56752
rect 251406 56541 251466 56747
rect 251406 56536 251515 56541
rect 251406 56480 251454 56536
rect 251510 56480 251515 56536
rect 251406 56478 251515 56480
rect 251449 56475 251515 56478
rect 583520 52716 584960 52956
rect -960 50146 480 50236
rect 4061 50146 4127 50149
rect -960 50144 4127 50146
rect -960 50088 4066 50144
rect 4122 50088 4127 50144
rect -960 50086 4127 50088
rect -960 49996 480 50086
rect 4061 50083 4127 50086
rect 336917 48242 336983 48245
rect 336782 48240 336983 48242
rect 336782 48184 336922 48240
rect 336978 48184 336983 48240
rect 336782 48182 336983 48184
rect 336782 48106 336842 48182
rect 336917 48179 336983 48182
rect 434253 48244 434319 48245
rect 434253 48240 434300 48244
rect 434364 48242 434370 48244
rect 434253 48184 434258 48240
rect 434253 48180 434300 48184
rect 434364 48182 434410 48242
rect 434364 48180 434370 48182
rect 434253 48179 434319 48180
rect 337009 48106 337075 48109
rect 336782 48104 337075 48106
rect 336782 48048 337014 48104
rect 337070 48048 337075 48104
rect 336782 48046 337075 48048
rect 337009 48043 337075 48046
rect 347957 45522 348023 45525
rect 347822 45520 348023 45522
rect 347822 45464 347962 45520
rect 348018 45464 348023 45520
rect 347822 45462 348023 45464
rect 347822 45386 347882 45462
rect 347957 45459 348023 45462
rect 348049 45386 348115 45389
rect 347822 45384 348115 45386
rect 347822 45328 348054 45384
rect 348110 45328 348115 45384
rect 347822 45326 348115 45328
rect 348049 45323 348115 45326
rect 307937 44162 308003 44165
rect 308213 44162 308279 44165
rect 307937 44160 308279 44162
rect 307937 44104 307942 44160
rect 307998 44104 308218 44160
rect 308274 44104 308279 44160
rect 307937 44102 308279 44104
rect 307937 44099 308003 44102
rect 308213 44099 308279 44102
rect 434294 41244 434300 41308
rect 434364 41306 434370 41308
rect 434437 41306 434503 41309
rect 434364 41304 434503 41306
rect 434364 41248 434442 41304
rect 434498 41248 434503 41304
rect 434364 41246 434503 41248
rect 434364 41244 434370 41246
rect 434437 41243 434503 41246
rect 583520 41034 584960 41124
rect 583342 40974 584960 41034
rect 453982 40700 453988 40764
rect 454052 40762 454058 40764
rect 460841 40762 460907 40765
rect 454052 40760 460907 40762
rect 454052 40704 460846 40760
rect 460902 40704 460907 40760
rect 454052 40702 460907 40704
rect 454052 40700 454058 40702
rect 460841 40699 460907 40702
rect 328361 40626 328427 40629
rect 337929 40626 337995 40629
rect 328361 40624 337995 40626
rect 328361 40568 328366 40624
rect 328422 40568 337934 40624
rect 337990 40568 337995 40624
rect 328361 40566 337995 40568
rect 328361 40563 328427 40566
rect 337929 40563 337995 40566
rect 447225 40490 447291 40493
rect 453982 40490 453988 40492
rect 376710 40430 386338 40490
rect 249742 40292 249748 40356
rect 249812 40354 249818 40356
rect 270493 40354 270559 40357
rect 249812 40352 270559 40354
rect 249812 40296 270498 40352
rect 270554 40296 270559 40352
rect 249812 40294 270559 40296
rect 249812 40292 249818 40294
rect 270493 40291 270559 40294
rect 280521 40354 280587 40357
rect 297541 40354 297607 40357
rect 280521 40352 289738 40354
rect 280521 40296 280526 40352
rect 280582 40296 289738 40352
rect 280521 40294 289738 40296
rect 280521 40291 280587 40294
rect 289678 40218 289738 40294
rect 289862 40352 297607 40354
rect 289862 40296 297546 40352
rect 297602 40296 297607 40352
rect 289862 40294 297607 40296
rect 289862 40218 289922 40294
rect 297541 40291 297607 40294
rect 328361 40218 328427 40221
rect 356053 40218 356119 40221
rect 376710 40218 376770 40430
rect 289678 40158 289922 40218
rect 312494 40216 328427 40218
rect 312494 40160 328366 40216
rect 328422 40160 328427 40216
rect 312494 40158 328427 40160
rect 232998 40020 233004 40084
rect 233068 40082 233074 40084
rect 249742 40082 249748 40084
rect 233068 40022 249748 40082
rect 233068 40020 233074 40022
rect 249742 40020 249748 40022
rect 249812 40020 249818 40084
rect 297541 40082 297607 40085
rect 312494 40082 312554 40158
rect 328361 40155 328427 40158
rect 350582 40216 356119 40218
rect 350582 40160 356058 40216
rect 356114 40160 356119 40216
rect 350582 40158 356119 40160
rect 297541 40080 312554 40082
rect 297541 40024 297546 40080
rect 297602 40024 312554 40080
rect 297541 40022 312554 40024
rect 337929 40082 337995 40085
rect 350582 40082 350642 40158
rect 356053 40155 356119 40158
rect 369902 40158 376770 40218
rect 337929 40080 350642 40082
rect 337929 40024 337934 40080
rect 337990 40024 350642 40080
rect 337929 40022 350642 40024
rect 365621 40082 365687 40085
rect 369902 40082 369962 40158
rect 365621 40080 369962 40082
rect 365621 40024 365626 40080
rect 365682 40024 369962 40080
rect 365621 40022 369962 40024
rect 386278 40082 386338 40430
rect 447225 40488 453988 40490
rect 447225 40432 447230 40488
rect 447286 40432 453988 40488
rect 447225 40430 453988 40432
rect 447225 40427 447291 40430
rect 453982 40428 453988 40430
rect 454052 40428 454058 40492
rect 460841 40354 460907 40357
rect 460841 40352 470610 40354
rect 460841 40296 460846 40352
rect 460902 40296 470610 40352
rect 460841 40294 470610 40296
rect 460841 40291 460907 40294
rect 398465 40218 398531 40221
rect 389222 40216 398531 40218
rect 389222 40160 398470 40216
rect 398526 40160 398531 40216
rect 389222 40158 398531 40160
rect 389222 40082 389282 40158
rect 398465 40155 398531 40158
rect 399017 40218 399083 40221
rect 417877 40218 417943 40221
rect 399017 40216 405658 40218
rect 399017 40160 399022 40216
rect 399078 40160 405658 40216
rect 399017 40158 405658 40160
rect 399017 40155 399083 40158
rect 386278 40022 389282 40082
rect 405598 40082 405658 40158
rect 408542 40216 417943 40218
rect 408542 40160 417882 40216
rect 417938 40160 417943 40216
rect 408542 40158 417943 40160
rect 408542 40082 408602 40158
rect 417877 40155 417943 40158
rect 418337 40218 418403 40221
rect 447133 40218 447199 40221
rect 418337 40216 424978 40218
rect 418337 40160 418342 40216
rect 418398 40160 424978 40216
rect 418337 40158 424978 40160
rect 418337 40155 418403 40158
rect 405598 40022 408602 40082
rect 424918 40082 424978 40158
rect 427862 40216 447199 40218
rect 427862 40160 447138 40216
rect 447194 40160 447199 40216
rect 427862 40158 447199 40160
rect 470550 40218 470610 40294
rect 480302 40294 489930 40354
rect 470550 40158 480178 40218
rect 427862 40082 427922 40158
rect 447133 40155 447199 40158
rect 424918 40022 427922 40082
rect 480118 40082 480178 40158
rect 480302 40082 480362 40294
rect 489870 40218 489930 40294
rect 499622 40294 509250 40354
rect 489870 40158 499498 40218
rect 480118 40022 480362 40082
rect 499438 40082 499498 40158
rect 499622 40082 499682 40294
rect 509190 40218 509250 40294
rect 518942 40294 528570 40354
rect 509190 40158 518818 40218
rect 499438 40022 499682 40082
rect 518758 40082 518818 40158
rect 518942 40082 519002 40294
rect 528510 40218 528570 40294
rect 538262 40294 547890 40354
rect 528510 40158 538138 40218
rect 518758 40022 519002 40082
rect 538078 40082 538138 40158
rect 538262 40082 538322 40294
rect 547830 40218 547890 40294
rect 557582 40294 567210 40354
rect 547830 40158 557458 40218
rect 538078 40022 538322 40082
rect 557398 40082 557458 40158
rect 557582 40082 557642 40294
rect 567150 40218 567210 40294
rect 583342 40218 583402 40974
rect 583520 40884 584960 40974
rect 567150 40158 576778 40218
rect 557398 40022 557642 40082
rect 576718 40082 576778 40158
rect 576902 40158 583402 40218
rect 576902 40082 576962 40158
rect 576718 40022 576962 40082
rect 297541 40019 297607 40022
rect 337929 40019 337995 40022
rect 365621 40019 365687 40022
rect 299749 36002 299815 36005
rect 299933 36002 299999 36005
rect 299749 36000 299999 36002
rect -960 35866 480 35956
rect 299749 35944 299754 36000
rect 299810 35944 299938 36000
rect 299994 35944 299999 36000
rect 299749 35942 299999 35944
rect 299749 35939 299815 35942
rect 299933 35939 299999 35942
rect 444414 35866 444420 35868
rect -960 35806 444420 35866
rect -960 35716 480 35806
rect 444414 35804 444420 35806
rect 444484 35804 444490 35868
rect 234470 32540 234476 32604
rect 234540 32602 234546 32604
rect 238661 32602 238727 32605
rect 234540 32600 238727 32602
rect 234540 32544 238666 32600
rect 238722 32544 238727 32600
rect 234540 32542 238727 32544
rect 234540 32540 234546 32542
rect 238661 32539 238727 32542
rect 291837 29610 291903 29613
rect 291837 29608 296730 29610
rect 291837 29552 291842 29608
rect 291898 29552 296730 29608
rect 291837 29550 296730 29552
rect 291837 29547 291903 29550
rect 296670 29474 296730 29550
rect 315982 29548 315988 29612
rect 316052 29610 316058 29612
rect 325601 29610 325667 29613
rect 316052 29608 325667 29610
rect 316052 29552 325606 29608
rect 325662 29552 325667 29608
rect 316052 29550 325667 29552
rect 316052 29548 316058 29550
rect 325601 29547 325667 29550
rect 306281 29474 306347 29477
rect 249750 29414 263794 29474
rect 296670 29472 306347 29474
rect 296670 29416 306286 29472
rect 306342 29416 306347 29472
rect 296670 29414 306347 29416
rect 249750 29341 249810 29414
rect 249701 29338 249810 29341
rect 249620 29336 249810 29338
rect 249620 29280 249706 29336
rect 249762 29280 249810 29336
rect 249620 29278 249810 29280
rect 249701 29275 249767 29278
rect 238661 29202 238727 29205
rect 263734 29202 263794 29414
rect 306281 29411 306347 29414
rect 350582 29414 360026 29474
rect 273989 29338 274055 29341
rect 284937 29338 285003 29341
rect 273989 29336 285003 29338
rect 273989 29280 273994 29336
rect 274050 29280 284942 29336
rect 284998 29280 285003 29336
rect 273989 29278 285003 29280
rect 273989 29275 274055 29278
rect 284937 29275 285003 29278
rect 325601 29338 325667 29341
rect 325601 29336 327090 29338
rect 325601 29280 325606 29336
rect 325662 29280 327090 29336
rect 325601 29278 327090 29280
rect 325601 29275 325667 29278
rect 270493 29202 270559 29205
rect 238661 29200 240242 29202
rect 238661 29144 238666 29200
rect 238722 29144 240242 29200
rect 238661 29142 240242 29144
rect 263734 29200 270559 29202
rect 263734 29144 270498 29200
rect 270554 29144 270559 29200
rect 263734 29142 270559 29144
rect 238661 29139 238727 29142
rect 240182 28930 240242 29142
rect 270493 29139 270559 29142
rect 306281 29202 306347 29205
rect 315941 29204 316007 29205
rect 327030 29204 327090 29278
rect 306281 29200 306482 29202
rect 306281 29144 306286 29200
rect 306342 29144 306482 29200
rect 306281 29142 306482 29144
rect 306281 29139 306347 29142
rect 284937 29066 285003 29069
rect 291837 29066 291903 29069
rect 284937 29064 291903 29066
rect 284937 29008 284942 29064
rect 284998 29008 291842 29064
rect 291898 29008 291903 29064
rect 284937 29006 291903 29008
rect 306422 29066 306482 29142
rect 315941 29200 315988 29204
rect 316052 29202 316058 29204
rect 315941 29144 315946 29200
rect 315941 29140 315988 29144
rect 316052 29142 316134 29202
rect 316052 29140 316058 29142
rect 327022 29140 327028 29204
rect 327092 29140 327098 29204
rect 327206 29140 327212 29204
rect 327276 29202 327282 29204
rect 350582 29202 350642 29414
rect 327276 29142 350642 29202
rect 359966 29202 360026 29414
rect 376710 29414 386338 29474
rect 366950 29338 366956 29340
rect 360334 29278 366956 29338
rect 360334 29202 360394 29278
rect 366950 29276 366956 29278
rect 367020 29276 367026 29340
rect 376710 29202 376770 29414
rect 359966 29142 360394 29202
rect 369902 29142 376770 29202
rect 327276 29140 327282 29142
rect 315941 29139 316007 29140
rect 315941 29066 316007 29069
rect 306422 29064 316007 29066
rect 306422 29008 315946 29064
rect 316002 29008 316007 29064
rect 306422 29006 316007 29008
rect 284937 29003 285003 29006
rect 291837 29003 291903 29006
rect 315941 29003 316007 29006
rect 366950 29004 366956 29068
rect 367020 29066 367026 29068
rect 369902 29066 369962 29142
rect 367020 29006 369962 29066
rect 386278 29066 386338 29414
rect 462262 29412 462268 29476
rect 462332 29474 462338 29476
rect 471881 29474 471947 29477
rect 462332 29472 471947 29474
rect 462332 29416 471886 29472
rect 471942 29416 471947 29472
rect 462332 29414 471947 29416
rect 462332 29412 462338 29414
rect 471881 29411 471947 29414
rect 449249 29338 449315 29341
rect 482921 29338 482987 29341
rect 583520 29338 584960 29428
rect 427678 29278 437490 29338
rect 398465 29202 398531 29205
rect 389222 29200 398531 29202
rect 389222 29144 398470 29200
rect 398526 29144 398531 29200
rect 389222 29142 398531 29144
rect 389222 29066 389282 29142
rect 398465 29139 398531 29142
rect 399017 29202 399083 29205
rect 417877 29202 417943 29205
rect 399017 29200 405658 29202
rect 399017 29144 399022 29200
rect 399078 29144 405658 29200
rect 399017 29142 405658 29144
rect 399017 29139 399083 29142
rect 386278 29006 389282 29066
rect 405598 29066 405658 29142
rect 408542 29200 417943 29202
rect 408542 29144 417882 29200
rect 417938 29144 417943 29200
rect 408542 29142 417943 29144
rect 408542 29066 408602 29142
rect 417877 29139 417943 29142
rect 418153 29202 418219 29205
rect 418153 29200 424978 29202
rect 418153 29144 418158 29200
rect 418214 29144 424978 29200
rect 418153 29142 424978 29144
rect 418153 29139 418219 29142
rect 405598 29006 408602 29066
rect 424918 29066 424978 29142
rect 427678 29066 427738 29278
rect 424918 29006 427738 29066
rect 437430 29066 437490 29278
rect 449249 29336 458834 29338
rect 449249 29280 449254 29336
rect 449310 29280 458834 29336
rect 449249 29278 458834 29280
rect 449249 29275 449315 29278
rect 458774 29202 458834 29278
rect 482921 29336 489930 29338
rect 482921 29280 482926 29336
rect 482982 29280 489930 29336
rect 482921 29278 489930 29280
rect 482921 29275 482987 29278
rect 462262 29202 462268 29204
rect 458774 29142 462268 29202
rect 462262 29140 462268 29142
rect 462332 29140 462338 29204
rect 476021 29202 476087 29205
rect 473310 29200 476087 29202
rect 473310 29144 476026 29200
rect 476082 29144 476087 29200
rect 473310 29142 476087 29144
rect 489870 29202 489930 29278
rect 499622 29278 509250 29338
rect 489870 29142 499498 29202
rect 444373 29066 444439 29069
rect 437430 29064 444439 29066
rect 437430 29008 444378 29064
rect 444434 29008 444439 29064
rect 437430 29006 444439 29008
rect 367020 29004 367026 29006
rect 444373 29003 444439 29006
rect 471881 29066 471947 29069
rect 473310 29066 473370 29142
rect 476021 29139 476087 29142
rect 471881 29064 473370 29066
rect 471881 29008 471886 29064
rect 471942 29008 473370 29064
rect 471881 29006 473370 29008
rect 499438 29066 499498 29142
rect 499622 29066 499682 29278
rect 509190 29202 509250 29278
rect 518942 29278 528570 29338
rect 509190 29142 518818 29202
rect 499438 29006 499682 29066
rect 518758 29066 518818 29142
rect 518942 29066 519002 29278
rect 528510 29202 528570 29278
rect 538262 29278 547890 29338
rect 528510 29142 538138 29202
rect 518758 29006 519002 29066
rect 538078 29066 538138 29142
rect 538262 29066 538322 29278
rect 547830 29202 547890 29278
rect 557582 29278 567210 29338
rect 547830 29142 557458 29202
rect 538078 29006 538322 29066
rect 557398 29066 557458 29142
rect 557582 29066 557642 29278
rect 567150 29202 567210 29278
rect 583342 29278 584960 29338
rect 583342 29202 583402 29278
rect 567150 29142 576778 29202
rect 557398 29006 557642 29066
rect 576718 29066 576778 29142
rect 576902 29142 583402 29202
rect 583520 29188 584960 29278
rect 576902 29066 576962 29142
rect 576718 29006 576962 29066
rect 471881 29003 471947 29006
rect 249701 28930 249767 28933
rect 287237 28930 287303 28933
rect 240182 28928 249767 28930
rect 240182 28872 249706 28928
rect 249762 28872 249767 28928
rect 240182 28870 249767 28872
rect 249701 28867 249767 28870
rect 287102 28928 287303 28930
rect 287102 28872 287242 28928
rect 287298 28872 287303 28928
rect 287102 28870 287303 28872
rect 287102 28794 287162 28870
rect 287237 28867 287303 28870
rect 287329 28794 287395 28797
rect 287102 28792 287395 28794
rect 287102 28736 287334 28792
rect 287390 28736 287395 28792
rect 287102 28734 287395 28736
rect 287329 28731 287395 28734
rect 348049 26210 348115 26213
rect 348233 26210 348299 26213
rect 348049 26208 348299 26210
rect 348049 26152 348054 26208
rect 348110 26152 348238 26208
rect 348294 26152 348299 26208
rect 348049 26150 348299 26152
rect 348049 26147 348115 26150
rect 348233 26147 348299 26150
rect 348049 24850 348115 24853
rect 348233 24850 348299 24853
rect 348049 24848 348299 24850
rect 348049 24792 348054 24848
rect 348110 24792 348238 24848
rect 348294 24792 348299 24848
rect 348049 24790 348299 24792
rect 348049 24787 348115 24790
rect 348233 24787 348299 24790
rect 229369 22268 229435 22269
rect 229318 22266 229324 22268
rect 229278 22206 229324 22266
rect 229388 22264 229435 22268
rect 229430 22208 229435 22264
rect 229318 22204 229324 22206
rect 229388 22204 229435 22208
rect 229369 22203 229435 22204
rect 448462 21994 448468 21996
rect 614 21934 448468 21994
rect -960 21450 480 21540
rect 614 21450 674 21934
rect 448462 21932 448468 21934
rect 448532 21932 448538 21996
rect -960 21390 674 21450
rect -960 21300 480 21390
rect 266997 19274 267063 19277
rect 266862 19272 267063 19274
rect 266862 19216 267002 19272
rect 267058 19216 267063 19272
rect 266862 19214 267063 19216
rect 266862 19138 266922 19214
rect 266997 19211 267063 19214
rect 267273 19138 267339 19141
rect 266862 19136 267339 19138
rect 266862 19080 267278 19136
rect 267334 19080 267339 19136
rect 266862 19078 267339 19080
rect 267273 19075 267339 19078
rect 240409 18186 240475 18189
rect 241789 18186 241855 18189
rect 240182 18184 240475 18186
rect 240182 18128 240414 18184
rect 240470 18128 240475 18184
rect 240182 18126 240475 18128
rect 229369 18052 229435 18053
rect 229318 17988 229324 18052
rect 229388 18050 229435 18052
rect 240182 18050 240242 18126
rect 240409 18123 240475 18126
rect 241608 18184 241855 18186
rect 241608 18128 241794 18184
rect 241850 18128 241855 18184
rect 241608 18126 241855 18128
rect 241608 18053 241668 18126
rect 241789 18123 241855 18126
rect 240317 18050 240383 18053
rect 229388 18048 229480 18050
rect 229430 17992 229480 18048
rect 229388 17990 229480 17992
rect 240182 18048 240383 18050
rect 240182 17992 240322 18048
rect 240378 17992 240383 18048
rect 240182 17990 240383 17992
rect 229388 17988 229435 17990
rect 229369 17987 229435 17988
rect 240317 17987 240383 17990
rect 241605 18048 241671 18053
rect 241605 17992 241610 18048
rect 241666 17992 241671 18048
rect 241605 17987 241671 17992
rect 583520 17642 584960 17732
rect 583342 17582 584960 17642
rect 376710 17038 386338 17098
rect 360009 16826 360075 16829
rect 350582 16824 360075 16826
rect 350582 16768 360014 16824
rect 360070 16768 360075 16824
rect 350582 16766 360075 16768
rect 231710 16628 231716 16692
rect 231780 16690 231786 16692
rect 350582 16690 350642 16766
rect 360009 16763 360075 16766
rect 361113 16826 361179 16829
rect 376710 16826 376770 17038
rect 361113 16824 367018 16826
rect 361113 16768 361118 16824
rect 361174 16768 367018 16824
rect 361113 16766 367018 16768
rect 361113 16763 361179 16766
rect 231780 16630 350642 16690
rect 366958 16690 367018 16766
rect 369902 16766 376770 16826
rect 369902 16690 369962 16766
rect 366958 16630 369962 16690
rect 386278 16690 386338 17038
rect 462262 17036 462268 17100
rect 462332 17098 462338 17100
rect 471881 17098 471947 17101
rect 462332 17096 471947 17098
rect 462332 17040 471886 17096
rect 471942 17040 471947 17096
rect 462332 17038 471947 17040
rect 462332 17036 462338 17038
rect 471881 17035 471947 17038
rect 434621 16962 434687 16965
rect 447225 16962 447291 16965
rect 482921 16962 482987 16965
rect 434621 16960 437490 16962
rect 434621 16904 434626 16960
rect 434682 16904 437490 16960
rect 434621 16902 437490 16904
rect 434621 16899 434687 16902
rect 398465 16826 398531 16829
rect 389222 16824 398531 16826
rect 389222 16768 398470 16824
rect 398526 16768 398531 16824
rect 389222 16766 398531 16768
rect 389222 16690 389282 16766
rect 398465 16763 398531 16766
rect 399017 16826 399083 16829
rect 417877 16826 417943 16829
rect 399017 16824 405658 16826
rect 399017 16768 399022 16824
rect 399078 16768 405658 16824
rect 399017 16766 405658 16768
rect 399017 16763 399083 16766
rect 386278 16630 389282 16690
rect 405598 16690 405658 16766
rect 408542 16824 417943 16826
rect 408542 16768 417882 16824
rect 417938 16768 417943 16824
rect 408542 16766 417943 16768
rect 408542 16690 408602 16766
rect 417877 16763 417943 16766
rect 425053 16690 425119 16693
rect 405598 16630 408602 16690
rect 424918 16688 425119 16690
rect 424918 16632 425058 16688
rect 425114 16632 425119 16688
rect 424918 16630 425119 16632
rect 437430 16690 437490 16902
rect 447225 16960 458834 16962
rect 447225 16904 447230 16960
rect 447286 16904 458834 16960
rect 447225 16902 458834 16904
rect 447225 16899 447291 16902
rect 458774 16826 458834 16902
rect 482921 16960 489930 16962
rect 482921 16904 482926 16960
rect 482982 16904 489930 16960
rect 482921 16902 489930 16904
rect 482921 16899 482987 16902
rect 462262 16826 462268 16828
rect 458774 16766 462268 16826
rect 462262 16764 462268 16766
rect 462332 16764 462338 16828
rect 476021 16826 476087 16829
rect 473310 16824 476087 16826
rect 473310 16768 476026 16824
rect 476082 16768 476087 16824
rect 473310 16766 476087 16768
rect 489870 16826 489930 16902
rect 499622 16902 509250 16962
rect 489870 16766 499498 16826
rect 444373 16690 444439 16693
rect 437430 16688 444439 16690
rect 437430 16632 444378 16688
rect 444434 16632 444439 16688
rect 437430 16630 444439 16632
rect 231780 16628 231786 16630
rect 417877 16418 417943 16421
rect 424918 16418 424978 16630
rect 425053 16627 425119 16630
rect 444373 16627 444439 16630
rect 471881 16690 471947 16693
rect 473310 16690 473370 16766
rect 476021 16763 476087 16766
rect 471881 16688 473370 16690
rect 471881 16632 471886 16688
rect 471942 16632 473370 16688
rect 471881 16630 473370 16632
rect 499438 16690 499498 16766
rect 499622 16690 499682 16902
rect 509190 16826 509250 16902
rect 518942 16902 528570 16962
rect 509190 16766 518818 16826
rect 499438 16630 499682 16690
rect 518758 16690 518818 16766
rect 518942 16690 519002 16902
rect 528510 16826 528570 16902
rect 538262 16902 547890 16962
rect 528510 16766 538138 16826
rect 518758 16630 519002 16690
rect 538078 16690 538138 16766
rect 538262 16690 538322 16902
rect 547830 16826 547890 16902
rect 557582 16902 567210 16962
rect 547830 16766 557458 16826
rect 538078 16630 538322 16690
rect 557398 16690 557458 16766
rect 557582 16690 557642 16902
rect 567150 16826 567210 16902
rect 583342 16826 583402 17582
rect 583520 17492 584960 17582
rect 567150 16766 576778 16826
rect 557398 16630 557642 16690
rect 576718 16690 576778 16766
rect 576902 16766 583402 16826
rect 576902 16690 576962 16766
rect 576718 16630 576962 16690
rect 471881 16627 471947 16630
rect 417877 16416 424978 16418
rect 417877 16360 417882 16416
rect 417938 16360 424978 16416
rect 417877 16358 424978 16360
rect 417877 16355 417943 16358
rect 305177 15194 305243 15197
rect 305361 15194 305427 15197
rect 305177 15192 305427 15194
rect 305177 15136 305182 15192
rect 305238 15136 305366 15192
rect 305422 15136 305427 15192
rect 305177 15134 305427 15136
rect 305177 15131 305243 15134
rect 305361 15131 305427 15134
rect 132585 8938 132651 8941
rect 278957 8938 279023 8941
rect 132585 8936 279023 8938
rect 132585 8880 132590 8936
rect 132646 8880 278962 8936
rect 279018 8880 279023 8936
rect 132585 8878 279023 8880
rect 132585 8875 132651 8878
rect 278957 8875 279023 8878
rect 251357 8394 251423 8397
rect 251541 8394 251607 8397
rect 251357 8392 251607 8394
rect 251357 8336 251362 8392
rect 251418 8336 251546 8392
rect 251602 8336 251607 8392
rect 251357 8334 251607 8336
rect 251357 8331 251423 8334
rect 251541 8331 251607 8334
rect 4061 8258 4127 8261
rect 445702 8258 445708 8260
rect 4061 8256 445708 8258
rect 4061 8200 4066 8256
rect 4122 8200 445708 8256
rect 4061 8198 445708 8200
rect 4061 8195 4127 8198
rect 445702 8196 445708 8198
rect 445772 8196 445778 8260
rect 3969 7578 4035 7581
rect 230565 7578 230631 7581
rect 3969 7576 230631 7578
rect 3969 7520 3974 7576
rect 4030 7520 230570 7576
rect 230626 7520 230631 7576
rect 3969 7518 230631 7520
rect 3969 7515 4035 7518
rect 230565 7515 230631 7518
rect -960 7170 480 7260
rect 4061 7170 4127 7173
rect -960 7168 4127 7170
rect -960 7112 4066 7168
rect 4122 7112 4127 7168
rect -960 7110 4127 7112
rect -960 7020 480 7110
rect 4061 7107 4127 7110
rect 55213 6218 55279 6221
rect 249977 6218 250043 6221
rect 55213 6216 250043 6218
rect 55213 6160 55218 6216
rect 55274 6160 249982 6216
rect 250038 6160 250043 6216
rect 55213 6158 250043 6160
rect 55213 6155 55279 6158
rect 249977 6155 250043 6158
rect 583520 5796 584960 6036
rect 205081 4858 205147 4861
rect 306373 4858 306439 4861
rect 205081 4856 306439 4858
rect 205081 4800 205086 4856
rect 205142 4800 306378 4856
rect 306434 4800 306439 4856
rect 205081 4798 306439 4800
rect 205081 4795 205147 4798
rect 306373 4795 306439 4798
rect 449801 4858 449867 4861
rect 579797 4858 579863 4861
rect 449801 4856 579863 4858
rect 449801 4800 449806 4856
rect 449862 4800 579802 4856
rect 579858 4800 579863 4856
rect 449801 4798 579863 4800
rect 449801 4795 449867 4798
rect 579797 4795 579863 4798
rect 6453 3362 6519 3365
rect 232129 3362 232195 3365
rect 6453 3360 232195 3362
rect 6453 3304 6458 3360
rect 6514 3304 232134 3360
rect 232190 3304 232195 3360
rect 6453 3302 232195 3304
rect 6453 3299 6519 3302
rect 232129 3299 232195 3302
<< via3 >>
rect 357388 563076 357452 563140
rect 366956 563076 367020 563140
rect 237788 562940 237852 563004
rect 252508 562940 252572 563004
rect 253612 562940 253676 563004
rect 266308 562940 266372 563004
rect 275876 562940 275940 563004
rect 446260 562940 446324 563004
rect 236868 562804 236932 562868
rect 5212 562668 5276 562732
rect 125548 562668 125612 562732
rect 135116 562668 135180 562732
rect 164188 562668 164252 562732
rect 167316 562668 167380 562732
rect 183508 562668 183572 562732
rect 193076 562668 193140 562732
rect 205036 562668 205100 562732
rect 207612 562668 207676 562732
rect 236500 562668 236564 562732
rect 424364 562668 424428 562732
rect 428412 562668 428476 562732
rect 436140 562668 436204 562732
rect 237972 562396 238036 562460
rect 288388 561580 288452 561644
rect 293172 561580 293236 561644
rect 50476 561308 50540 561372
rect 51580 561308 51644 561372
rect 85620 561308 85684 561372
rect 90220 561308 90284 561372
rect 108436 561308 108500 561372
rect 109724 561308 109788 561372
rect 117636 561308 117700 561372
rect 120764 561308 120828 561372
rect 135668 561308 135732 561372
rect 140084 561308 140148 561372
rect 147444 561308 147508 561372
rect 154436 561308 154500 561372
rect 154988 561308 155052 561372
rect 159404 561308 159468 561372
rect 176148 561308 176212 561372
rect 178724 561308 178788 561372
rect 193628 561308 193692 561372
rect 196756 561308 196820 561372
rect 223620 561308 223684 561372
rect 225460 561308 225524 561372
rect 325740 561308 325804 561372
rect 335124 561308 335188 561372
rect 393268 561308 393332 561372
rect 406332 561308 406396 561372
rect 335124 560900 335188 560964
rect 376708 560900 376772 560964
rect 280108 560764 280172 560828
rect 280108 560492 280172 560556
rect 357388 560824 357452 560828
rect 357388 560768 357402 560824
rect 357402 560768 357452 560824
rect 357388 560764 357452 560768
rect 308996 560492 309060 560556
rect 308996 560356 309060 560420
rect 335308 560628 335372 560692
rect 357388 560552 357452 560556
rect 357388 560496 357402 560552
rect 357402 560496 357452 560552
rect 357388 560492 357452 560496
rect 376708 560492 376772 560556
rect 447732 560220 447796 560284
rect 299428 559812 299492 559876
rect 299428 559540 299492 559604
rect 222148 559404 222212 559468
rect 231716 559268 231780 559332
rect 233004 559268 233068 559332
rect 234292 559268 234356 559332
rect 222148 559132 222212 559196
rect 236684 559404 236748 559468
rect 237236 559268 237300 559332
rect 238156 559328 238220 559332
rect 238156 559272 238206 559328
rect 238206 559272 238220 559328
rect 238156 559268 238220 559272
rect 252508 559132 252572 559196
rect 307708 559404 307772 559468
rect 299428 559268 299492 559332
rect 307892 559268 307956 559332
rect 383148 559328 383212 559332
rect 383148 559272 383198 559328
rect 383198 559272 383212 559328
rect 383148 559268 383212 559272
rect 384068 559404 384132 559468
rect 311940 559132 312004 559196
rect 244044 558996 244108 559060
rect 299428 558996 299492 559060
rect 311756 558996 311820 559060
rect 318748 558996 318812 559060
rect 244044 558724 244108 558788
rect 252508 558724 252572 558788
rect 318748 558724 318812 558788
rect 352052 559132 352116 559196
rect 338068 558996 338132 559060
rect 338068 558724 338132 558788
rect 351868 558996 351932 559060
rect 384068 559132 384132 559196
rect 409092 559404 409156 559468
rect 396028 559268 396092 559332
rect 396028 558996 396092 559060
rect 444420 559268 444484 559332
rect 445708 559268 445772 559332
rect 448468 559328 448532 559332
rect 448468 559272 448518 559328
rect 448518 559272 448532 559328
rect 448468 559268 448532 559272
rect 409092 558996 409156 559060
rect 383148 558180 383212 558244
rect 446260 486100 446324 486164
rect 236868 337996 236932 338060
rect 236684 309028 236748 309092
rect 434484 299372 434548 299436
rect 434484 289852 434548 289916
rect 434484 280060 434548 280124
rect 434484 270540 434548 270604
rect 434484 260748 434548 260812
rect 236500 252452 236564 252516
rect 434484 251228 434548 251292
rect 447732 204580 447796 204644
rect 357388 181460 357452 181524
rect 237788 181052 237852 181116
rect 241468 181052 241532 181116
rect 241468 180780 241532 180844
rect 299244 181188 299308 181252
rect 299428 181052 299492 181116
rect 357388 181188 357452 181252
rect 434300 173904 434364 173908
rect 434300 173848 434350 173904
rect 434350 173848 434364 173904
rect 434300 173844 434364 173848
rect 434300 164188 434364 164252
rect 327396 138272 327460 138276
rect 327396 138216 327446 138272
rect 327446 138216 327460 138272
rect 327396 138212 327460 138216
rect 327396 135280 327460 135284
rect 327396 135224 327410 135280
rect 327410 135224 327460 135280
rect 327396 135220 327460 135224
rect 453988 134540 454052 134604
rect 237972 133860 238036 133924
rect 453988 134268 454052 134332
rect 238156 91156 238220 91220
rect 299428 87484 299492 87548
rect 269068 87212 269132 87276
rect 299428 87212 299492 87276
rect 453988 87484 454052 87548
rect 366956 87348 367020 87412
rect 317460 87212 317524 87276
rect 269068 86940 269132 87004
rect 317460 86940 317524 87004
rect 366956 86940 367020 87004
rect 453988 87212 454052 87276
rect 473308 87212 473372 87276
rect 473308 86940 473372 87004
rect 453988 64228 454052 64292
rect 343588 63956 343652 64020
rect 237236 63548 237300 63612
rect 343588 63684 343652 63748
rect 453988 63956 454052 64020
rect 434300 48240 434364 48244
rect 434300 48184 434314 48240
rect 434314 48184 434364 48240
rect 434300 48180 434364 48184
rect 434300 41244 434364 41308
rect 453988 40700 454052 40764
rect 249748 40292 249812 40356
rect 233004 40020 233068 40084
rect 249748 40020 249812 40084
rect 453988 40428 454052 40492
rect 444420 35804 444484 35868
rect 234476 32540 234540 32604
rect 315988 29548 316052 29612
rect 315988 29200 316052 29204
rect 315988 29144 316002 29200
rect 316002 29144 316052 29200
rect 315988 29140 316052 29144
rect 327028 29140 327092 29204
rect 327212 29140 327276 29204
rect 366956 29276 367020 29340
rect 366956 29004 367020 29068
rect 462268 29412 462332 29476
rect 462268 29140 462332 29204
rect 229324 22264 229388 22268
rect 229324 22208 229374 22264
rect 229374 22208 229388 22264
rect 229324 22204 229388 22208
rect 448468 21932 448532 21996
rect 229324 18048 229388 18052
rect 229324 17992 229374 18048
rect 229374 17992 229388 18048
rect 229324 17988 229388 17992
rect 231716 16628 231780 16692
rect 462268 17036 462332 17100
rect 462268 16764 462332 16828
rect 445708 8196 445772 8260
<< metal4 >>
rect -8436 711278 -7836 711300
rect -8436 711042 -8254 711278
rect -8018 711042 -7836 711278
rect -8436 710958 -7836 711042
rect -8436 710722 -8254 710958
rect -8018 710722 -7836 710958
rect -8436 679254 -7836 710722
rect -8436 679018 -8254 679254
rect -8018 679018 -7836 679254
rect -8436 678934 -7836 679018
rect -8436 678698 -8254 678934
rect -8018 678698 -7836 678934
rect -8436 643254 -7836 678698
rect -8436 643018 -8254 643254
rect -8018 643018 -7836 643254
rect -8436 642934 -7836 643018
rect -8436 642698 -8254 642934
rect -8018 642698 -7836 642934
rect -8436 607254 -7836 642698
rect -8436 607018 -8254 607254
rect -8018 607018 -7836 607254
rect -8436 606934 -7836 607018
rect -8436 606698 -8254 606934
rect -8018 606698 -7836 606934
rect -8436 571254 -7836 606698
rect -8436 571018 -8254 571254
rect -8018 571018 -7836 571254
rect -8436 570934 -7836 571018
rect -8436 570698 -8254 570934
rect -8018 570698 -7836 570934
rect -8436 535254 -7836 570698
rect -8436 535018 -8254 535254
rect -8018 535018 -7836 535254
rect -8436 534934 -7836 535018
rect -8436 534698 -8254 534934
rect -8018 534698 -7836 534934
rect -8436 499254 -7836 534698
rect -8436 499018 -8254 499254
rect -8018 499018 -7836 499254
rect -8436 498934 -7836 499018
rect -8436 498698 -8254 498934
rect -8018 498698 -7836 498934
rect -8436 463254 -7836 498698
rect -8436 463018 -8254 463254
rect -8018 463018 -7836 463254
rect -8436 462934 -7836 463018
rect -8436 462698 -8254 462934
rect -8018 462698 -7836 462934
rect -8436 427254 -7836 462698
rect -8436 427018 -8254 427254
rect -8018 427018 -7836 427254
rect -8436 426934 -7836 427018
rect -8436 426698 -8254 426934
rect -8018 426698 -7836 426934
rect -8436 391254 -7836 426698
rect -8436 391018 -8254 391254
rect -8018 391018 -7836 391254
rect -8436 390934 -7836 391018
rect -8436 390698 -8254 390934
rect -8018 390698 -7836 390934
rect -8436 355254 -7836 390698
rect -8436 355018 -8254 355254
rect -8018 355018 -7836 355254
rect -8436 354934 -7836 355018
rect -8436 354698 -8254 354934
rect -8018 354698 -7836 354934
rect -8436 319254 -7836 354698
rect -8436 319018 -8254 319254
rect -8018 319018 -7836 319254
rect -8436 318934 -7836 319018
rect -8436 318698 -8254 318934
rect -8018 318698 -7836 318934
rect -8436 283254 -7836 318698
rect -8436 283018 -8254 283254
rect -8018 283018 -7836 283254
rect -8436 282934 -7836 283018
rect -8436 282698 -8254 282934
rect -8018 282698 -7836 282934
rect -8436 247254 -7836 282698
rect -8436 247018 -8254 247254
rect -8018 247018 -7836 247254
rect -8436 246934 -7836 247018
rect -8436 246698 -8254 246934
rect -8018 246698 -7836 246934
rect -8436 211254 -7836 246698
rect -8436 211018 -8254 211254
rect -8018 211018 -7836 211254
rect -8436 210934 -7836 211018
rect -8436 210698 -8254 210934
rect -8018 210698 -7836 210934
rect -8436 175254 -7836 210698
rect -8436 175018 -8254 175254
rect -8018 175018 -7836 175254
rect -8436 174934 -7836 175018
rect -8436 174698 -8254 174934
rect -8018 174698 -7836 174934
rect -8436 139254 -7836 174698
rect -8436 139018 -8254 139254
rect -8018 139018 -7836 139254
rect -8436 138934 -7836 139018
rect -8436 138698 -8254 138934
rect -8018 138698 -7836 138934
rect -8436 103254 -7836 138698
rect -8436 103018 -8254 103254
rect -8018 103018 -7836 103254
rect -8436 102934 -7836 103018
rect -8436 102698 -8254 102934
rect -8018 102698 -7836 102934
rect -8436 67254 -7836 102698
rect -8436 67018 -8254 67254
rect -8018 67018 -7836 67254
rect -8436 66934 -7836 67018
rect -8436 66698 -8254 66934
rect -8018 66698 -7836 66934
rect -8436 31254 -7836 66698
rect -8436 31018 -8254 31254
rect -8018 31018 -7836 31254
rect -8436 30934 -7836 31018
rect -8436 30698 -8254 30934
rect -8018 30698 -7836 30934
rect -8436 -6786 -7836 30698
rect -7516 710358 -6916 710380
rect -7516 710122 -7334 710358
rect -7098 710122 -6916 710358
rect -7516 710038 -6916 710122
rect -7516 709802 -7334 710038
rect -7098 709802 -6916 710038
rect -7516 697254 -6916 709802
rect 11604 710358 12204 711300
rect 11604 710122 11786 710358
rect 12022 710122 12204 710358
rect 11604 710038 12204 710122
rect 11604 709802 11786 710038
rect 12022 709802 12204 710038
rect -7516 697018 -7334 697254
rect -7098 697018 -6916 697254
rect -7516 696934 -6916 697018
rect -7516 696698 -7334 696934
rect -7098 696698 -6916 696934
rect -7516 661254 -6916 696698
rect -7516 661018 -7334 661254
rect -7098 661018 -6916 661254
rect -7516 660934 -6916 661018
rect -7516 660698 -7334 660934
rect -7098 660698 -6916 660934
rect -7516 625254 -6916 660698
rect -7516 625018 -7334 625254
rect -7098 625018 -6916 625254
rect -7516 624934 -6916 625018
rect -7516 624698 -7334 624934
rect -7098 624698 -6916 624934
rect -7516 589254 -6916 624698
rect -7516 589018 -7334 589254
rect -7098 589018 -6916 589254
rect -7516 588934 -6916 589018
rect -7516 588698 -7334 588934
rect -7098 588698 -6916 588934
rect -7516 553254 -6916 588698
rect -7516 553018 -7334 553254
rect -7098 553018 -6916 553254
rect -7516 552934 -6916 553018
rect -7516 552698 -7334 552934
rect -7098 552698 -6916 552934
rect -7516 517254 -6916 552698
rect -7516 517018 -7334 517254
rect -7098 517018 -6916 517254
rect -7516 516934 -6916 517018
rect -7516 516698 -7334 516934
rect -7098 516698 -6916 516934
rect -7516 481254 -6916 516698
rect -7516 481018 -7334 481254
rect -7098 481018 -6916 481254
rect -7516 480934 -6916 481018
rect -7516 480698 -7334 480934
rect -7098 480698 -6916 480934
rect -7516 445254 -6916 480698
rect -7516 445018 -7334 445254
rect -7098 445018 -6916 445254
rect -7516 444934 -6916 445018
rect -7516 444698 -7334 444934
rect -7098 444698 -6916 444934
rect -7516 409254 -6916 444698
rect -7516 409018 -7334 409254
rect -7098 409018 -6916 409254
rect -7516 408934 -6916 409018
rect -7516 408698 -7334 408934
rect -7098 408698 -6916 408934
rect -7516 373254 -6916 408698
rect -7516 373018 -7334 373254
rect -7098 373018 -6916 373254
rect -7516 372934 -6916 373018
rect -7516 372698 -7334 372934
rect -7098 372698 -6916 372934
rect -7516 337254 -6916 372698
rect -7516 337018 -7334 337254
rect -7098 337018 -6916 337254
rect -7516 336934 -6916 337018
rect -7516 336698 -7334 336934
rect -7098 336698 -6916 336934
rect -7516 301254 -6916 336698
rect -7516 301018 -7334 301254
rect -7098 301018 -6916 301254
rect -7516 300934 -6916 301018
rect -7516 300698 -7334 300934
rect -7098 300698 -6916 300934
rect -7516 265254 -6916 300698
rect -7516 265018 -7334 265254
rect -7098 265018 -6916 265254
rect -7516 264934 -6916 265018
rect -7516 264698 -7334 264934
rect -7098 264698 -6916 264934
rect -7516 229254 -6916 264698
rect -7516 229018 -7334 229254
rect -7098 229018 -6916 229254
rect -7516 228934 -6916 229018
rect -7516 228698 -7334 228934
rect -7098 228698 -6916 228934
rect -7516 193254 -6916 228698
rect -7516 193018 -7334 193254
rect -7098 193018 -6916 193254
rect -7516 192934 -6916 193018
rect -7516 192698 -7334 192934
rect -7098 192698 -6916 192934
rect -7516 157254 -6916 192698
rect -7516 157018 -7334 157254
rect -7098 157018 -6916 157254
rect -7516 156934 -6916 157018
rect -7516 156698 -7334 156934
rect -7098 156698 -6916 156934
rect -7516 121254 -6916 156698
rect -7516 121018 -7334 121254
rect -7098 121018 -6916 121254
rect -7516 120934 -6916 121018
rect -7516 120698 -7334 120934
rect -7098 120698 -6916 120934
rect -7516 85254 -6916 120698
rect -7516 85018 -7334 85254
rect -7098 85018 -6916 85254
rect -7516 84934 -6916 85018
rect -7516 84698 -7334 84934
rect -7098 84698 -6916 84934
rect -7516 49254 -6916 84698
rect -7516 49018 -7334 49254
rect -7098 49018 -6916 49254
rect -7516 48934 -6916 49018
rect -7516 48698 -7334 48934
rect -7098 48698 -6916 48934
rect -7516 13254 -6916 48698
rect -7516 13018 -7334 13254
rect -7098 13018 -6916 13254
rect -7516 12934 -6916 13018
rect -7516 12698 -7334 12934
rect -7098 12698 -6916 12934
rect -7516 -5866 -6916 12698
rect -6596 709438 -5996 709460
rect -6596 709202 -6414 709438
rect -6178 709202 -5996 709438
rect -6596 709118 -5996 709202
rect -6596 708882 -6414 709118
rect -6178 708882 -5996 709118
rect -6596 675654 -5996 708882
rect -6596 675418 -6414 675654
rect -6178 675418 -5996 675654
rect -6596 675334 -5996 675418
rect -6596 675098 -6414 675334
rect -6178 675098 -5996 675334
rect -6596 639654 -5996 675098
rect -6596 639418 -6414 639654
rect -6178 639418 -5996 639654
rect -6596 639334 -5996 639418
rect -6596 639098 -6414 639334
rect -6178 639098 -5996 639334
rect -6596 603654 -5996 639098
rect -6596 603418 -6414 603654
rect -6178 603418 -5996 603654
rect -6596 603334 -5996 603418
rect -6596 603098 -6414 603334
rect -6178 603098 -5996 603334
rect -6596 567654 -5996 603098
rect -6596 567418 -6414 567654
rect -6178 567418 -5996 567654
rect -6596 567334 -5996 567418
rect -6596 567098 -6414 567334
rect -6178 567098 -5996 567334
rect -6596 531654 -5996 567098
rect -6596 531418 -6414 531654
rect -6178 531418 -5996 531654
rect -6596 531334 -5996 531418
rect -6596 531098 -6414 531334
rect -6178 531098 -5996 531334
rect -6596 495654 -5996 531098
rect -6596 495418 -6414 495654
rect -6178 495418 -5996 495654
rect -6596 495334 -5996 495418
rect -6596 495098 -6414 495334
rect -6178 495098 -5996 495334
rect -6596 459654 -5996 495098
rect -6596 459418 -6414 459654
rect -6178 459418 -5996 459654
rect -6596 459334 -5996 459418
rect -6596 459098 -6414 459334
rect -6178 459098 -5996 459334
rect -6596 423654 -5996 459098
rect -6596 423418 -6414 423654
rect -6178 423418 -5996 423654
rect -6596 423334 -5996 423418
rect -6596 423098 -6414 423334
rect -6178 423098 -5996 423334
rect -6596 387654 -5996 423098
rect -6596 387418 -6414 387654
rect -6178 387418 -5996 387654
rect -6596 387334 -5996 387418
rect -6596 387098 -6414 387334
rect -6178 387098 -5996 387334
rect -6596 351654 -5996 387098
rect -6596 351418 -6414 351654
rect -6178 351418 -5996 351654
rect -6596 351334 -5996 351418
rect -6596 351098 -6414 351334
rect -6178 351098 -5996 351334
rect -6596 315654 -5996 351098
rect -6596 315418 -6414 315654
rect -6178 315418 -5996 315654
rect -6596 315334 -5996 315418
rect -6596 315098 -6414 315334
rect -6178 315098 -5996 315334
rect -6596 279654 -5996 315098
rect -6596 279418 -6414 279654
rect -6178 279418 -5996 279654
rect -6596 279334 -5996 279418
rect -6596 279098 -6414 279334
rect -6178 279098 -5996 279334
rect -6596 243654 -5996 279098
rect -6596 243418 -6414 243654
rect -6178 243418 -5996 243654
rect -6596 243334 -5996 243418
rect -6596 243098 -6414 243334
rect -6178 243098 -5996 243334
rect -6596 207654 -5996 243098
rect -6596 207418 -6414 207654
rect -6178 207418 -5996 207654
rect -6596 207334 -5996 207418
rect -6596 207098 -6414 207334
rect -6178 207098 -5996 207334
rect -6596 171654 -5996 207098
rect -6596 171418 -6414 171654
rect -6178 171418 -5996 171654
rect -6596 171334 -5996 171418
rect -6596 171098 -6414 171334
rect -6178 171098 -5996 171334
rect -6596 135654 -5996 171098
rect -6596 135418 -6414 135654
rect -6178 135418 -5996 135654
rect -6596 135334 -5996 135418
rect -6596 135098 -6414 135334
rect -6178 135098 -5996 135334
rect -6596 99654 -5996 135098
rect -6596 99418 -6414 99654
rect -6178 99418 -5996 99654
rect -6596 99334 -5996 99418
rect -6596 99098 -6414 99334
rect -6178 99098 -5996 99334
rect -6596 63654 -5996 99098
rect -6596 63418 -6414 63654
rect -6178 63418 -5996 63654
rect -6596 63334 -5996 63418
rect -6596 63098 -6414 63334
rect -6178 63098 -5996 63334
rect -6596 27654 -5996 63098
rect -6596 27418 -6414 27654
rect -6178 27418 -5996 27654
rect -6596 27334 -5996 27418
rect -6596 27098 -6414 27334
rect -6178 27098 -5996 27334
rect -6596 -4946 -5996 27098
rect -5676 708518 -5076 708540
rect -5676 708282 -5494 708518
rect -5258 708282 -5076 708518
rect -5676 708198 -5076 708282
rect -5676 707962 -5494 708198
rect -5258 707962 -5076 708198
rect -5676 693654 -5076 707962
rect 8004 708518 8604 709460
rect 8004 708282 8186 708518
rect 8422 708282 8604 708518
rect 8004 708198 8604 708282
rect 8004 707962 8186 708198
rect 8422 707962 8604 708198
rect -5676 693418 -5494 693654
rect -5258 693418 -5076 693654
rect -5676 693334 -5076 693418
rect -5676 693098 -5494 693334
rect -5258 693098 -5076 693334
rect -5676 657654 -5076 693098
rect -5676 657418 -5494 657654
rect -5258 657418 -5076 657654
rect -5676 657334 -5076 657418
rect -5676 657098 -5494 657334
rect -5258 657098 -5076 657334
rect -5676 621654 -5076 657098
rect -5676 621418 -5494 621654
rect -5258 621418 -5076 621654
rect -5676 621334 -5076 621418
rect -5676 621098 -5494 621334
rect -5258 621098 -5076 621334
rect -5676 585654 -5076 621098
rect -5676 585418 -5494 585654
rect -5258 585418 -5076 585654
rect -5676 585334 -5076 585418
rect -5676 585098 -5494 585334
rect -5258 585098 -5076 585334
rect -5676 549654 -5076 585098
rect -5676 549418 -5494 549654
rect -5258 549418 -5076 549654
rect -5676 549334 -5076 549418
rect -5676 549098 -5494 549334
rect -5258 549098 -5076 549334
rect -5676 513654 -5076 549098
rect -5676 513418 -5494 513654
rect -5258 513418 -5076 513654
rect -5676 513334 -5076 513418
rect -5676 513098 -5494 513334
rect -5258 513098 -5076 513334
rect -5676 477654 -5076 513098
rect -5676 477418 -5494 477654
rect -5258 477418 -5076 477654
rect -5676 477334 -5076 477418
rect -5676 477098 -5494 477334
rect -5258 477098 -5076 477334
rect -5676 441654 -5076 477098
rect -5676 441418 -5494 441654
rect -5258 441418 -5076 441654
rect -5676 441334 -5076 441418
rect -5676 441098 -5494 441334
rect -5258 441098 -5076 441334
rect -5676 405654 -5076 441098
rect -5676 405418 -5494 405654
rect -5258 405418 -5076 405654
rect -5676 405334 -5076 405418
rect -5676 405098 -5494 405334
rect -5258 405098 -5076 405334
rect -5676 369654 -5076 405098
rect -5676 369418 -5494 369654
rect -5258 369418 -5076 369654
rect -5676 369334 -5076 369418
rect -5676 369098 -5494 369334
rect -5258 369098 -5076 369334
rect -5676 333654 -5076 369098
rect -5676 333418 -5494 333654
rect -5258 333418 -5076 333654
rect -5676 333334 -5076 333418
rect -5676 333098 -5494 333334
rect -5258 333098 -5076 333334
rect -5676 297654 -5076 333098
rect -5676 297418 -5494 297654
rect -5258 297418 -5076 297654
rect -5676 297334 -5076 297418
rect -5676 297098 -5494 297334
rect -5258 297098 -5076 297334
rect -5676 261654 -5076 297098
rect -5676 261418 -5494 261654
rect -5258 261418 -5076 261654
rect -5676 261334 -5076 261418
rect -5676 261098 -5494 261334
rect -5258 261098 -5076 261334
rect -5676 225654 -5076 261098
rect -5676 225418 -5494 225654
rect -5258 225418 -5076 225654
rect -5676 225334 -5076 225418
rect -5676 225098 -5494 225334
rect -5258 225098 -5076 225334
rect -5676 189654 -5076 225098
rect -5676 189418 -5494 189654
rect -5258 189418 -5076 189654
rect -5676 189334 -5076 189418
rect -5676 189098 -5494 189334
rect -5258 189098 -5076 189334
rect -5676 153654 -5076 189098
rect -5676 153418 -5494 153654
rect -5258 153418 -5076 153654
rect -5676 153334 -5076 153418
rect -5676 153098 -5494 153334
rect -5258 153098 -5076 153334
rect -5676 117654 -5076 153098
rect -5676 117418 -5494 117654
rect -5258 117418 -5076 117654
rect -5676 117334 -5076 117418
rect -5676 117098 -5494 117334
rect -5258 117098 -5076 117334
rect -5676 81654 -5076 117098
rect -5676 81418 -5494 81654
rect -5258 81418 -5076 81654
rect -5676 81334 -5076 81418
rect -5676 81098 -5494 81334
rect -5258 81098 -5076 81334
rect -5676 45654 -5076 81098
rect -5676 45418 -5494 45654
rect -5258 45418 -5076 45654
rect -5676 45334 -5076 45418
rect -5676 45098 -5494 45334
rect -5258 45098 -5076 45334
rect -5676 9654 -5076 45098
rect -5676 9418 -5494 9654
rect -5258 9418 -5076 9654
rect -5676 9334 -5076 9418
rect -5676 9098 -5494 9334
rect -5258 9098 -5076 9334
rect -5676 -4026 -5076 9098
rect -4756 707598 -4156 707620
rect -4756 707362 -4574 707598
rect -4338 707362 -4156 707598
rect -4756 707278 -4156 707362
rect -4756 707042 -4574 707278
rect -4338 707042 -4156 707278
rect -4756 672054 -4156 707042
rect -4756 671818 -4574 672054
rect -4338 671818 -4156 672054
rect -4756 671734 -4156 671818
rect -4756 671498 -4574 671734
rect -4338 671498 -4156 671734
rect -4756 636054 -4156 671498
rect -4756 635818 -4574 636054
rect -4338 635818 -4156 636054
rect -4756 635734 -4156 635818
rect -4756 635498 -4574 635734
rect -4338 635498 -4156 635734
rect -4756 600054 -4156 635498
rect -4756 599818 -4574 600054
rect -4338 599818 -4156 600054
rect -4756 599734 -4156 599818
rect -4756 599498 -4574 599734
rect -4338 599498 -4156 599734
rect -4756 564054 -4156 599498
rect -4756 563818 -4574 564054
rect -4338 563818 -4156 564054
rect -4756 563734 -4156 563818
rect -4756 563498 -4574 563734
rect -4338 563498 -4156 563734
rect -4756 528054 -4156 563498
rect -4756 527818 -4574 528054
rect -4338 527818 -4156 528054
rect -4756 527734 -4156 527818
rect -4756 527498 -4574 527734
rect -4338 527498 -4156 527734
rect -4756 492054 -4156 527498
rect -4756 491818 -4574 492054
rect -4338 491818 -4156 492054
rect -4756 491734 -4156 491818
rect -4756 491498 -4574 491734
rect -4338 491498 -4156 491734
rect -4756 456054 -4156 491498
rect -4756 455818 -4574 456054
rect -4338 455818 -4156 456054
rect -4756 455734 -4156 455818
rect -4756 455498 -4574 455734
rect -4338 455498 -4156 455734
rect -4756 420054 -4156 455498
rect -4756 419818 -4574 420054
rect -4338 419818 -4156 420054
rect -4756 419734 -4156 419818
rect -4756 419498 -4574 419734
rect -4338 419498 -4156 419734
rect -4756 384054 -4156 419498
rect -4756 383818 -4574 384054
rect -4338 383818 -4156 384054
rect -4756 383734 -4156 383818
rect -4756 383498 -4574 383734
rect -4338 383498 -4156 383734
rect -4756 348054 -4156 383498
rect -4756 347818 -4574 348054
rect -4338 347818 -4156 348054
rect -4756 347734 -4156 347818
rect -4756 347498 -4574 347734
rect -4338 347498 -4156 347734
rect -4756 312054 -4156 347498
rect -4756 311818 -4574 312054
rect -4338 311818 -4156 312054
rect -4756 311734 -4156 311818
rect -4756 311498 -4574 311734
rect -4338 311498 -4156 311734
rect -4756 276054 -4156 311498
rect -4756 275818 -4574 276054
rect -4338 275818 -4156 276054
rect -4756 275734 -4156 275818
rect -4756 275498 -4574 275734
rect -4338 275498 -4156 275734
rect -4756 240054 -4156 275498
rect -4756 239818 -4574 240054
rect -4338 239818 -4156 240054
rect -4756 239734 -4156 239818
rect -4756 239498 -4574 239734
rect -4338 239498 -4156 239734
rect -4756 204054 -4156 239498
rect -4756 203818 -4574 204054
rect -4338 203818 -4156 204054
rect -4756 203734 -4156 203818
rect -4756 203498 -4574 203734
rect -4338 203498 -4156 203734
rect -4756 168054 -4156 203498
rect -4756 167818 -4574 168054
rect -4338 167818 -4156 168054
rect -4756 167734 -4156 167818
rect -4756 167498 -4574 167734
rect -4338 167498 -4156 167734
rect -4756 132054 -4156 167498
rect -4756 131818 -4574 132054
rect -4338 131818 -4156 132054
rect -4756 131734 -4156 131818
rect -4756 131498 -4574 131734
rect -4338 131498 -4156 131734
rect -4756 96054 -4156 131498
rect -4756 95818 -4574 96054
rect -4338 95818 -4156 96054
rect -4756 95734 -4156 95818
rect -4756 95498 -4574 95734
rect -4338 95498 -4156 95734
rect -4756 60054 -4156 95498
rect -4756 59818 -4574 60054
rect -4338 59818 -4156 60054
rect -4756 59734 -4156 59818
rect -4756 59498 -4574 59734
rect -4338 59498 -4156 59734
rect -4756 24054 -4156 59498
rect -4756 23818 -4574 24054
rect -4338 23818 -4156 24054
rect -4756 23734 -4156 23818
rect -4756 23498 -4574 23734
rect -4338 23498 -4156 23734
rect -4756 -3106 -4156 23498
rect -3836 706678 -3236 706700
rect -3836 706442 -3654 706678
rect -3418 706442 -3236 706678
rect -3836 706358 -3236 706442
rect -3836 706122 -3654 706358
rect -3418 706122 -3236 706358
rect -3836 690054 -3236 706122
rect 4404 706678 5004 707620
rect 4404 706442 4586 706678
rect 4822 706442 5004 706678
rect 4404 706358 5004 706442
rect 4404 706122 4586 706358
rect 4822 706122 5004 706358
rect -3836 689818 -3654 690054
rect -3418 689818 -3236 690054
rect -3836 689734 -3236 689818
rect -3836 689498 -3654 689734
rect -3418 689498 -3236 689734
rect -3836 654054 -3236 689498
rect -3836 653818 -3654 654054
rect -3418 653818 -3236 654054
rect -3836 653734 -3236 653818
rect -3836 653498 -3654 653734
rect -3418 653498 -3236 653734
rect -3836 618054 -3236 653498
rect -3836 617818 -3654 618054
rect -3418 617818 -3236 618054
rect -3836 617734 -3236 617818
rect -3836 617498 -3654 617734
rect -3418 617498 -3236 617734
rect -3836 582054 -3236 617498
rect -3836 581818 -3654 582054
rect -3418 581818 -3236 582054
rect -3836 581734 -3236 581818
rect -3836 581498 -3654 581734
rect -3418 581498 -3236 581734
rect -3836 546054 -3236 581498
rect -3836 545818 -3654 546054
rect -3418 545818 -3236 546054
rect -3836 545734 -3236 545818
rect -3836 545498 -3654 545734
rect -3418 545498 -3236 545734
rect -3836 510054 -3236 545498
rect -3836 509818 -3654 510054
rect -3418 509818 -3236 510054
rect -3836 509734 -3236 509818
rect -3836 509498 -3654 509734
rect -3418 509498 -3236 509734
rect -3836 474054 -3236 509498
rect -3836 473818 -3654 474054
rect -3418 473818 -3236 474054
rect -3836 473734 -3236 473818
rect -3836 473498 -3654 473734
rect -3418 473498 -3236 473734
rect -3836 438054 -3236 473498
rect -3836 437818 -3654 438054
rect -3418 437818 -3236 438054
rect -3836 437734 -3236 437818
rect -3836 437498 -3654 437734
rect -3418 437498 -3236 437734
rect -3836 402054 -3236 437498
rect -3836 401818 -3654 402054
rect -3418 401818 -3236 402054
rect -3836 401734 -3236 401818
rect -3836 401498 -3654 401734
rect -3418 401498 -3236 401734
rect -3836 366054 -3236 401498
rect -3836 365818 -3654 366054
rect -3418 365818 -3236 366054
rect -3836 365734 -3236 365818
rect -3836 365498 -3654 365734
rect -3418 365498 -3236 365734
rect -3836 330054 -3236 365498
rect -3836 329818 -3654 330054
rect -3418 329818 -3236 330054
rect -3836 329734 -3236 329818
rect -3836 329498 -3654 329734
rect -3418 329498 -3236 329734
rect -3836 294054 -3236 329498
rect -3836 293818 -3654 294054
rect -3418 293818 -3236 294054
rect -3836 293734 -3236 293818
rect -3836 293498 -3654 293734
rect -3418 293498 -3236 293734
rect -3836 258054 -3236 293498
rect -3836 257818 -3654 258054
rect -3418 257818 -3236 258054
rect -3836 257734 -3236 257818
rect -3836 257498 -3654 257734
rect -3418 257498 -3236 257734
rect -3836 222054 -3236 257498
rect -3836 221818 -3654 222054
rect -3418 221818 -3236 222054
rect -3836 221734 -3236 221818
rect -3836 221498 -3654 221734
rect -3418 221498 -3236 221734
rect -3836 186054 -3236 221498
rect -3836 185818 -3654 186054
rect -3418 185818 -3236 186054
rect -3836 185734 -3236 185818
rect -3836 185498 -3654 185734
rect -3418 185498 -3236 185734
rect -3836 150054 -3236 185498
rect -3836 149818 -3654 150054
rect -3418 149818 -3236 150054
rect -3836 149734 -3236 149818
rect -3836 149498 -3654 149734
rect -3418 149498 -3236 149734
rect -3836 114054 -3236 149498
rect -3836 113818 -3654 114054
rect -3418 113818 -3236 114054
rect -3836 113734 -3236 113818
rect -3836 113498 -3654 113734
rect -3418 113498 -3236 113734
rect -3836 78054 -3236 113498
rect -3836 77818 -3654 78054
rect -3418 77818 -3236 78054
rect -3836 77734 -3236 77818
rect -3836 77498 -3654 77734
rect -3418 77498 -3236 77734
rect -3836 42054 -3236 77498
rect -3836 41818 -3654 42054
rect -3418 41818 -3236 42054
rect -3836 41734 -3236 41818
rect -3836 41498 -3654 41734
rect -3418 41498 -3236 41734
rect -3836 6054 -3236 41498
rect -3836 5818 -3654 6054
rect -3418 5818 -3236 6054
rect -3836 5734 -3236 5818
rect -3836 5498 -3654 5734
rect -3418 5498 -3236 5734
rect -3836 -2186 -3236 5498
rect -2916 705758 -2316 705780
rect -2916 705522 -2734 705758
rect -2498 705522 -2316 705758
rect -2916 705438 -2316 705522
rect -2916 705202 -2734 705438
rect -2498 705202 -2316 705438
rect -2916 668454 -2316 705202
rect -2916 668218 -2734 668454
rect -2498 668218 -2316 668454
rect -2916 668134 -2316 668218
rect -2916 667898 -2734 668134
rect -2498 667898 -2316 668134
rect -2916 632454 -2316 667898
rect -2916 632218 -2734 632454
rect -2498 632218 -2316 632454
rect -2916 632134 -2316 632218
rect -2916 631898 -2734 632134
rect -2498 631898 -2316 632134
rect -2916 596454 -2316 631898
rect -2916 596218 -2734 596454
rect -2498 596218 -2316 596454
rect -2916 596134 -2316 596218
rect -2916 595898 -2734 596134
rect -2498 595898 -2316 596134
rect -2916 560454 -2316 595898
rect -2916 560218 -2734 560454
rect -2498 560218 -2316 560454
rect -2916 560134 -2316 560218
rect -2916 559898 -2734 560134
rect -2498 559898 -2316 560134
rect -2916 524454 -2316 559898
rect -2916 524218 -2734 524454
rect -2498 524218 -2316 524454
rect -2916 524134 -2316 524218
rect -2916 523898 -2734 524134
rect -2498 523898 -2316 524134
rect -2916 488454 -2316 523898
rect -2916 488218 -2734 488454
rect -2498 488218 -2316 488454
rect -2916 488134 -2316 488218
rect -2916 487898 -2734 488134
rect -2498 487898 -2316 488134
rect -2916 452454 -2316 487898
rect -2916 452218 -2734 452454
rect -2498 452218 -2316 452454
rect -2916 452134 -2316 452218
rect -2916 451898 -2734 452134
rect -2498 451898 -2316 452134
rect -2916 416454 -2316 451898
rect -2916 416218 -2734 416454
rect -2498 416218 -2316 416454
rect -2916 416134 -2316 416218
rect -2916 415898 -2734 416134
rect -2498 415898 -2316 416134
rect -2916 380454 -2316 415898
rect -2916 380218 -2734 380454
rect -2498 380218 -2316 380454
rect -2916 380134 -2316 380218
rect -2916 379898 -2734 380134
rect -2498 379898 -2316 380134
rect -2916 344454 -2316 379898
rect -2916 344218 -2734 344454
rect -2498 344218 -2316 344454
rect -2916 344134 -2316 344218
rect -2916 343898 -2734 344134
rect -2498 343898 -2316 344134
rect -2916 308454 -2316 343898
rect -2916 308218 -2734 308454
rect -2498 308218 -2316 308454
rect -2916 308134 -2316 308218
rect -2916 307898 -2734 308134
rect -2498 307898 -2316 308134
rect -2916 272454 -2316 307898
rect -2916 272218 -2734 272454
rect -2498 272218 -2316 272454
rect -2916 272134 -2316 272218
rect -2916 271898 -2734 272134
rect -2498 271898 -2316 272134
rect -2916 236454 -2316 271898
rect -2916 236218 -2734 236454
rect -2498 236218 -2316 236454
rect -2916 236134 -2316 236218
rect -2916 235898 -2734 236134
rect -2498 235898 -2316 236134
rect -2916 200454 -2316 235898
rect -2916 200218 -2734 200454
rect -2498 200218 -2316 200454
rect -2916 200134 -2316 200218
rect -2916 199898 -2734 200134
rect -2498 199898 -2316 200134
rect -2916 164454 -2316 199898
rect -2916 164218 -2734 164454
rect -2498 164218 -2316 164454
rect -2916 164134 -2316 164218
rect -2916 163898 -2734 164134
rect -2498 163898 -2316 164134
rect -2916 128454 -2316 163898
rect -2916 128218 -2734 128454
rect -2498 128218 -2316 128454
rect -2916 128134 -2316 128218
rect -2916 127898 -2734 128134
rect -2498 127898 -2316 128134
rect -2916 92454 -2316 127898
rect -2916 92218 -2734 92454
rect -2498 92218 -2316 92454
rect -2916 92134 -2316 92218
rect -2916 91898 -2734 92134
rect -2498 91898 -2316 92134
rect -2916 56454 -2316 91898
rect -2916 56218 -2734 56454
rect -2498 56218 -2316 56454
rect -2916 56134 -2316 56218
rect -2916 55898 -2734 56134
rect -2498 55898 -2316 56134
rect -2916 20454 -2316 55898
rect -2916 20218 -2734 20454
rect -2498 20218 -2316 20454
rect -2916 20134 -2316 20218
rect -2916 19898 -2734 20134
rect -2498 19898 -2316 20134
rect -2916 -1266 -2316 19898
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 686454 -1396 704282
rect -1996 686218 -1814 686454
rect -1578 686218 -1396 686454
rect -1996 686134 -1396 686218
rect -1996 685898 -1814 686134
rect -1578 685898 -1396 686134
rect -1996 650454 -1396 685898
rect -1996 650218 -1814 650454
rect -1578 650218 -1396 650454
rect -1996 650134 -1396 650218
rect -1996 649898 -1814 650134
rect -1578 649898 -1396 650134
rect -1996 614454 -1396 649898
rect -1996 614218 -1814 614454
rect -1578 614218 -1396 614454
rect -1996 614134 -1396 614218
rect -1996 613898 -1814 614134
rect -1578 613898 -1396 614134
rect -1996 578454 -1396 613898
rect -1996 578218 -1814 578454
rect -1578 578218 -1396 578454
rect -1996 578134 -1396 578218
rect -1996 577898 -1814 578134
rect -1578 577898 -1396 578134
rect -1996 542454 -1396 577898
rect -1996 542218 -1814 542454
rect -1578 542218 -1396 542454
rect -1996 542134 -1396 542218
rect -1996 541898 -1814 542134
rect -1578 541898 -1396 542134
rect -1996 506454 -1396 541898
rect -1996 506218 -1814 506454
rect -1578 506218 -1396 506454
rect -1996 506134 -1396 506218
rect -1996 505898 -1814 506134
rect -1578 505898 -1396 506134
rect -1996 470454 -1396 505898
rect -1996 470218 -1814 470454
rect -1578 470218 -1396 470454
rect -1996 470134 -1396 470218
rect -1996 469898 -1814 470134
rect -1578 469898 -1396 470134
rect -1996 434454 -1396 469898
rect -1996 434218 -1814 434454
rect -1578 434218 -1396 434454
rect -1996 434134 -1396 434218
rect -1996 433898 -1814 434134
rect -1578 433898 -1396 434134
rect -1996 398454 -1396 433898
rect -1996 398218 -1814 398454
rect -1578 398218 -1396 398454
rect -1996 398134 -1396 398218
rect -1996 397898 -1814 398134
rect -1578 397898 -1396 398134
rect -1996 362454 -1396 397898
rect -1996 362218 -1814 362454
rect -1578 362218 -1396 362454
rect -1996 362134 -1396 362218
rect -1996 361898 -1814 362134
rect -1578 361898 -1396 362134
rect -1996 326454 -1396 361898
rect -1996 326218 -1814 326454
rect -1578 326218 -1396 326454
rect -1996 326134 -1396 326218
rect -1996 325898 -1814 326134
rect -1578 325898 -1396 326134
rect -1996 290454 -1396 325898
rect -1996 290218 -1814 290454
rect -1578 290218 -1396 290454
rect -1996 290134 -1396 290218
rect -1996 289898 -1814 290134
rect -1578 289898 -1396 290134
rect -1996 254454 -1396 289898
rect -1996 254218 -1814 254454
rect -1578 254218 -1396 254454
rect -1996 254134 -1396 254218
rect -1996 253898 -1814 254134
rect -1578 253898 -1396 254134
rect -1996 218454 -1396 253898
rect -1996 218218 -1814 218454
rect -1578 218218 -1396 218454
rect -1996 218134 -1396 218218
rect -1996 217898 -1814 218134
rect -1578 217898 -1396 218134
rect -1996 182454 -1396 217898
rect -1996 182218 -1814 182454
rect -1578 182218 -1396 182454
rect -1996 182134 -1396 182218
rect -1996 181898 -1814 182134
rect -1578 181898 -1396 182134
rect -1996 146454 -1396 181898
rect -1996 146218 -1814 146454
rect -1578 146218 -1396 146454
rect -1996 146134 -1396 146218
rect -1996 145898 -1814 146134
rect -1578 145898 -1396 146134
rect -1996 110454 -1396 145898
rect -1996 110218 -1814 110454
rect -1578 110218 -1396 110454
rect -1996 110134 -1396 110218
rect -1996 109898 -1814 110134
rect -1578 109898 -1396 110134
rect -1996 74454 -1396 109898
rect -1996 74218 -1814 74454
rect -1578 74218 -1396 74454
rect -1996 74134 -1396 74218
rect -1996 73898 -1814 74134
rect -1578 73898 -1396 74134
rect -1996 38454 -1396 73898
rect -1996 38218 -1814 38454
rect -1578 38218 -1396 38454
rect -1996 38134 -1396 38218
rect -1996 37898 -1814 38134
rect -1578 37898 -1396 38134
rect -1996 2454 -1396 37898
rect -1996 2218 -1814 2454
rect -1578 2218 -1396 2454
rect -1996 2134 -1396 2218
rect -1996 1898 -1814 2134
rect -1578 1898 -1396 2134
rect -1996 -346 -1396 1898
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 804 704838 1404 705780
rect 804 704602 986 704838
rect 1222 704602 1404 704838
rect 804 704518 1404 704602
rect 804 704282 986 704518
rect 1222 704282 1404 704518
rect 804 686454 1404 704282
rect 804 686218 986 686454
rect 1222 686218 1404 686454
rect 804 686134 1404 686218
rect 804 685898 986 686134
rect 1222 685898 1404 686134
rect 804 650454 1404 685898
rect 804 650218 986 650454
rect 1222 650218 1404 650454
rect 804 650134 1404 650218
rect 804 649898 986 650134
rect 1222 649898 1404 650134
rect 804 614454 1404 649898
rect 804 614218 986 614454
rect 1222 614218 1404 614454
rect 804 614134 1404 614218
rect 804 613898 986 614134
rect 1222 613898 1404 614134
rect 804 578454 1404 613898
rect 804 578218 986 578454
rect 1222 578218 1404 578454
rect 804 578134 1404 578218
rect 804 577898 986 578134
rect 1222 577898 1404 578134
rect 804 542454 1404 577898
rect 804 542218 986 542454
rect 1222 542218 1404 542454
rect 804 542134 1404 542218
rect 804 541898 986 542134
rect 1222 541898 1404 542134
rect 804 506454 1404 541898
rect 804 506218 986 506454
rect 1222 506218 1404 506454
rect 804 506134 1404 506218
rect 804 505898 986 506134
rect 1222 505898 1404 506134
rect 804 470454 1404 505898
rect 804 470218 986 470454
rect 1222 470218 1404 470454
rect 804 470134 1404 470218
rect 804 469898 986 470134
rect 1222 469898 1404 470134
rect 804 434454 1404 469898
rect 804 434218 986 434454
rect 1222 434218 1404 434454
rect 804 434134 1404 434218
rect 804 433898 986 434134
rect 1222 433898 1404 434134
rect 804 398454 1404 433898
rect 804 398218 986 398454
rect 1222 398218 1404 398454
rect 804 398134 1404 398218
rect 804 397898 986 398134
rect 1222 397898 1404 398134
rect 804 362454 1404 397898
rect 804 362218 986 362454
rect 1222 362218 1404 362454
rect 804 362134 1404 362218
rect 804 361898 986 362134
rect 1222 361898 1404 362134
rect 804 326454 1404 361898
rect 804 326218 986 326454
rect 1222 326218 1404 326454
rect 804 326134 1404 326218
rect 804 325898 986 326134
rect 1222 325898 1404 326134
rect 804 290454 1404 325898
rect 804 290218 986 290454
rect 1222 290218 1404 290454
rect 804 290134 1404 290218
rect 804 289898 986 290134
rect 1222 289898 1404 290134
rect 804 254454 1404 289898
rect 804 254218 986 254454
rect 1222 254218 1404 254454
rect 804 254134 1404 254218
rect 804 253898 986 254134
rect 1222 253898 1404 254134
rect 804 218454 1404 253898
rect 804 218218 986 218454
rect 1222 218218 1404 218454
rect 804 218134 1404 218218
rect 804 217898 986 218134
rect 1222 217898 1404 218134
rect 804 182454 1404 217898
rect 804 182218 986 182454
rect 1222 182218 1404 182454
rect 804 182134 1404 182218
rect 804 181898 986 182134
rect 1222 181898 1404 182134
rect 804 146454 1404 181898
rect 804 146218 986 146454
rect 1222 146218 1404 146454
rect 804 146134 1404 146218
rect 804 145898 986 146134
rect 1222 145898 1404 146134
rect 804 110454 1404 145898
rect 804 110218 986 110454
rect 1222 110218 1404 110454
rect 804 110134 1404 110218
rect 804 109898 986 110134
rect 1222 109898 1404 110134
rect 804 74454 1404 109898
rect 804 74218 986 74454
rect 1222 74218 1404 74454
rect 804 74134 1404 74218
rect 804 73898 986 74134
rect 1222 73898 1404 74134
rect 804 38454 1404 73898
rect 804 38218 986 38454
rect 1222 38218 1404 38454
rect 804 38134 1404 38218
rect 804 37898 986 38134
rect 1222 37898 1404 38134
rect 804 2454 1404 37898
rect 804 2218 986 2454
rect 1222 2218 1404 2454
rect 804 2134 1404 2218
rect 804 1898 986 2134
rect 1222 1898 1404 2134
rect 804 -346 1404 1898
rect 804 -582 986 -346
rect 1222 -582 1404 -346
rect 804 -666 1404 -582
rect 804 -902 986 -666
rect 1222 -902 1404 -666
rect -2916 -1502 -2734 -1266
rect -2498 -1502 -2316 -1266
rect -2916 -1586 -2316 -1502
rect -2916 -1822 -2734 -1586
rect -2498 -1822 -2316 -1586
rect -2916 -1844 -2316 -1822
rect 804 -1844 1404 -902
rect 4404 690054 5004 706122
rect 4404 689818 4586 690054
rect 4822 689818 5004 690054
rect 4404 689734 5004 689818
rect 4404 689498 4586 689734
rect 4822 689498 5004 689734
rect 4404 654054 5004 689498
rect 4404 653818 4586 654054
rect 4822 653818 5004 654054
rect 4404 653734 5004 653818
rect 4404 653498 4586 653734
rect 4822 653498 5004 653734
rect 4404 618054 5004 653498
rect 4404 617818 4586 618054
rect 4822 617818 5004 618054
rect 4404 617734 5004 617818
rect 4404 617498 4586 617734
rect 4822 617498 5004 617734
rect 4404 582054 5004 617498
rect 4404 581818 4586 582054
rect 4822 581818 5004 582054
rect 4404 581734 5004 581818
rect 4404 581498 4586 581734
rect 4822 581498 5004 581734
rect 4404 546054 5004 581498
rect 8004 693654 8604 707962
rect 8004 693418 8186 693654
rect 8422 693418 8604 693654
rect 8004 693334 8604 693418
rect 8004 693098 8186 693334
rect 8422 693098 8604 693334
rect 8004 657654 8604 693098
rect 8004 657418 8186 657654
rect 8422 657418 8604 657654
rect 8004 657334 8604 657418
rect 8004 657098 8186 657334
rect 8422 657098 8604 657334
rect 8004 621654 8604 657098
rect 8004 621418 8186 621654
rect 8422 621418 8604 621654
rect 8004 621334 8604 621418
rect 8004 621098 8186 621334
rect 8422 621098 8604 621334
rect 8004 585654 8604 621098
rect 8004 585418 8186 585654
rect 8422 585418 8604 585654
rect 8004 585334 8604 585418
rect 8004 585098 8186 585334
rect 8422 585098 8604 585334
rect 4404 545818 4586 546054
rect 4822 545818 5004 546054
rect 4404 545734 5004 545818
rect 4404 545498 4586 545734
rect 4822 545498 5004 545734
rect 4404 510054 5004 545498
rect 4404 509818 4586 510054
rect 4822 509818 5004 510054
rect 4404 509734 5004 509818
rect 4404 509498 4586 509734
rect 4822 509498 5004 509734
rect 4404 474054 5004 509498
rect 4404 473818 4586 474054
rect 4822 473818 5004 474054
rect 4404 473734 5004 473818
rect 4404 473498 4586 473734
rect 4822 473498 5004 473734
rect 4404 438054 5004 473498
rect 4404 437818 4586 438054
rect 4822 437818 5004 438054
rect 4404 437734 5004 437818
rect 4404 437498 4586 437734
rect 4822 437498 5004 437734
rect 4404 402054 5004 437498
rect 4404 401818 4586 402054
rect 4822 401818 5004 402054
rect 4404 401734 5004 401818
rect 4404 401498 4586 401734
rect 4822 401498 5004 401734
rect 4404 366054 5004 401498
rect 4404 365818 4586 366054
rect 4822 365818 5004 366054
rect 4404 365734 5004 365818
rect 4404 365498 4586 365734
rect 4822 365498 5004 365734
rect 4404 330054 5004 365498
rect 4404 329818 4586 330054
rect 4822 329818 5004 330054
rect 4404 329734 5004 329818
rect 4404 329498 4586 329734
rect 4822 329498 5004 329734
rect 4404 294054 5004 329498
rect 4404 293818 4586 294054
rect 4822 293818 5004 294054
rect 4404 293734 5004 293818
rect 4404 293498 4586 293734
rect 4822 293498 5004 293734
rect 4404 258054 5004 293498
rect 4404 257818 4586 258054
rect 4822 257818 5004 258054
rect 4404 257734 5004 257818
rect 4404 257498 4586 257734
rect 4822 257498 5004 257734
rect 4404 222054 5004 257498
rect 4404 221818 4586 222054
rect 4822 221818 5004 222054
rect 4404 221734 5004 221818
rect 4404 221498 4586 221734
rect 4822 221498 5004 221734
rect 4404 186054 5004 221498
rect 4404 185818 4586 186054
rect 4822 185818 5004 186054
rect 4404 185734 5004 185818
rect 4404 185498 4586 185734
rect 4822 185498 5004 185734
rect 4404 150054 5004 185498
rect 4404 149818 4586 150054
rect 4822 149818 5004 150054
rect 4404 149734 5004 149818
rect 4404 149498 4586 149734
rect 4822 149498 5004 149734
rect 4404 114054 5004 149498
rect 4404 113818 4586 114054
rect 4822 113818 5004 114054
rect 4404 113734 5004 113818
rect 4404 113498 4586 113734
rect 4822 113498 5004 113734
rect 4404 78054 5004 113498
rect 4404 77818 4586 78054
rect 4822 77818 5004 78054
rect 4404 77734 5004 77818
rect 4404 77498 4586 77734
rect 4822 77498 5004 77734
rect 4404 42054 5004 77498
rect 4404 41818 4586 42054
rect 4822 41818 5004 42054
rect 4404 41734 5004 41818
rect 4404 41498 4586 41734
rect 4822 41498 5004 41734
rect 4404 6054 5004 41498
rect 4404 5818 4586 6054
rect 4822 5818 5004 6054
rect 4404 5734 5004 5818
rect 4404 5498 4586 5734
rect 4822 5498 5004 5734
rect -3836 -2422 -3654 -2186
rect -3418 -2422 -3236 -2186
rect -3836 -2506 -3236 -2422
rect -3836 -2742 -3654 -2506
rect -3418 -2742 -3236 -2506
rect -3836 -2764 -3236 -2742
rect 4404 -2186 5004 5498
rect 4404 -2422 4586 -2186
rect 4822 -2422 5004 -2186
rect 4404 -2506 5004 -2422
rect 4404 -2742 4586 -2506
rect 4822 -2742 5004 -2506
rect -4756 -3342 -4574 -3106
rect -4338 -3342 -4156 -3106
rect -4756 -3426 -4156 -3342
rect -4756 -3662 -4574 -3426
rect -4338 -3662 -4156 -3426
rect -4756 -3684 -4156 -3662
rect 4404 -3684 5004 -2742
rect 8004 549654 8604 585098
rect 8004 549418 8186 549654
rect 8422 549418 8604 549654
rect 8004 549334 8604 549418
rect 8004 549098 8186 549334
rect 8422 549098 8604 549334
rect 8004 513654 8604 549098
rect 8004 513418 8186 513654
rect 8422 513418 8604 513654
rect 8004 513334 8604 513418
rect 8004 513098 8186 513334
rect 8422 513098 8604 513334
rect 8004 477654 8604 513098
rect 8004 477418 8186 477654
rect 8422 477418 8604 477654
rect 8004 477334 8604 477418
rect 8004 477098 8186 477334
rect 8422 477098 8604 477334
rect 8004 441654 8604 477098
rect 8004 441418 8186 441654
rect 8422 441418 8604 441654
rect 8004 441334 8604 441418
rect 8004 441098 8186 441334
rect 8422 441098 8604 441334
rect 8004 405654 8604 441098
rect 8004 405418 8186 405654
rect 8422 405418 8604 405654
rect 8004 405334 8604 405418
rect 8004 405098 8186 405334
rect 8422 405098 8604 405334
rect 8004 369654 8604 405098
rect 8004 369418 8186 369654
rect 8422 369418 8604 369654
rect 8004 369334 8604 369418
rect 8004 369098 8186 369334
rect 8422 369098 8604 369334
rect 8004 333654 8604 369098
rect 8004 333418 8186 333654
rect 8422 333418 8604 333654
rect 8004 333334 8604 333418
rect 8004 333098 8186 333334
rect 8422 333098 8604 333334
rect 8004 297654 8604 333098
rect 8004 297418 8186 297654
rect 8422 297418 8604 297654
rect 8004 297334 8604 297418
rect 8004 297098 8186 297334
rect 8422 297098 8604 297334
rect 8004 261654 8604 297098
rect 8004 261418 8186 261654
rect 8422 261418 8604 261654
rect 8004 261334 8604 261418
rect 8004 261098 8186 261334
rect 8422 261098 8604 261334
rect 8004 225654 8604 261098
rect 8004 225418 8186 225654
rect 8422 225418 8604 225654
rect 8004 225334 8604 225418
rect 8004 225098 8186 225334
rect 8422 225098 8604 225334
rect 8004 189654 8604 225098
rect 8004 189418 8186 189654
rect 8422 189418 8604 189654
rect 8004 189334 8604 189418
rect 8004 189098 8186 189334
rect 8422 189098 8604 189334
rect 8004 153654 8604 189098
rect 8004 153418 8186 153654
rect 8422 153418 8604 153654
rect 8004 153334 8604 153418
rect 8004 153098 8186 153334
rect 8422 153098 8604 153334
rect 8004 117654 8604 153098
rect 8004 117418 8186 117654
rect 8422 117418 8604 117654
rect 8004 117334 8604 117418
rect 8004 117098 8186 117334
rect 8422 117098 8604 117334
rect 8004 81654 8604 117098
rect 8004 81418 8186 81654
rect 8422 81418 8604 81654
rect 8004 81334 8604 81418
rect 8004 81098 8186 81334
rect 8422 81098 8604 81334
rect 8004 45654 8604 81098
rect 8004 45418 8186 45654
rect 8422 45418 8604 45654
rect 8004 45334 8604 45418
rect 8004 45098 8186 45334
rect 8422 45098 8604 45334
rect 8004 9654 8604 45098
rect 8004 9418 8186 9654
rect 8422 9418 8604 9654
rect 8004 9334 8604 9418
rect 8004 9098 8186 9334
rect 8422 9098 8604 9334
rect -5676 -4262 -5494 -4026
rect -5258 -4262 -5076 -4026
rect -5676 -4346 -5076 -4262
rect -5676 -4582 -5494 -4346
rect -5258 -4582 -5076 -4346
rect -5676 -4604 -5076 -4582
rect 8004 -4026 8604 9098
rect 8004 -4262 8186 -4026
rect 8422 -4262 8604 -4026
rect 8004 -4346 8604 -4262
rect 8004 -4582 8186 -4346
rect 8422 -4582 8604 -4346
rect -6596 -5182 -6414 -4946
rect -6178 -5182 -5996 -4946
rect -6596 -5266 -5996 -5182
rect -6596 -5502 -6414 -5266
rect -6178 -5502 -5996 -5266
rect -6596 -5524 -5996 -5502
rect 8004 -5524 8604 -4582
rect 11604 697254 12204 709802
rect 29604 711278 30204 711300
rect 29604 711042 29786 711278
rect 30022 711042 30204 711278
rect 29604 710958 30204 711042
rect 29604 710722 29786 710958
rect 30022 710722 30204 710958
rect 26004 709438 26604 709460
rect 26004 709202 26186 709438
rect 26422 709202 26604 709438
rect 26004 709118 26604 709202
rect 26004 708882 26186 709118
rect 26422 708882 26604 709118
rect 22404 707598 23004 707620
rect 22404 707362 22586 707598
rect 22822 707362 23004 707598
rect 22404 707278 23004 707362
rect 22404 707042 22586 707278
rect 22822 707042 23004 707278
rect 11604 697018 11786 697254
rect 12022 697018 12204 697254
rect 11604 696934 12204 697018
rect 11604 696698 11786 696934
rect 12022 696698 12204 696934
rect 11604 661254 12204 696698
rect 11604 661018 11786 661254
rect 12022 661018 12204 661254
rect 11604 660934 12204 661018
rect 11604 660698 11786 660934
rect 12022 660698 12204 660934
rect 11604 625254 12204 660698
rect 11604 625018 11786 625254
rect 12022 625018 12204 625254
rect 11604 624934 12204 625018
rect 11604 624698 11786 624934
rect 12022 624698 12204 624934
rect 11604 589254 12204 624698
rect 11604 589018 11786 589254
rect 12022 589018 12204 589254
rect 11604 588934 12204 589018
rect 11604 588698 11786 588934
rect 12022 588698 12204 588934
rect 11604 553254 12204 588698
rect 11604 553018 11786 553254
rect 12022 553018 12204 553254
rect 11604 552934 12204 553018
rect 11604 552698 11786 552934
rect 12022 552698 12204 552934
rect 11604 517254 12204 552698
rect 11604 517018 11786 517254
rect 12022 517018 12204 517254
rect 11604 516934 12204 517018
rect 11604 516698 11786 516934
rect 12022 516698 12204 516934
rect 11604 481254 12204 516698
rect 11604 481018 11786 481254
rect 12022 481018 12204 481254
rect 11604 480934 12204 481018
rect 11604 480698 11786 480934
rect 12022 480698 12204 480934
rect 11604 445254 12204 480698
rect 11604 445018 11786 445254
rect 12022 445018 12204 445254
rect 11604 444934 12204 445018
rect 11604 444698 11786 444934
rect 12022 444698 12204 444934
rect 11604 409254 12204 444698
rect 11604 409018 11786 409254
rect 12022 409018 12204 409254
rect 11604 408934 12204 409018
rect 11604 408698 11786 408934
rect 12022 408698 12204 408934
rect 11604 373254 12204 408698
rect 11604 373018 11786 373254
rect 12022 373018 12204 373254
rect 11604 372934 12204 373018
rect 11604 372698 11786 372934
rect 12022 372698 12204 372934
rect 11604 337254 12204 372698
rect 11604 337018 11786 337254
rect 12022 337018 12204 337254
rect 11604 336934 12204 337018
rect 11604 336698 11786 336934
rect 12022 336698 12204 336934
rect 11604 301254 12204 336698
rect 11604 301018 11786 301254
rect 12022 301018 12204 301254
rect 11604 300934 12204 301018
rect 11604 300698 11786 300934
rect 12022 300698 12204 300934
rect 11604 265254 12204 300698
rect 11604 265018 11786 265254
rect 12022 265018 12204 265254
rect 11604 264934 12204 265018
rect 11604 264698 11786 264934
rect 12022 264698 12204 264934
rect 11604 229254 12204 264698
rect 11604 229018 11786 229254
rect 12022 229018 12204 229254
rect 11604 228934 12204 229018
rect 11604 228698 11786 228934
rect 12022 228698 12204 228934
rect 11604 193254 12204 228698
rect 11604 193018 11786 193254
rect 12022 193018 12204 193254
rect 11604 192934 12204 193018
rect 11604 192698 11786 192934
rect 12022 192698 12204 192934
rect 11604 157254 12204 192698
rect 11604 157018 11786 157254
rect 12022 157018 12204 157254
rect 11604 156934 12204 157018
rect 11604 156698 11786 156934
rect 12022 156698 12204 156934
rect 11604 121254 12204 156698
rect 11604 121018 11786 121254
rect 12022 121018 12204 121254
rect 11604 120934 12204 121018
rect 11604 120698 11786 120934
rect 12022 120698 12204 120934
rect 11604 85254 12204 120698
rect 11604 85018 11786 85254
rect 12022 85018 12204 85254
rect 11604 84934 12204 85018
rect 11604 84698 11786 84934
rect 12022 84698 12204 84934
rect 11604 49254 12204 84698
rect 11604 49018 11786 49254
rect 12022 49018 12204 49254
rect 11604 48934 12204 49018
rect 11604 48698 11786 48934
rect 12022 48698 12204 48934
rect 11604 13254 12204 48698
rect 11604 13018 11786 13254
rect 12022 13018 12204 13254
rect 11604 12934 12204 13018
rect 11604 12698 11786 12934
rect 12022 12698 12204 12934
rect -7516 -6102 -7334 -5866
rect -7098 -6102 -6916 -5866
rect -7516 -6186 -6916 -6102
rect -7516 -6422 -7334 -6186
rect -7098 -6422 -6916 -6186
rect -7516 -6444 -6916 -6422
rect 11604 -5866 12204 12698
rect 18804 705758 19404 705780
rect 18804 705522 18986 705758
rect 19222 705522 19404 705758
rect 18804 705438 19404 705522
rect 18804 705202 18986 705438
rect 19222 705202 19404 705438
rect 18804 668454 19404 705202
rect 18804 668218 18986 668454
rect 19222 668218 19404 668454
rect 18804 668134 19404 668218
rect 18804 667898 18986 668134
rect 19222 667898 19404 668134
rect 18804 632454 19404 667898
rect 18804 632218 18986 632454
rect 19222 632218 19404 632454
rect 18804 632134 19404 632218
rect 18804 631898 18986 632134
rect 19222 631898 19404 632134
rect 18804 596454 19404 631898
rect 18804 596218 18986 596454
rect 19222 596218 19404 596454
rect 18804 596134 19404 596218
rect 18804 595898 18986 596134
rect 19222 595898 19404 596134
rect 18804 560454 19404 595898
rect 18804 560218 18986 560454
rect 19222 560218 19404 560454
rect 18804 560134 19404 560218
rect 18804 559898 18986 560134
rect 19222 559898 19404 560134
rect 18804 524454 19404 559898
rect 18804 524218 18986 524454
rect 19222 524218 19404 524454
rect 18804 524134 19404 524218
rect 18804 523898 18986 524134
rect 19222 523898 19404 524134
rect 18804 488454 19404 523898
rect 18804 488218 18986 488454
rect 19222 488218 19404 488454
rect 18804 488134 19404 488218
rect 18804 487898 18986 488134
rect 19222 487898 19404 488134
rect 18804 452454 19404 487898
rect 18804 452218 18986 452454
rect 19222 452218 19404 452454
rect 18804 452134 19404 452218
rect 18804 451898 18986 452134
rect 19222 451898 19404 452134
rect 18804 416454 19404 451898
rect 18804 416218 18986 416454
rect 19222 416218 19404 416454
rect 18804 416134 19404 416218
rect 18804 415898 18986 416134
rect 19222 415898 19404 416134
rect 18804 380454 19404 415898
rect 18804 380218 18986 380454
rect 19222 380218 19404 380454
rect 18804 380134 19404 380218
rect 18804 379898 18986 380134
rect 19222 379898 19404 380134
rect 18804 344454 19404 379898
rect 18804 344218 18986 344454
rect 19222 344218 19404 344454
rect 18804 344134 19404 344218
rect 18804 343898 18986 344134
rect 19222 343898 19404 344134
rect 18804 308454 19404 343898
rect 18804 308218 18986 308454
rect 19222 308218 19404 308454
rect 18804 308134 19404 308218
rect 18804 307898 18986 308134
rect 19222 307898 19404 308134
rect 18804 272454 19404 307898
rect 18804 272218 18986 272454
rect 19222 272218 19404 272454
rect 18804 272134 19404 272218
rect 18804 271898 18986 272134
rect 19222 271898 19404 272134
rect 18804 236454 19404 271898
rect 18804 236218 18986 236454
rect 19222 236218 19404 236454
rect 18804 236134 19404 236218
rect 18804 235898 18986 236134
rect 19222 235898 19404 236134
rect 18804 200454 19404 235898
rect 18804 200218 18986 200454
rect 19222 200218 19404 200454
rect 18804 200134 19404 200218
rect 18804 199898 18986 200134
rect 19222 199898 19404 200134
rect 18804 164454 19404 199898
rect 18804 164218 18986 164454
rect 19222 164218 19404 164454
rect 18804 164134 19404 164218
rect 18804 163898 18986 164134
rect 19222 163898 19404 164134
rect 18804 128454 19404 163898
rect 18804 128218 18986 128454
rect 19222 128218 19404 128454
rect 18804 128134 19404 128218
rect 18804 127898 18986 128134
rect 19222 127898 19404 128134
rect 18804 92454 19404 127898
rect 18804 92218 18986 92454
rect 19222 92218 19404 92454
rect 18804 92134 19404 92218
rect 18804 91898 18986 92134
rect 19222 91898 19404 92134
rect 18804 56454 19404 91898
rect 18804 56218 18986 56454
rect 19222 56218 19404 56454
rect 18804 56134 19404 56218
rect 18804 55898 18986 56134
rect 19222 55898 19404 56134
rect 18804 20454 19404 55898
rect 18804 20218 18986 20454
rect 19222 20218 19404 20454
rect 18804 20134 19404 20218
rect 18804 19898 18986 20134
rect 19222 19898 19404 20134
rect 18804 -1266 19404 19898
rect 18804 -1502 18986 -1266
rect 19222 -1502 19404 -1266
rect 18804 -1586 19404 -1502
rect 18804 -1822 18986 -1586
rect 19222 -1822 19404 -1586
rect 18804 -1844 19404 -1822
rect 22404 672054 23004 707042
rect 22404 671818 22586 672054
rect 22822 671818 23004 672054
rect 22404 671734 23004 671818
rect 22404 671498 22586 671734
rect 22822 671498 23004 671734
rect 22404 636054 23004 671498
rect 22404 635818 22586 636054
rect 22822 635818 23004 636054
rect 22404 635734 23004 635818
rect 22404 635498 22586 635734
rect 22822 635498 23004 635734
rect 22404 600054 23004 635498
rect 22404 599818 22586 600054
rect 22822 599818 23004 600054
rect 22404 599734 23004 599818
rect 22404 599498 22586 599734
rect 22822 599498 23004 599734
rect 22404 564054 23004 599498
rect 22404 563818 22586 564054
rect 22822 563818 23004 564054
rect 22404 563734 23004 563818
rect 22404 563498 22586 563734
rect 22822 563498 23004 563734
rect 22404 528054 23004 563498
rect 22404 527818 22586 528054
rect 22822 527818 23004 528054
rect 22404 527734 23004 527818
rect 22404 527498 22586 527734
rect 22822 527498 23004 527734
rect 22404 492054 23004 527498
rect 22404 491818 22586 492054
rect 22822 491818 23004 492054
rect 22404 491734 23004 491818
rect 22404 491498 22586 491734
rect 22822 491498 23004 491734
rect 22404 456054 23004 491498
rect 22404 455818 22586 456054
rect 22822 455818 23004 456054
rect 22404 455734 23004 455818
rect 22404 455498 22586 455734
rect 22822 455498 23004 455734
rect 22404 420054 23004 455498
rect 22404 419818 22586 420054
rect 22822 419818 23004 420054
rect 22404 419734 23004 419818
rect 22404 419498 22586 419734
rect 22822 419498 23004 419734
rect 22404 384054 23004 419498
rect 22404 383818 22586 384054
rect 22822 383818 23004 384054
rect 22404 383734 23004 383818
rect 22404 383498 22586 383734
rect 22822 383498 23004 383734
rect 22404 348054 23004 383498
rect 22404 347818 22586 348054
rect 22822 347818 23004 348054
rect 22404 347734 23004 347818
rect 22404 347498 22586 347734
rect 22822 347498 23004 347734
rect 22404 312054 23004 347498
rect 22404 311818 22586 312054
rect 22822 311818 23004 312054
rect 22404 311734 23004 311818
rect 22404 311498 22586 311734
rect 22822 311498 23004 311734
rect 22404 276054 23004 311498
rect 22404 275818 22586 276054
rect 22822 275818 23004 276054
rect 22404 275734 23004 275818
rect 22404 275498 22586 275734
rect 22822 275498 23004 275734
rect 22404 240054 23004 275498
rect 22404 239818 22586 240054
rect 22822 239818 23004 240054
rect 22404 239734 23004 239818
rect 22404 239498 22586 239734
rect 22822 239498 23004 239734
rect 22404 204054 23004 239498
rect 22404 203818 22586 204054
rect 22822 203818 23004 204054
rect 22404 203734 23004 203818
rect 22404 203498 22586 203734
rect 22822 203498 23004 203734
rect 22404 168054 23004 203498
rect 22404 167818 22586 168054
rect 22822 167818 23004 168054
rect 22404 167734 23004 167818
rect 22404 167498 22586 167734
rect 22822 167498 23004 167734
rect 22404 132054 23004 167498
rect 22404 131818 22586 132054
rect 22822 131818 23004 132054
rect 22404 131734 23004 131818
rect 22404 131498 22586 131734
rect 22822 131498 23004 131734
rect 22404 96054 23004 131498
rect 22404 95818 22586 96054
rect 22822 95818 23004 96054
rect 22404 95734 23004 95818
rect 22404 95498 22586 95734
rect 22822 95498 23004 95734
rect 22404 60054 23004 95498
rect 22404 59818 22586 60054
rect 22822 59818 23004 60054
rect 22404 59734 23004 59818
rect 22404 59498 22586 59734
rect 22822 59498 23004 59734
rect 22404 24054 23004 59498
rect 22404 23818 22586 24054
rect 22822 23818 23004 24054
rect 22404 23734 23004 23818
rect 22404 23498 22586 23734
rect 22822 23498 23004 23734
rect 22404 -3106 23004 23498
rect 22404 -3342 22586 -3106
rect 22822 -3342 23004 -3106
rect 22404 -3426 23004 -3342
rect 22404 -3662 22586 -3426
rect 22822 -3662 23004 -3426
rect 22404 -3684 23004 -3662
rect 26004 675654 26604 708882
rect 26004 675418 26186 675654
rect 26422 675418 26604 675654
rect 26004 675334 26604 675418
rect 26004 675098 26186 675334
rect 26422 675098 26604 675334
rect 26004 639654 26604 675098
rect 26004 639418 26186 639654
rect 26422 639418 26604 639654
rect 26004 639334 26604 639418
rect 26004 639098 26186 639334
rect 26422 639098 26604 639334
rect 26004 603654 26604 639098
rect 26004 603418 26186 603654
rect 26422 603418 26604 603654
rect 26004 603334 26604 603418
rect 26004 603098 26186 603334
rect 26422 603098 26604 603334
rect 26004 567654 26604 603098
rect 26004 567418 26186 567654
rect 26422 567418 26604 567654
rect 26004 567334 26604 567418
rect 26004 567098 26186 567334
rect 26422 567098 26604 567334
rect 26004 531654 26604 567098
rect 26004 531418 26186 531654
rect 26422 531418 26604 531654
rect 26004 531334 26604 531418
rect 26004 531098 26186 531334
rect 26422 531098 26604 531334
rect 26004 495654 26604 531098
rect 26004 495418 26186 495654
rect 26422 495418 26604 495654
rect 26004 495334 26604 495418
rect 26004 495098 26186 495334
rect 26422 495098 26604 495334
rect 26004 459654 26604 495098
rect 26004 459418 26186 459654
rect 26422 459418 26604 459654
rect 26004 459334 26604 459418
rect 26004 459098 26186 459334
rect 26422 459098 26604 459334
rect 26004 423654 26604 459098
rect 26004 423418 26186 423654
rect 26422 423418 26604 423654
rect 26004 423334 26604 423418
rect 26004 423098 26186 423334
rect 26422 423098 26604 423334
rect 26004 387654 26604 423098
rect 26004 387418 26186 387654
rect 26422 387418 26604 387654
rect 26004 387334 26604 387418
rect 26004 387098 26186 387334
rect 26422 387098 26604 387334
rect 26004 351654 26604 387098
rect 26004 351418 26186 351654
rect 26422 351418 26604 351654
rect 26004 351334 26604 351418
rect 26004 351098 26186 351334
rect 26422 351098 26604 351334
rect 26004 315654 26604 351098
rect 26004 315418 26186 315654
rect 26422 315418 26604 315654
rect 26004 315334 26604 315418
rect 26004 315098 26186 315334
rect 26422 315098 26604 315334
rect 26004 279654 26604 315098
rect 26004 279418 26186 279654
rect 26422 279418 26604 279654
rect 26004 279334 26604 279418
rect 26004 279098 26186 279334
rect 26422 279098 26604 279334
rect 26004 243654 26604 279098
rect 26004 243418 26186 243654
rect 26422 243418 26604 243654
rect 26004 243334 26604 243418
rect 26004 243098 26186 243334
rect 26422 243098 26604 243334
rect 26004 207654 26604 243098
rect 26004 207418 26186 207654
rect 26422 207418 26604 207654
rect 26004 207334 26604 207418
rect 26004 207098 26186 207334
rect 26422 207098 26604 207334
rect 26004 171654 26604 207098
rect 26004 171418 26186 171654
rect 26422 171418 26604 171654
rect 26004 171334 26604 171418
rect 26004 171098 26186 171334
rect 26422 171098 26604 171334
rect 26004 135654 26604 171098
rect 26004 135418 26186 135654
rect 26422 135418 26604 135654
rect 26004 135334 26604 135418
rect 26004 135098 26186 135334
rect 26422 135098 26604 135334
rect 26004 99654 26604 135098
rect 26004 99418 26186 99654
rect 26422 99418 26604 99654
rect 26004 99334 26604 99418
rect 26004 99098 26186 99334
rect 26422 99098 26604 99334
rect 26004 63654 26604 99098
rect 26004 63418 26186 63654
rect 26422 63418 26604 63654
rect 26004 63334 26604 63418
rect 26004 63098 26186 63334
rect 26422 63098 26604 63334
rect 26004 27654 26604 63098
rect 26004 27418 26186 27654
rect 26422 27418 26604 27654
rect 26004 27334 26604 27418
rect 26004 27098 26186 27334
rect 26422 27098 26604 27334
rect 26004 -4946 26604 27098
rect 26004 -5182 26186 -4946
rect 26422 -5182 26604 -4946
rect 26004 -5266 26604 -5182
rect 26004 -5502 26186 -5266
rect 26422 -5502 26604 -5266
rect 26004 -5524 26604 -5502
rect 29604 679254 30204 710722
rect 47604 710358 48204 711300
rect 47604 710122 47786 710358
rect 48022 710122 48204 710358
rect 47604 710038 48204 710122
rect 47604 709802 47786 710038
rect 48022 709802 48204 710038
rect 44004 708518 44604 709460
rect 44004 708282 44186 708518
rect 44422 708282 44604 708518
rect 44004 708198 44604 708282
rect 44004 707962 44186 708198
rect 44422 707962 44604 708198
rect 40404 706678 41004 707620
rect 40404 706442 40586 706678
rect 40822 706442 41004 706678
rect 40404 706358 41004 706442
rect 40404 706122 40586 706358
rect 40822 706122 41004 706358
rect 29604 679018 29786 679254
rect 30022 679018 30204 679254
rect 29604 678934 30204 679018
rect 29604 678698 29786 678934
rect 30022 678698 30204 678934
rect 29604 643254 30204 678698
rect 29604 643018 29786 643254
rect 30022 643018 30204 643254
rect 29604 642934 30204 643018
rect 29604 642698 29786 642934
rect 30022 642698 30204 642934
rect 29604 607254 30204 642698
rect 29604 607018 29786 607254
rect 30022 607018 30204 607254
rect 29604 606934 30204 607018
rect 29604 606698 29786 606934
rect 30022 606698 30204 606934
rect 29604 571254 30204 606698
rect 29604 571018 29786 571254
rect 30022 571018 30204 571254
rect 29604 570934 30204 571018
rect 29604 570698 29786 570934
rect 30022 570698 30204 570934
rect 29604 535254 30204 570698
rect 29604 535018 29786 535254
rect 30022 535018 30204 535254
rect 29604 534934 30204 535018
rect 29604 534698 29786 534934
rect 30022 534698 30204 534934
rect 29604 499254 30204 534698
rect 29604 499018 29786 499254
rect 30022 499018 30204 499254
rect 29604 498934 30204 499018
rect 29604 498698 29786 498934
rect 30022 498698 30204 498934
rect 29604 463254 30204 498698
rect 29604 463018 29786 463254
rect 30022 463018 30204 463254
rect 29604 462934 30204 463018
rect 29604 462698 29786 462934
rect 30022 462698 30204 462934
rect 29604 427254 30204 462698
rect 29604 427018 29786 427254
rect 30022 427018 30204 427254
rect 29604 426934 30204 427018
rect 29604 426698 29786 426934
rect 30022 426698 30204 426934
rect 29604 391254 30204 426698
rect 29604 391018 29786 391254
rect 30022 391018 30204 391254
rect 29604 390934 30204 391018
rect 29604 390698 29786 390934
rect 30022 390698 30204 390934
rect 29604 355254 30204 390698
rect 29604 355018 29786 355254
rect 30022 355018 30204 355254
rect 29604 354934 30204 355018
rect 29604 354698 29786 354934
rect 30022 354698 30204 354934
rect 29604 319254 30204 354698
rect 29604 319018 29786 319254
rect 30022 319018 30204 319254
rect 29604 318934 30204 319018
rect 29604 318698 29786 318934
rect 30022 318698 30204 318934
rect 29604 283254 30204 318698
rect 29604 283018 29786 283254
rect 30022 283018 30204 283254
rect 29604 282934 30204 283018
rect 29604 282698 29786 282934
rect 30022 282698 30204 282934
rect 29604 247254 30204 282698
rect 29604 247018 29786 247254
rect 30022 247018 30204 247254
rect 29604 246934 30204 247018
rect 29604 246698 29786 246934
rect 30022 246698 30204 246934
rect 29604 211254 30204 246698
rect 29604 211018 29786 211254
rect 30022 211018 30204 211254
rect 29604 210934 30204 211018
rect 29604 210698 29786 210934
rect 30022 210698 30204 210934
rect 29604 175254 30204 210698
rect 29604 175018 29786 175254
rect 30022 175018 30204 175254
rect 29604 174934 30204 175018
rect 29604 174698 29786 174934
rect 30022 174698 30204 174934
rect 29604 139254 30204 174698
rect 29604 139018 29786 139254
rect 30022 139018 30204 139254
rect 29604 138934 30204 139018
rect 29604 138698 29786 138934
rect 30022 138698 30204 138934
rect 29604 103254 30204 138698
rect 29604 103018 29786 103254
rect 30022 103018 30204 103254
rect 29604 102934 30204 103018
rect 29604 102698 29786 102934
rect 30022 102698 30204 102934
rect 29604 67254 30204 102698
rect 29604 67018 29786 67254
rect 30022 67018 30204 67254
rect 29604 66934 30204 67018
rect 29604 66698 29786 66934
rect 30022 66698 30204 66934
rect 29604 31254 30204 66698
rect 29604 31018 29786 31254
rect 30022 31018 30204 31254
rect 29604 30934 30204 31018
rect 29604 30698 29786 30934
rect 30022 30698 30204 30934
rect 11604 -6102 11786 -5866
rect 12022 -6102 12204 -5866
rect 11604 -6186 12204 -6102
rect 11604 -6422 11786 -6186
rect 12022 -6422 12204 -6186
rect -8436 -7022 -8254 -6786
rect -8018 -7022 -7836 -6786
rect -8436 -7106 -7836 -7022
rect -8436 -7342 -8254 -7106
rect -8018 -7342 -7836 -7106
rect -8436 -7364 -7836 -7342
rect 11604 -7364 12204 -6422
rect 29604 -6786 30204 30698
rect 36804 704838 37404 705780
rect 36804 704602 36986 704838
rect 37222 704602 37404 704838
rect 36804 704518 37404 704602
rect 36804 704282 36986 704518
rect 37222 704282 37404 704518
rect 36804 686454 37404 704282
rect 36804 686218 36986 686454
rect 37222 686218 37404 686454
rect 36804 686134 37404 686218
rect 36804 685898 36986 686134
rect 37222 685898 37404 686134
rect 36804 650454 37404 685898
rect 36804 650218 36986 650454
rect 37222 650218 37404 650454
rect 36804 650134 37404 650218
rect 36804 649898 36986 650134
rect 37222 649898 37404 650134
rect 36804 614454 37404 649898
rect 36804 614218 36986 614454
rect 37222 614218 37404 614454
rect 36804 614134 37404 614218
rect 36804 613898 36986 614134
rect 37222 613898 37404 614134
rect 36804 578454 37404 613898
rect 36804 578218 36986 578454
rect 37222 578218 37404 578454
rect 36804 578134 37404 578218
rect 36804 577898 36986 578134
rect 37222 577898 37404 578134
rect 36804 542454 37404 577898
rect 36804 542218 36986 542454
rect 37222 542218 37404 542454
rect 36804 542134 37404 542218
rect 36804 541898 36986 542134
rect 37222 541898 37404 542134
rect 36804 506454 37404 541898
rect 36804 506218 36986 506454
rect 37222 506218 37404 506454
rect 36804 506134 37404 506218
rect 36804 505898 36986 506134
rect 37222 505898 37404 506134
rect 36804 470454 37404 505898
rect 36804 470218 36986 470454
rect 37222 470218 37404 470454
rect 36804 470134 37404 470218
rect 36804 469898 36986 470134
rect 37222 469898 37404 470134
rect 36804 434454 37404 469898
rect 36804 434218 36986 434454
rect 37222 434218 37404 434454
rect 36804 434134 37404 434218
rect 36804 433898 36986 434134
rect 37222 433898 37404 434134
rect 36804 398454 37404 433898
rect 36804 398218 36986 398454
rect 37222 398218 37404 398454
rect 36804 398134 37404 398218
rect 36804 397898 36986 398134
rect 37222 397898 37404 398134
rect 36804 362454 37404 397898
rect 36804 362218 36986 362454
rect 37222 362218 37404 362454
rect 36804 362134 37404 362218
rect 36804 361898 36986 362134
rect 37222 361898 37404 362134
rect 36804 326454 37404 361898
rect 36804 326218 36986 326454
rect 37222 326218 37404 326454
rect 36804 326134 37404 326218
rect 36804 325898 36986 326134
rect 37222 325898 37404 326134
rect 36804 290454 37404 325898
rect 36804 290218 36986 290454
rect 37222 290218 37404 290454
rect 36804 290134 37404 290218
rect 36804 289898 36986 290134
rect 37222 289898 37404 290134
rect 36804 254454 37404 289898
rect 36804 254218 36986 254454
rect 37222 254218 37404 254454
rect 36804 254134 37404 254218
rect 36804 253898 36986 254134
rect 37222 253898 37404 254134
rect 36804 218454 37404 253898
rect 36804 218218 36986 218454
rect 37222 218218 37404 218454
rect 36804 218134 37404 218218
rect 36804 217898 36986 218134
rect 37222 217898 37404 218134
rect 36804 182454 37404 217898
rect 36804 182218 36986 182454
rect 37222 182218 37404 182454
rect 36804 182134 37404 182218
rect 36804 181898 36986 182134
rect 37222 181898 37404 182134
rect 36804 146454 37404 181898
rect 36804 146218 36986 146454
rect 37222 146218 37404 146454
rect 36804 146134 37404 146218
rect 36804 145898 36986 146134
rect 37222 145898 37404 146134
rect 36804 110454 37404 145898
rect 36804 110218 36986 110454
rect 37222 110218 37404 110454
rect 36804 110134 37404 110218
rect 36804 109898 36986 110134
rect 37222 109898 37404 110134
rect 36804 74454 37404 109898
rect 36804 74218 36986 74454
rect 37222 74218 37404 74454
rect 36804 74134 37404 74218
rect 36804 73898 36986 74134
rect 37222 73898 37404 74134
rect 36804 38454 37404 73898
rect 36804 38218 36986 38454
rect 37222 38218 37404 38454
rect 36804 38134 37404 38218
rect 36804 37898 36986 38134
rect 37222 37898 37404 38134
rect 36804 2454 37404 37898
rect 36804 2218 36986 2454
rect 37222 2218 37404 2454
rect 36804 2134 37404 2218
rect 36804 1898 36986 2134
rect 37222 1898 37404 2134
rect 36804 -346 37404 1898
rect 36804 -582 36986 -346
rect 37222 -582 37404 -346
rect 36804 -666 37404 -582
rect 36804 -902 36986 -666
rect 37222 -902 37404 -666
rect 36804 -1844 37404 -902
rect 40404 690054 41004 706122
rect 40404 689818 40586 690054
rect 40822 689818 41004 690054
rect 40404 689734 41004 689818
rect 40404 689498 40586 689734
rect 40822 689498 41004 689734
rect 40404 654054 41004 689498
rect 40404 653818 40586 654054
rect 40822 653818 41004 654054
rect 40404 653734 41004 653818
rect 40404 653498 40586 653734
rect 40822 653498 41004 653734
rect 40404 618054 41004 653498
rect 40404 617818 40586 618054
rect 40822 617818 41004 618054
rect 40404 617734 41004 617818
rect 40404 617498 40586 617734
rect 40822 617498 41004 617734
rect 40404 582054 41004 617498
rect 40404 581818 40586 582054
rect 40822 581818 41004 582054
rect 40404 581734 41004 581818
rect 40404 581498 40586 581734
rect 40822 581498 41004 581734
rect 40404 546054 41004 581498
rect 40404 545818 40586 546054
rect 40822 545818 41004 546054
rect 40404 545734 41004 545818
rect 40404 545498 40586 545734
rect 40822 545498 41004 545734
rect 40404 510054 41004 545498
rect 40404 509818 40586 510054
rect 40822 509818 41004 510054
rect 40404 509734 41004 509818
rect 40404 509498 40586 509734
rect 40822 509498 41004 509734
rect 40404 474054 41004 509498
rect 40404 473818 40586 474054
rect 40822 473818 41004 474054
rect 40404 473734 41004 473818
rect 40404 473498 40586 473734
rect 40822 473498 41004 473734
rect 40404 438054 41004 473498
rect 40404 437818 40586 438054
rect 40822 437818 41004 438054
rect 40404 437734 41004 437818
rect 40404 437498 40586 437734
rect 40822 437498 41004 437734
rect 40404 402054 41004 437498
rect 40404 401818 40586 402054
rect 40822 401818 41004 402054
rect 40404 401734 41004 401818
rect 40404 401498 40586 401734
rect 40822 401498 41004 401734
rect 40404 366054 41004 401498
rect 40404 365818 40586 366054
rect 40822 365818 41004 366054
rect 40404 365734 41004 365818
rect 40404 365498 40586 365734
rect 40822 365498 41004 365734
rect 40404 330054 41004 365498
rect 40404 329818 40586 330054
rect 40822 329818 41004 330054
rect 40404 329734 41004 329818
rect 40404 329498 40586 329734
rect 40822 329498 41004 329734
rect 40404 294054 41004 329498
rect 40404 293818 40586 294054
rect 40822 293818 41004 294054
rect 40404 293734 41004 293818
rect 40404 293498 40586 293734
rect 40822 293498 41004 293734
rect 40404 258054 41004 293498
rect 40404 257818 40586 258054
rect 40822 257818 41004 258054
rect 40404 257734 41004 257818
rect 40404 257498 40586 257734
rect 40822 257498 41004 257734
rect 40404 222054 41004 257498
rect 40404 221818 40586 222054
rect 40822 221818 41004 222054
rect 40404 221734 41004 221818
rect 40404 221498 40586 221734
rect 40822 221498 41004 221734
rect 40404 186054 41004 221498
rect 40404 185818 40586 186054
rect 40822 185818 41004 186054
rect 40404 185734 41004 185818
rect 40404 185498 40586 185734
rect 40822 185498 41004 185734
rect 40404 150054 41004 185498
rect 40404 149818 40586 150054
rect 40822 149818 41004 150054
rect 40404 149734 41004 149818
rect 40404 149498 40586 149734
rect 40822 149498 41004 149734
rect 40404 114054 41004 149498
rect 40404 113818 40586 114054
rect 40822 113818 41004 114054
rect 40404 113734 41004 113818
rect 40404 113498 40586 113734
rect 40822 113498 41004 113734
rect 40404 78054 41004 113498
rect 40404 77818 40586 78054
rect 40822 77818 41004 78054
rect 40404 77734 41004 77818
rect 40404 77498 40586 77734
rect 40822 77498 41004 77734
rect 40404 42054 41004 77498
rect 40404 41818 40586 42054
rect 40822 41818 41004 42054
rect 40404 41734 41004 41818
rect 40404 41498 40586 41734
rect 40822 41498 41004 41734
rect 40404 6054 41004 41498
rect 40404 5818 40586 6054
rect 40822 5818 41004 6054
rect 40404 5734 41004 5818
rect 40404 5498 40586 5734
rect 40822 5498 41004 5734
rect 40404 -2186 41004 5498
rect 40404 -2422 40586 -2186
rect 40822 -2422 41004 -2186
rect 40404 -2506 41004 -2422
rect 40404 -2742 40586 -2506
rect 40822 -2742 41004 -2506
rect 40404 -3684 41004 -2742
rect 44004 693654 44604 707962
rect 44004 693418 44186 693654
rect 44422 693418 44604 693654
rect 44004 693334 44604 693418
rect 44004 693098 44186 693334
rect 44422 693098 44604 693334
rect 44004 657654 44604 693098
rect 44004 657418 44186 657654
rect 44422 657418 44604 657654
rect 44004 657334 44604 657418
rect 44004 657098 44186 657334
rect 44422 657098 44604 657334
rect 44004 621654 44604 657098
rect 44004 621418 44186 621654
rect 44422 621418 44604 621654
rect 44004 621334 44604 621418
rect 44004 621098 44186 621334
rect 44422 621098 44604 621334
rect 44004 585654 44604 621098
rect 44004 585418 44186 585654
rect 44422 585418 44604 585654
rect 44004 585334 44604 585418
rect 44004 585098 44186 585334
rect 44422 585098 44604 585334
rect 44004 549654 44604 585098
rect 44004 549418 44186 549654
rect 44422 549418 44604 549654
rect 44004 549334 44604 549418
rect 44004 549098 44186 549334
rect 44422 549098 44604 549334
rect 44004 513654 44604 549098
rect 44004 513418 44186 513654
rect 44422 513418 44604 513654
rect 44004 513334 44604 513418
rect 44004 513098 44186 513334
rect 44422 513098 44604 513334
rect 44004 477654 44604 513098
rect 44004 477418 44186 477654
rect 44422 477418 44604 477654
rect 44004 477334 44604 477418
rect 44004 477098 44186 477334
rect 44422 477098 44604 477334
rect 44004 441654 44604 477098
rect 44004 441418 44186 441654
rect 44422 441418 44604 441654
rect 44004 441334 44604 441418
rect 44004 441098 44186 441334
rect 44422 441098 44604 441334
rect 44004 405654 44604 441098
rect 44004 405418 44186 405654
rect 44422 405418 44604 405654
rect 44004 405334 44604 405418
rect 44004 405098 44186 405334
rect 44422 405098 44604 405334
rect 44004 369654 44604 405098
rect 44004 369418 44186 369654
rect 44422 369418 44604 369654
rect 44004 369334 44604 369418
rect 44004 369098 44186 369334
rect 44422 369098 44604 369334
rect 44004 333654 44604 369098
rect 44004 333418 44186 333654
rect 44422 333418 44604 333654
rect 44004 333334 44604 333418
rect 44004 333098 44186 333334
rect 44422 333098 44604 333334
rect 44004 297654 44604 333098
rect 44004 297418 44186 297654
rect 44422 297418 44604 297654
rect 44004 297334 44604 297418
rect 44004 297098 44186 297334
rect 44422 297098 44604 297334
rect 44004 261654 44604 297098
rect 44004 261418 44186 261654
rect 44422 261418 44604 261654
rect 44004 261334 44604 261418
rect 44004 261098 44186 261334
rect 44422 261098 44604 261334
rect 44004 225654 44604 261098
rect 44004 225418 44186 225654
rect 44422 225418 44604 225654
rect 44004 225334 44604 225418
rect 44004 225098 44186 225334
rect 44422 225098 44604 225334
rect 44004 189654 44604 225098
rect 44004 189418 44186 189654
rect 44422 189418 44604 189654
rect 44004 189334 44604 189418
rect 44004 189098 44186 189334
rect 44422 189098 44604 189334
rect 44004 153654 44604 189098
rect 44004 153418 44186 153654
rect 44422 153418 44604 153654
rect 44004 153334 44604 153418
rect 44004 153098 44186 153334
rect 44422 153098 44604 153334
rect 44004 117654 44604 153098
rect 44004 117418 44186 117654
rect 44422 117418 44604 117654
rect 44004 117334 44604 117418
rect 44004 117098 44186 117334
rect 44422 117098 44604 117334
rect 44004 81654 44604 117098
rect 44004 81418 44186 81654
rect 44422 81418 44604 81654
rect 44004 81334 44604 81418
rect 44004 81098 44186 81334
rect 44422 81098 44604 81334
rect 44004 45654 44604 81098
rect 44004 45418 44186 45654
rect 44422 45418 44604 45654
rect 44004 45334 44604 45418
rect 44004 45098 44186 45334
rect 44422 45098 44604 45334
rect 44004 9654 44604 45098
rect 44004 9418 44186 9654
rect 44422 9418 44604 9654
rect 44004 9334 44604 9418
rect 44004 9098 44186 9334
rect 44422 9098 44604 9334
rect 44004 -4026 44604 9098
rect 44004 -4262 44186 -4026
rect 44422 -4262 44604 -4026
rect 44004 -4346 44604 -4262
rect 44004 -4582 44186 -4346
rect 44422 -4582 44604 -4346
rect 44004 -5524 44604 -4582
rect 47604 697254 48204 709802
rect 65604 711278 66204 711300
rect 65604 711042 65786 711278
rect 66022 711042 66204 711278
rect 65604 710958 66204 711042
rect 65604 710722 65786 710958
rect 66022 710722 66204 710958
rect 62004 709438 62604 709460
rect 62004 709202 62186 709438
rect 62422 709202 62604 709438
rect 62004 709118 62604 709202
rect 62004 708882 62186 709118
rect 62422 708882 62604 709118
rect 58404 707598 59004 707620
rect 58404 707362 58586 707598
rect 58822 707362 59004 707598
rect 58404 707278 59004 707362
rect 58404 707042 58586 707278
rect 58822 707042 59004 707278
rect 47604 697018 47786 697254
rect 48022 697018 48204 697254
rect 47604 696934 48204 697018
rect 47604 696698 47786 696934
rect 48022 696698 48204 696934
rect 47604 661254 48204 696698
rect 47604 661018 47786 661254
rect 48022 661018 48204 661254
rect 47604 660934 48204 661018
rect 47604 660698 47786 660934
rect 48022 660698 48204 660934
rect 47604 625254 48204 660698
rect 47604 625018 47786 625254
rect 48022 625018 48204 625254
rect 47604 624934 48204 625018
rect 47604 624698 47786 624934
rect 48022 624698 48204 624934
rect 47604 589254 48204 624698
rect 47604 589018 47786 589254
rect 48022 589018 48204 589254
rect 47604 588934 48204 589018
rect 47604 588698 47786 588934
rect 48022 588698 48204 588934
rect 47604 553254 48204 588698
rect 54804 705758 55404 705780
rect 54804 705522 54986 705758
rect 55222 705522 55404 705758
rect 54804 705438 55404 705522
rect 54804 705202 54986 705438
rect 55222 705202 55404 705438
rect 54804 668454 55404 705202
rect 54804 668218 54986 668454
rect 55222 668218 55404 668454
rect 54804 668134 55404 668218
rect 54804 667898 54986 668134
rect 55222 667898 55404 668134
rect 54804 632454 55404 667898
rect 54804 632218 54986 632454
rect 55222 632218 55404 632454
rect 54804 632134 55404 632218
rect 54804 631898 54986 632134
rect 55222 631898 55404 632134
rect 54804 596454 55404 631898
rect 54804 596218 54986 596454
rect 55222 596218 55404 596454
rect 54804 596134 55404 596218
rect 54804 595898 54986 596134
rect 55222 595898 55404 596134
rect 47604 553018 47786 553254
rect 48022 553018 48204 553254
rect 47604 552934 48204 553018
rect 47604 552698 47786 552934
rect 48022 552698 48204 552934
rect 47604 517254 48204 552698
rect 47604 517018 47786 517254
rect 48022 517018 48204 517254
rect 47604 516934 48204 517018
rect 47604 516698 47786 516934
rect 48022 516698 48204 516934
rect 47604 481254 48204 516698
rect 47604 481018 47786 481254
rect 48022 481018 48204 481254
rect 47604 480934 48204 481018
rect 47604 480698 47786 480934
rect 48022 480698 48204 480934
rect 47604 445254 48204 480698
rect 47604 445018 47786 445254
rect 48022 445018 48204 445254
rect 47604 444934 48204 445018
rect 47604 444698 47786 444934
rect 48022 444698 48204 444934
rect 47604 409254 48204 444698
rect 47604 409018 47786 409254
rect 48022 409018 48204 409254
rect 47604 408934 48204 409018
rect 47604 408698 47786 408934
rect 48022 408698 48204 408934
rect 47604 373254 48204 408698
rect 47604 373018 47786 373254
rect 48022 373018 48204 373254
rect 47604 372934 48204 373018
rect 47604 372698 47786 372934
rect 48022 372698 48204 372934
rect 47604 337254 48204 372698
rect 47604 337018 47786 337254
rect 48022 337018 48204 337254
rect 47604 336934 48204 337018
rect 47604 336698 47786 336934
rect 48022 336698 48204 336934
rect 47604 301254 48204 336698
rect 47604 301018 47786 301254
rect 48022 301018 48204 301254
rect 47604 300934 48204 301018
rect 47604 300698 47786 300934
rect 48022 300698 48204 300934
rect 47604 265254 48204 300698
rect 47604 265018 47786 265254
rect 48022 265018 48204 265254
rect 47604 264934 48204 265018
rect 47604 264698 47786 264934
rect 48022 264698 48204 264934
rect 47604 229254 48204 264698
rect 47604 229018 47786 229254
rect 48022 229018 48204 229254
rect 47604 228934 48204 229018
rect 47604 228698 47786 228934
rect 48022 228698 48204 228934
rect 47604 193254 48204 228698
rect 47604 193018 47786 193254
rect 48022 193018 48204 193254
rect 47604 192934 48204 193018
rect 47604 192698 47786 192934
rect 48022 192698 48204 192934
rect 47604 157254 48204 192698
rect 47604 157018 47786 157254
rect 48022 157018 48204 157254
rect 47604 156934 48204 157018
rect 47604 156698 47786 156934
rect 48022 156698 48204 156934
rect 47604 121254 48204 156698
rect 47604 121018 47786 121254
rect 48022 121018 48204 121254
rect 47604 120934 48204 121018
rect 47604 120698 47786 120934
rect 48022 120698 48204 120934
rect 47604 85254 48204 120698
rect 47604 85018 47786 85254
rect 48022 85018 48204 85254
rect 47604 84934 48204 85018
rect 47604 84698 47786 84934
rect 48022 84698 48204 84934
rect 47604 49254 48204 84698
rect 47604 49018 47786 49254
rect 48022 49018 48204 49254
rect 47604 48934 48204 49018
rect 47604 48698 47786 48934
rect 48022 48698 48204 48934
rect 47604 13254 48204 48698
rect 47604 13018 47786 13254
rect 48022 13018 48204 13254
rect 47604 12934 48204 13018
rect 47604 12698 47786 12934
rect 48022 12698 48204 12934
rect 29604 -7022 29786 -6786
rect 30022 -7022 30204 -6786
rect 29604 -7106 30204 -7022
rect 29604 -7342 29786 -7106
rect 30022 -7342 30204 -7106
rect 29604 -7364 30204 -7342
rect 47604 -5866 48204 12698
rect 54804 560454 55404 595898
rect 54804 560218 54986 560454
rect 55222 560218 55404 560454
rect 54804 560134 55404 560218
rect 54804 559898 54986 560134
rect 55222 559898 55404 560134
rect 54804 524454 55404 559898
rect 54804 524218 54986 524454
rect 55222 524218 55404 524454
rect 54804 524134 55404 524218
rect 54804 523898 54986 524134
rect 55222 523898 55404 524134
rect 54804 488454 55404 523898
rect 54804 488218 54986 488454
rect 55222 488218 55404 488454
rect 54804 488134 55404 488218
rect 54804 487898 54986 488134
rect 55222 487898 55404 488134
rect 54804 452454 55404 487898
rect 54804 452218 54986 452454
rect 55222 452218 55404 452454
rect 54804 452134 55404 452218
rect 54804 451898 54986 452134
rect 55222 451898 55404 452134
rect 54804 416454 55404 451898
rect 54804 416218 54986 416454
rect 55222 416218 55404 416454
rect 54804 416134 55404 416218
rect 54804 415898 54986 416134
rect 55222 415898 55404 416134
rect 54804 380454 55404 415898
rect 54804 380218 54986 380454
rect 55222 380218 55404 380454
rect 54804 380134 55404 380218
rect 54804 379898 54986 380134
rect 55222 379898 55404 380134
rect 54804 344454 55404 379898
rect 54804 344218 54986 344454
rect 55222 344218 55404 344454
rect 54804 344134 55404 344218
rect 54804 343898 54986 344134
rect 55222 343898 55404 344134
rect 54804 308454 55404 343898
rect 54804 308218 54986 308454
rect 55222 308218 55404 308454
rect 54804 308134 55404 308218
rect 54804 307898 54986 308134
rect 55222 307898 55404 308134
rect 54804 272454 55404 307898
rect 54804 272218 54986 272454
rect 55222 272218 55404 272454
rect 54804 272134 55404 272218
rect 54804 271898 54986 272134
rect 55222 271898 55404 272134
rect 54804 236454 55404 271898
rect 54804 236218 54986 236454
rect 55222 236218 55404 236454
rect 54804 236134 55404 236218
rect 54804 235898 54986 236134
rect 55222 235898 55404 236134
rect 54804 200454 55404 235898
rect 54804 200218 54986 200454
rect 55222 200218 55404 200454
rect 54804 200134 55404 200218
rect 54804 199898 54986 200134
rect 55222 199898 55404 200134
rect 54804 164454 55404 199898
rect 54804 164218 54986 164454
rect 55222 164218 55404 164454
rect 54804 164134 55404 164218
rect 54804 163898 54986 164134
rect 55222 163898 55404 164134
rect 54804 128454 55404 163898
rect 54804 128218 54986 128454
rect 55222 128218 55404 128454
rect 54804 128134 55404 128218
rect 54804 127898 54986 128134
rect 55222 127898 55404 128134
rect 54804 92454 55404 127898
rect 54804 92218 54986 92454
rect 55222 92218 55404 92454
rect 54804 92134 55404 92218
rect 54804 91898 54986 92134
rect 55222 91898 55404 92134
rect 54804 56454 55404 91898
rect 54804 56218 54986 56454
rect 55222 56218 55404 56454
rect 54804 56134 55404 56218
rect 54804 55898 54986 56134
rect 55222 55898 55404 56134
rect 54804 20454 55404 55898
rect 54804 20218 54986 20454
rect 55222 20218 55404 20454
rect 54804 20134 55404 20218
rect 54804 19898 54986 20134
rect 55222 19898 55404 20134
rect 54804 -1266 55404 19898
rect 54804 -1502 54986 -1266
rect 55222 -1502 55404 -1266
rect 54804 -1586 55404 -1502
rect 54804 -1822 54986 -1586
rect 55222 -1822 55404 -1586
rect 54804 -1844 55404 -1822
rect 58404 672054 59004 707042
rect 58404 671818 58586 672054
rect 58822 671818 59004 672054
rect 58404 671734 59004 671818
rect 58404 671498 58586 671734
rect 58822 671498 59004 671734
rect 58404 636054 59004 671498
rect 58404 635818 58586 636054
rect 58822 635818 59004 636054
rect 58404 635734 59004 635818
rect 58404 635498 58586 635734
rect 58822 635498 59004 635734
rect 58404 600054 59004 635498
rect 58404 599818 58586 600054
rect 58822 599818 59004 600054
rect 58404 599734 59004 599818
rect 58404 599498 58586 599734
rect 58822 599498 59004 599734
rect 58404 564054 59004 599498
rect 58404 563818 58586 564054
rect 58822 563818 59004 564054
rect 58404 563734 59004 563818
rect 58404 563498 58586 563734
rect 58822 563498 59004 563734
rect 58404 528054 59004 563498
rect 58404 527818 58586 528054
rect 58822 527818 59004 528054
rect 58404 527734 59004 527818
rect 58404 527498 58586 527734
rect 58822 527498 59004 527734
rect 58404 492054 59004 527498
rect 58404 491818 58586 492054
rect 58822 491818 59004 492054
rect 58404 491734 59004 491818
rect 58404 491498 58586 491734
rect 58822 491498 59004 491734
rect 58404 456054 59004 491498
rect 58404 455818 58586 456054
rect 58822 455818 59004 456054
rect 58404 455734 59004 455818
rect 58404 455498 58586 455734
rect 58822 455498 59004 455734
rect 58404 420054 59004 455498
rect 58404 419818 58586 420054
rect 58822 419818 59004 420054
rect 58404 419734 59004 419818
rect 58404 419498 58586 419734
rect 58822 419498 59004 419734
rect 58404 384054 59004 419498
rect 58404 383818 58586 384054
rect 58822 383818 59004 384054
rect 58404 383734 59004 383818
rect 58404 383498 58586 383734
rect 58822 383498 59004 383734
rect 58404 348054 59004 383498
rect 58404 347818 58586 348054
rect 58822 347818 59004 348054
rect 58404 347734 59004 347818
rect 58404 347498 58586 347734
rect 58822 347498 59004 347734
rect 58404 312054 59004 347498
rect 58404 311818 58586 312054
rect 58822 311818 59004 312054
rect 58404 311734 59004 311818
rect 58404 311498 58586 311734
rect 58822 311498 59004 311734
rect 58404 276054 59004 311498
rect 58404 275818 58586 276054
rect 58822 275818 59004 276054
rect 58404 275734 59004 275818
rect 58404 275498 58586 275734
rect 58822 275498 59004 275734
rect 58404 240054 59004 275498
rect 58404 239818 58586 240054
rect 58822 239818 59004 240054
rect 58404 239734 59004 239818
rect 58404 239498 58586 239734
rect 58822 239498 59004 239734
rect 58404 204054 59004 239498
rect 58404 203818 58586 204054
rect 58822 203818 59004 204054
rect 58404 203734 59004 203818
rect 58404 203498 58586 203734
rect 58822 203498 59004 203734
rect 58404 168054 59004 203498
rect 58404 167818 58586 168054
rect 58822 167818 59004 168054
rect 58404 167734 59004 167818
rect 58404 167498 58586 167734
rect 58822 167498 59004 167734
rect 58404 132054 59004 167498
rect 58404 131818 58586 132054
rect 58822 131818 59004 132054
rect 58404 131734 59004 131818
rect 58404 131498 58586 131734
rect 58822 131498 59004 131734
rect 58404 96054 59004 131498
rect 58404 95818 58586 96054
rect 58822 95818 59004 96054
rect 58404 95734 59004 95818
rect 58404 95498 58586 95734
rect 58822 95498 59004 95734
rect 58404 60054 59004 95498
rect 58404 59818 58586 60054
rect 58822 59818 59004 60054
rect 58404 59734 59004 59818
rect 58404 59498 58586 59734
rect 58822 59498 59004 59734
rect 58404 24054 59004 59498
rect 58404 23818 58586 24054
rect 58822 23818 59004 24054
rect 58404 23734 59004 23818
rect 58404 23498 58586 23734
rect 58822 23498 59004 23734
rect 58404 -3106 59004 23498
rect 58404 -3342 58586 -3106
rect 58822 -3342 59004 -3106
rect 58404 -3426 59004 -3342
rect 58404 -3662 58586 -3426
rect 58822 -3662 59004 -3426
rect 58404 -3684 59004 -3662
rect 62004 675654 62604 708882
rect 62004 675418 62186 675654
rect 62422 675418 62604 675654
rect 62004 675334 62604 675418
rect 62004 675098 62186 675334
rect 62422 675098 62604 675334
rect 62004 639654 62604 675098
rect 62004 639418 62186 639654
rect 62422 639418 62604 639654
rect 62004 639334 62604 639418
rect 62004 639098 62186 639334
rect 62422 639098 62604 639334
rect 62004 603654 62604 639098
rect 62004 603418 62186 603654
rect 62422 603418 62604 603654
rect 62004 603334 62604 603418
rect 62004 603098 62186 603334
rect 62422 603098 62604 603334
rect 62004 567654 62604 603098
rect 62004 567418 62186 567654
rect 62422 567418 62604 567654
rect 62004 567334 62604 567418
rect 62004 567098 62186 567334
rect 62422 567098 62604 567334
rect 62004 531654 62604 567098
rect 62004 531418 62186 531654
rect 62422 531418 62604 531654
rect 62004 531334 62604 531418
rect 62004 531098 62186 531334
rect 62422 531098 62604 531334
rect 62004 495654 62604 531098
rect 62004 495418 62186 495654
rect 62422 495418 62604 495654
rect 62004 495334 62604 495418
rect 62004 495098 62186 495334
rect 62422 495098 62604 495334
rect 62004 459654 62604 495098
rect 62004 459418 62186 459654
rect 62422 459418 62604 459654
rect 62004 459334 62604 459418
rect 62004 459098 62186 459334
rect 62422 459098 62604 459334
rect 62004 423654 62604 459098
rect 62004 423418 62186 423654
rect 62422 423418 62604 423654
rect 62004 423334 62604 423418
rect 62004 423098 62186 423334
rect 62422 423098 62604 423334
rect 62004 387654 62604 423098
rect 62004 387418 62186 387654
rect 62422 387418 62604 387654
rect 62004 387334 62604 387418
rect 62004 387098 62186 387334
rect 62422 387098 62604 387334
rect 62004 351654 62604 387098
rect 62004 351418 62186 351654
rect 62422 351418 62604 351654
rect 62004 351334 62604 351418
rect 62004 351098 62186 351334
rect 62422 351098 62604 351334
rect 62004 315654 62604 351098
rect 62004 315418 62186 315654
rect 62422 315418 62604 315654
rect 62004 315334 62604 315418
rect 62004 315098 62186 315334
rect 62422 315098 62604 315334
rect 62004 279654 62604 315098
rect 62004 279418 62186 279654
rect 62422 279418 62604 279654
rect 62004 279334 62604 279418
rect 62004 279098 62186 279334
rect 62422 279098 62604 279334
rect 62004 243654 62604 279098
rect 62004 243418 62186 243654
rect 62422 243418 62604 243654
rect 62004 243334 62604 243418
rect 62004 243098 62186 243334
rect 62422 243098 62604 243334
rect 62004 207654 62604 243098
rect 62004 207418 62186 207654
rect 62422 207418 62604 207654
rect 62004 207334 62604 207418
rect 62004 207098 62186 207334
rect 62422 207098 62604 207334
rect 62004 171654 62604 207098
rect 62004 171418 62186 171654
rect 62422 171418 62604 171654
rect 62004 171334 62604 171418
rect 62004 171098 62186 171334
rect 62422 171098 62604 171334
rect 62004 135654 62604 171098
rect 62004 135418 62186 135654
rect 62422 135418 62604 135654
rect 62004 135334 62604 135418
rect 62004 135098 62186 135334
rect 62422 135098 62604 135334
rect 62004 99654 62604 135098
rect 62004 99418 62186 99654
rect 62422 99418 62604 99654
rect 62004 99334 62604 99418
rect 62004 99098 62186 99334
rect 62422 99098 62604 99334
rect 62004 63654 62604 99098
rect 62004 63418 62186 63654
rect 62422 63418 62604 63654
rect 62004 63334 62604 63418
rect 62004 63098 62186 63334
rect 62422 63098 62604 63334
rect 62004 27654 62604 63098
rect 62004 27418 62186 27654
rect 62422 27418 62604 27654
rect 62004 27334 62604 27418
rect 62004 27098 62186 27334
rect 62422 27098 62604 27334
rect 62004 -4946 62604 27098
rect 62004 -5182 62186 -4946
rect 62422 -5182 62604 -4946
rect 62004 -5266 62604 -5182
rect 62004 -5502 62186 -5266
rect 62422 -5502 62604 -5266
rect 62004 -5524 62604 -5502
rect 65604 679254 66204 710722
rect 83604 710358 84204 711300
rect 83604 710122 83786 710358
rect 84022 710122 84204 710358
rect 83604 710038 84204 710122
rect 83604 709802 83786 710038
rect 84022 709802 84204 710038
rect 80004 708518 80604 709460
rect 80004 708282 80186 708518
rect 80422 708282 80604 708518
rect 80004 708198 80604 708282
rect 80004 707962 80186 708198
rect 80422 707962 80604 708198
rect 76404 706678 77004 707620
rect 76404 706442 76586 706678
rect 76822 706442 77004 706678
rect 76404 706358 77004 706442
rect 76404 706122 76586 706358
rect 76822 706122 77004 706358
rect 65604 679018 65786 679254
rect 66022 679018 66204 679254
rect 65604 678934 66204 679018
rect 65604 678698 65786 678934
rect 66022 678698 66204 678934
rect 65604 643254 66204 678698
rect 65604 643018 65786 643254
rect 66022 643018 66204 643254
rect 65604 642934 66204 643018
rect 65604 642698 65786 642934
rect 66022 642698 66204 642934
rect 65604 607254 66204 642698
rect 65604 607018 65786 607254
rect 66022 607018 66204 607254
rect 65604 606934 66204 607018
rect 65604 606698 65786 606934
rect 66022 606698 66204 606934
rect 65604 571254 66204 606698
rect 65604 571018 65786 571254
rect 66022 571018 66204 571254
rect 65604 570934 66204 571018
rect 65604 570698 65786 570934
rect 66022 570698 66204 570934
rect 65604 535254 66204 570698
rect 65604 535018 65786 535254
rect 66022 535018 66204 535254
rect 65604 534934 66204 535018
rect 65604 534698 65786 534934
rect 66022 534698 66204 534934
rect 65604 499254 66204 534698
rect 65604 499018 65786 499254
rect 66022 499018 66204 499254
rect 65604 498934 66204 499018
rect 65604 498698 65786 498934
rect 66022 498698 66204 498934
rect 65604 463254 66204 498698
rect 65604 463018 65786 463254
rect 66022 463018 66204 463254
rect 65604 462934 66204 463018
rect 65604 462698 65786 462934
rect 66022 462698 66204 462934
rect 65604 427254 66204 462698
rect 65604 427018 65786 427254
rect 66022 427018 66204 427254
rect 65604 426934 66204 427018
rect 65604 426698 65786 426934
rect 66022 426698 66204 426934
rect 65604 391254 66204 426698
rect 65604 391018 65786 391254
rect 66022 391018 66204 391254
rect 65604 390934 66204 391018
rect 65604 390698 65786 390934
rect 66022 390698 66204 390934
rect 65604 355254 66204 390698
rect 65604 355018 65786 355254
rect 66022 355018 66204 355254
rect 65604 354934 66204 355018
rect 65604 354698 65786 354934
rect 66022 354698 66204 354934
rect 65604 319254 66204 354698
rect 65604 319018 65786 319254
rect 66022 319018 66204 319254
rect 65604 318934 66204 319018
rect 65604 318698 65786 318934
rect 66022 318698 66204 318934
rect 65604 283254 66204 318698
rect 65604 283018 65786 283254
rect 66022 283018 66204 283254
rect 65604 282934 66204 283018
rect 65604 282698 65786 282934
rect 66022 282698 66204 282934
rect 65604 247254 66204 282698
rect 65604 247018 65786 247254
rect 66022 247018 66204 247254
rect 65604 246934 66204 247018
rect 65604 246698 65786 246934
rect 66022 246698 66204 246934
rect 65604 211254 66204 246698
rect 65604 211018 65786 211254
rect 66022 211018 66204 211254
rect 65604 210934 66204 211018
rect 65604 210698 65786 210934
rect 66022 210698 66204 210934
rect 65604 175254 66204 210698
rect 65604 175018 65786 175254
rect 66022 175018 66204 175254
rect 65604 174934 66204 175018
rect 65604 174698 65786 174934
rect 66022 174698 66204 174934
rect 65604 139254 66204 174698
rect 65604 139018 65786 139254
rect 66022 139018 66204 139254
rect 65604 138934 66204 139018
rect 65604 138698 65786 138934
rect 66022 138698 66204 138934
rect 65604 103254 66204 138698
rect 65604 103018 65786 103254
rect 66022 103018 66204 103254
rect 65604 102934 66204 103018
rect 65604 102698 65786 102934
rect 66022 102698 66204 102934
rect 65604 67254 66204 102698
rect 65604 67018 65786 67254
rect 66022 67018 66204 67254
rect 65604 66934 66204 67018
rect 65604 66698 65786 66934
rect 66022 66698 66204 66934
rect 65604 31254 66204 66698
rect 65604 31018 65786 31254
rect 66022 31018 66204 31254
rect 65604 30934 66204 31018
rect 65604 30698 65786 30934
rect 66022 30698 66204 30934
rect 47604 -6102 47786 -5866
rect 48022 -6102 48204 -5866
rect 47604 -6186 48204 -6102
rect 47604 -6422 47786 -6186
rect 48022 -6422 48204 -6186
rect 47604 -7364 48204 -6422
rect 65604 -6786 66204 30698
rect 72804 704838 73404 705780
rect 72804 704602 72986 704838
rect 73222 704602 73404 704838
rect 72804 704518 73404 704602
rect 72804 704282 72986 704518
rect 73222 704282 73404 704518
rect 72804 686454 73404 704282
rect 72804 686218 72986 686454
rect 73222 686218 73404 686454
rect 72804 686134 73404 686218
rect 72804 685898 72986 686134
rect 73222 685898 73404 686134
rect 72804 650454 73404 685898
rect 72804 650218 72986 650454
rect 73222 650218 73404 650454
rect 72804 650134 73404 650218
rect 72804 649898 72986 650134
rect 73222 649898 73404 650134
rect 72804 614454 73404 649898
rect 72804 614218 72986 614454
rect 73222 614218 73404 614454
rect 72804 614134 73404 614218
rect 72804 613898 72986 614134
rect 73222 613898 73404 614134
rect 72804 578454 73404 613898
rect 72804 578218 72986 578454
rect 73222 578218 73404 578454
rect 72804 578134 73404 578218
rect 72804 577898 72986 578134
rect 73222 577898 73404 578134
rect 72804 542454 73404 577898
rect 72804 542218 72986 542454
rect 73222 542218 73404 542454
rect 72804 542134 73404 542218
rect 72804 541898 72986 542134
rect 73222 541898 73404 542134
rect 72804 506454 73404 541898
rect 72804 506218 72986 506454
rect 73222 506218 73404 506454
rect 72804 506134 73404 506218
rect 72804 505898 72986 506134
rect 73222 505898 73404 506134
rect 72804 470454 73404 505898
rect 72804 470218 72986 470454
rect 73222 470218 73404 470454
rect 72804 470134 73404 470218
rect 72804 469898 72986 470134
rect 73222 469898 73404 470134
rect 72804 434454 73404 469898
rect 72804 434218 72986 434454
rect 73222 434218 73404 434454
rect 72804 434134 73404 434218
rect 72804 433898 72986 434134
rect 73222 433898 73404 434134
rect 72804 398454 73404 433898
rect 72804 398218 72986 398454
rect 73222 398218 73404 398454
rect 72804 398134 73404 398218
rect 72804 397898 72986 398134
rect 73222 397898 73404 398134
rect 72804 362454 73404 397898
rect 72804 362218 72986 362454
rect 73222 362218 73404 362454
rect 72804 362134 73404 362218
rect 72804 361898 72986 362134
rect 73222 361898 73404 362134
rect 72804 326454 73404 361898
rect 72804 326218 72986 326454
rect 73222 326218 73404 326454
rect 72804 326134 73404 326218
rect 72804 325898 72986 326134
rect 73222 325898 73404 326134
rect 72804 290454 73404 325898
rect 72804 290218 72986 290454
rect 73222 290218 73404 290454
rect 72804 290134 73404 290218
rect 72804 289898 72986 290134
rect 73222 289898 73404 290134
rect 72804 254454 73404 289898
rect 72804 254218 72986 254454
rect 73222 254218 73404 254454
rect 72804 254134 73404 254218
rect 72804 253898 72986 254134
rect 73222 253898 73404 254134
rect 72804 218454 73404 253898
rect 72804 218218 72986 218454
rect 73222 218218 73404 218454
rect 72804 218134 73404 218218
rect 72804 217898 72986 218134
rect 73222 217898 73404 218134
rect 72804 182454 73404 217898
rect 72804 182218 72986 182454
rect 73222 182218 73404 182454
rect 72804 182134 73404 182218
rect 72804 181898 72986 182134
rect 73222 181898 73404 182134
rect 72804 146454 73404 181898
rect 72804 146218 72986 146454
rect 73222 146218 73404 146454
rect 72804 146134 73404 146218
rect 72804 145898 72986 146134
rect 73222 145898 73404 146134
rect 72804 110454 73404 145898
rect 72804 110218 72986 110454
rect 73222 110218 73404 110454
rect 72804 110134 73404 110218
rect 72804 109898 72986 110134
rect 73222 109898 73404 110134
rect 72804 74454 73404 109898
rect 72804 74218 72986 74454
rect 73222 74218 73404 74454
rect 72804 74134 73404 74218
rect 72804 73898 72986 74134
rect 73222 73898 73404 74134
rect 72804 38454 73404 73898
rect 72804 38218 72986 38454
rect 73222 38218 73404 38454
rect 72804 38134 73404 38218
rect 72804 37898 72986 38134
rect 73222 37898 73404 38134
rect 72804 2454 73404 37898
rect 72804 2218 72986 2454
rect 73222 2218 73404 2454
rect 72804 2134 73404 2218
rect 72804 1898 72986 2134
rect 73222 1898 73404 2134
rect 72804 -346 73404 1898
rect 72804 -582 72986 -346
rect 73222 -582 73404 -346
rect 72804 -666 73404 -582
rect 72804 -902 72986 -666
rect 73222 -902 73404 -666
rect 72804 -1844 73404 -902
rect 76404 690054 77004 706122
rect 76404 689818 76586 690054
rect 76822 689818 77004 690054
rect 76404 689734 77004 689818
rect 76404 689498 76586 689734
rect 76822 689498 77004 689734
rect 76404 654054 77004 689498
rect 76404 653818 76586 654054
rect 76822 653818 77004 654054
rect 76404 653734 77004 653818
rect 76404 653498 76586 653734
rect 76822 653498 77004 653734
rect 76404 618054 77004 653498
rect 76404 617818 76586 618054
rect 76822 617818 77004 618054
rect 76404 617734 77004 617818
rect 76404 617498 76586 617734
rect 76822 617498 77004 617734
rect 76404 582054 77004 617498
rect 76404 581818 76586 582054
rect 76822 581818 77004 582054
rect 76404 581734 77004 581818
rect 76404 581498 76586 581734
rect 76822 581498 77004 581734
rect 76404 546054 77004 581498
rect 76404 545818 76586 546054
rect 76822 545818 77004 546054
rect 76404 545734 77004 545818
rect 76404 545498 76586 545734
rect 76822 545498 77004 545734
rect 76404 510054 77004 545498
rect 76404 509818 76586 510054
rect 76822 509818 77004 510054
rect 76404 509734 77004 509818
rect 76404 509498 76586 509734
rect 76822 509498 77004 509734
rect 76404 474054 77004 509498
rect 76404 473818 76586 474054
rect 76822 473818 77004 474054
rect 76404 473734 77004 473818
rect 76404 473498 76586 473734
rect 76822 473498 77004 473734
rect 76404 438054 77004 473498
rect 76404 437818 76586 438054
rect 76822 437818 77004 438054
rect 76404 437734 77004 437818
rect 76404 437498 76586 437734
rect 76822 437498 77004 437734
rect 76404 402054 77004 437498
rect 76404 401818 76586 402054
rect 76822 401818 77004 402054
rect 76404 401734 77004 401818
rect 76404 401498 76586 401734
rect 76822 401498 77004 401734
rect 76404 366054 77004 401498
rect 76404 365818 76586 366054
rect 76822 365818 77004 366054
rect 76404 365734 77004 365818
rect 76404 365498 76586 365734
rect 76822 365498 77004 365734
rect 76404 330054 77004 365498
rect 76404 329818 76586 330054
rect 76822 329818 77004 330054
rect 76404 329734 77004 329818
rect 76404 329498 76586 329734
rect 76822 329498 77004 329734
rect 76404 294054 77004 329498
rect 76404 293818 76586 294054
rect 76822 293818 77004 294054
rect 76404 293734 77004 293818
rect 76404 293498 76586 293734
rect 76822 293498 77004 293734
rect 76404 258054 77004 293498
rect 76404 257818 76586 258054
rect 76822 257818 77004 258054
rect 76404 257734 77004 257818
rect 76404 257498 76586 257734
rect 76822 257498 77004 257734
rect 76404 222054 77004 257498
rect 76404 221818 76586 222054
rect 76822 221818 77004 222054
rect 76404 221734 77004 221818
rect 76404 221498 76586 221734
rect 76822 221498 77004 221734
rect 76404 186054 77004 221498
rect 76404 185818 76586 186054
rect 76822 185818 77004 186054
rect 76404 185734 77004 185818
rect 76404 185498 76586 185734
rect 76822 185498 77004 185734
rect 76404 150054 77004 185498
rect 76404 149818 76586 150054
rect 76822 149818 77004 150054
rect 76404 149734 77004 149818
rect 76404 149498 76586 149734
rect 76822 149498 77004 149734
rect 76404 114054 77004 149498
rect 76404 113818 76586 114054
rect 76822 113818 77004 114054
rect 76404 113734 77004 113818
rect 76404 113498 76586 113734
rect 76822 113498 77004 113734
rect 76404 78054 77004 113498
rect 76404 77818 76586 78054
rect 76822 77818 77004 78054
rect 76404 77734 77004 77818
rect 76404 77498 76586 77734
rect 76822 77498 77004 77734
rect 76404 42054 77004 77498
rect 76404 41818 76586 42054
rect 76822 41818 77004 42054
rect 76404 41734 77004 41818
rect 76404 41498 76586 41734
rect 76822 41498 77004 41734
rect 76404 6054 77004 41498
rect 76404 5818 76586 6054
rect 76822 5818 77004 6054
rect 76404 5734 77004 5818
rect 76404 5498 76586 5734
rect 76822 5498 77004 5734
rect 76404 -2186 77004 5498
rect 76404 -2422 76586 -2186
rect 76822 -2422 77004 -2186
rect 76404 -2506 77004 -2422
rect 76404 -2742 76586 -2506
rect 76822 -2742 77004 -2506
rect 76404 -3684 77004 -2742
rect 80004 693654 80604 707962
rect 80004 693418 80186 693654
rect 80422 693418 80604 693654
rect 80004 693334 80604 693418
rect 80004 693098 80186 693334
rect 80422 693098 80604 693334
rect 80004 657654 80604 693098
rect 80004 657418 80186 657654
rect 80422 657418 80604 657654
rect 80004 657334 80604 657418
rect 80004 657098 80186 657334
rect 80422 657098 80604 657334
rect 80004 621654 80604 657098
rect 80004 621418 80186 621654
rect 80422 621418 80604 621654
rect 80004 621334 80604 621418
rect 80004 621098 80186 621334
rect 80422 621098 80604 621334
rect 80004 585654 80604 621098
rect 80004 585418 80186 585654
rect 80422 585418 80604 585654
rect 80004 585334 80604 585418
rect 80004 585098 80186 585334
rect 80422 585098 80604 585334
rect 80004 549654 80604 585098
rect 80004 549418 80186 549654
rect 80422 549418 80604 549654
rect 80004 549334 80604 549418
rect 80004 549098 80186 549334
rect 80422 549098 80604 549334
rect 80004 513654 80604 549098
rect 80004 513418 80186 513654
rect 80422 513418 80604 513654
rect 80004 513334 80604 513418
rect 80004 513098 80186 513334
rect 80422 513098 80604 513334
rect 80004 477654 80604 513098
rect 80004 477418 80186 477654
rect 80422 477418 80604 477654
rect 80004 477334 80604 477418
rect 80004 477098 80186 477334
rect 80422 477098 80604 477334
rect 80004 441654 80604 477098
rect 80004 441418 80186 441654
rect 80422 441418 80604 441654
rect 80004 441334 80604 441418
rect 80004 441098 80186 441334
rect 80422 441098 80604 441334
rect 80004 405654 80604 441098
rect 80004 405418 80186 405654
rect 80422 405418 80604 405654
rect 80004 405334 80604 405418
rect 80004 405098 80186 405334
rect 80422 405098 80604 405334
rect 80004 369654 80604 405098
rect 80004 369418 80186 369654
rect 80422 369418 80604 369654
rect 80004 369334 80604 369418
rect 80004 369098 80186 369334
rect 80422 369098 80604 369334
rect 80004 333654 80604 369098
rect 80004 333418 80186 333654
rect 80422 333418 80604 333654
rect 80004 333334 80604 333418
rect 80004 333098 80186 333334
rect 80422 333098 80604 333334
rect 80004 297654 80604 333098
rect 80004 297418 80186 297654
rect 80422 297418 80604 297654
rect 80004 297334 80604 297418
rect 80004 297098 80186 297334
rect 80422 297098 80604 297334
rect 80004 261654 80604 297098
rect 80004 261418 80186 261654
rect 80422 261418 80604 261654
rect 80004 261334 80604 261418
rect 80004 261098 80186 261334
rect 80422 261098 80604 261334
rect 80004 225654 80604 261098
rect 80004 225418 80186 225654
rect 80422 225418 80604 225654
rect 80004 225334 80604 225418
rect 80004 225098 80186 225334
rect 80422 225098 80604 225334
rect 80004 189654 80604 225098
rect 80004 189418 80186 189654
rect 80422 189418 80604 189654
rect 80004 189334 80604 189418
rect 80004 189098 80186 189334
rect 80422 189098 80604 189334
rect 80004 153654 80604 189098
rect 80004 153418 80186 153654
rect 80422 153418 80604 153654
rect 80004 153334 80604 153418
rect 80004 153098 80186 153334
rect 80422 153098 80604 153334
rect 80004 117654 80604 153098
rect 80004 117418 80186 117654
rect 80422 117418 80604 117654
rect 80004 117334 80604 117418
rect 80004 117098 80186 117334
rect 80422 117098 80604 117334
rect 80004 81654 80604 117098
rect 80004 81418 80186 81654
rect 80422 81418 80604 81654
rect 80004 81334 80604 81418
rect 80004 81098 80186 81334
rect 80422 81098 80604 81334
rect 80004 45654 80604 81098
rect 80004 45418 80186 45654
rect 80422 45418 80604 45654
rect 80004 45334 80604 45418
rect 80004 45098 80186 45334
rect 80422 45098 80604 45334
rect 80004 9654 80604 45098
rect 80004 9418 80186 9654
rect 80422 9418 80604 9654
rect 80004 9334 80604 9418
rect 80004 9098 80186 9334
rect 80422 9098 80604 9334
rect 80004 -4026 80604 9098
rect 80004 -4262 80186 -4026
rect 80422 -4262 80604 -4026
rect 80004 -4346 80604 -4262
rect 80004 -4582 80186 -4346
rect 80422 -4582 80604 -4346
rect 80004 -5524 80604 -4582
rect 83604 697254 84204 709802
rect 101604 711278 102204 711300
rect 101604 711042 101786 711278
rect 102022 711042 102204 711278
rect 101604 710958 102204 711042
rect 101604 710722 101786 710958
rect 102022 710722 102204 710958
rect 98004 709438 98604 709460
rect 98004 709202 98186 709438
rect 98422 709202 98604 709438
rect 98004 709118 98604 709202
rect 98004 708882 98186 709118
rect 98422 708882 98604 709118
rect 94404 707598 95004 707620
rect 94404 707362 94586 707598
rect 94822 707362 95004 707598
rect 94404 707278 95004 707362
rect 94404 707042 94586 707278
rect 94822 707042 95004 707278
rect 83604 697018 83786 697254
rect 84022 697018 84204 697254
rect 83604 696934 84204 697018
rect 83604 696698 83786 696934
rect 84022 696698 84204 696934
rect 83604 661254 84204 696698
rect 83604 661018 83786 661254
rect 84022 661018 84204 661254
rect 83604 660934 84204 661018
rect 83604 660698 83786 660934
rect 84022 660698 84204 660934
rect 83604 625254 84204 660698
rect 83604 625018 83786 625254
rect 84022 625018 84204 625254
rect 83604 624934 84204 625018
rect 83604 624698 83786 624934
rect 84022 624698 84204 624934
rect 83604 589254 84204 624698
rect 83604 589018 83786 589254
rect 84022 589018 84204 589254
rect 83604 588934 84204 589018
rect 83604 588698 83786 588934
rect 84022 588698 84204 588934
rect 83604 553254 84204 588698
rect 90804 705758 91404 705780
rect 90804 705522 90986 705758
rect 91222 705522 91404 705758
rect 90804 705438 91404 705522
rect 90804 705202 90986 705438
rect 91222 705202 91404 705438
rect 90804 668454 91404 705202
rect 90804 668218 90986 668454
rect 91222 668218 91404 668454
rect 90804 668134 91404 668218
rect 90804 667898 90986 668134
rect 91222 667898 91404 668134
rect 90804 632454 91404 667898
rect 90804 632218 90986 632454
rect 91222 632218 91404 632454
rect 90804 632134 91404 632218
rect 90804 631898 90986 632134
rect 91222 631898 91404 632134
rect 90804 596454 91404 631898
rect 90804 596218 90986 596454
rect 91222 596218 91404 596454
rect 90804 596134 91404 596218
rect 90804 595898 90986 596134
rect 91222 595898 91404 596134
rect 83604 553018 83786 553254
rect 84022 553018 84204 553254
rect 83604 552934 84204 553018
rect 83604 552698 83786 552934
rect 84022 552698 84204 552934
rect 83604 517254 84204 552698
rect 83604 517018 83786 517254
rect 84022 517018 84204 517254
rect 83604 516934 84204 517018
rect 83604 516698 83786 516934
rect 84022 516698 84204 516934
rect 83604 481254 84204 516698
rect 83604 481018 83786 481254
rect 84022 481018 84204 481254
rect 83604 480934 84204 481018
rect 83604 480698 83786 480934
rect 84022 480698 84204 480934
rect 83604 445254 84204 480698
rect 83604 445018 83786 445254
rect 84022 445018 84204 445254
rect 83604 444934 84204 445018
rect 83604 444698 83786 444934
rect 84022 444698 84204 444934
rect 83604 409254 84204 444698
rect 83604 409018 83786 409254
rect 84022 409018 84204 409254
rect 83604 408934 84204 409018
rect 83604 408698 83786 408934
rect 84022 408698 84204 408934
rect 83604 373254 84204 408698
rect 83604 373018 83786 373254
rect 84022 373018 84204 373254
rect 83604 372934 84204 373018
rect 83604 372698 83786 372934
rect 84022 372698 84204 372934
rect 83604 337254 84204 372698
rect 83604 337018 83786 337254
rect 84022 337018 84204 337254
rect 83604 336934 84204 337018
rect 83604 336698 83786 336934
rect 84022 336698 84204 336934
rect 83604 301254 84204 336698
rect 83604 301018 83786 301254
rect 84022 301018 84204 301254
rect 83604 300934 84204 301018
rect 83604 300698 83786 300934
rect 84022 300698 84204 300934
rect 83604 265254 84204 300698
rect 83604 265018 83786 265254
rect 84022 265018 84204 265254
rect 83604 264934 84204 265018
rect 83604 264698 83786 264934
rect 84022 264698 84204 264934
rect 83604 229254 84204 264698
rect 83604 229018 83786 229254
rect 84022 229018 84204 229254
rect 83604 228934 84204 229018
rect 83604 228698 83786 228934
rect 84022 228698 84204 228934
rect 83604 193254 84204 228698
rect 83604 193018 83786 193254
rect 84022 193018 84204 193254
rect 83604 192934 84204 193018
rect 83604 192698 83786 192934
rect 84022 192698 84204 192934
rect 83604 157254 84204 192698
rect 83604 157018 83786 157254
rect 84022 157018 84204 157254
rect 83604 156934 84204 157018
rect 83604 156698 83786 156934
rect 84022 156698 84204 156934
rect 83604 121254 84204 156698
rect 83604 121018 83786 121254
rect 84022 121018 84204 121254
rect 83604 120934 84204 121018
rect 83604 120698 83786 120934
rect 84022 120698 84204 120934
rect 83604 85254 84204 120698
rect 83604 85018 83786 85254
rect 84022 85018 84204 85254
rect 83604 84934 84204 85018
rect 83604 84698 83786 84934
rect 84022 84698 84204 84934
rect 83604 49254 84204 84698
rect 83604 49018 83786 49254
rect 84022 49018 84204 49254
rect 83604 48934 84204 49018
rect 83604 48698 83786 48934
rect 84022 48698 84204 48934
rect 83604 13254 84204 48698
rect 83604 13018 83786 13254
rect 84022 13018 84204 13254
rect 83604 12934 84204 13018
rect 83604 12698 83786 12934
rect 84022 12698 84204 12934
rect 65604 -7022 65786 -6786
rect 66022 -7022 66204 -6786
rect 65604 -7106 66204 -7022
rect 65604 -7342 65786 -7106
rect 66022 -7342 66204 -7106
rect 65604 -7364 66204 -7342
rect 83604 -5866 84204 12698
rect 90804 560454 91404 595898
rect 90804 560218 90986 560454
rect 91222 560218 91404 560454
rect 90804 560134 91404 560218
rect 90804 559898 90986 560134
rect 91222 559898 91404 560134
rect 90804 524454 91404 559898
rect 90804 524218 90986 524454
rect 91222 524218 91404 524454
rect 90804 524134 91404 524218
rect 90804 523898 90986 524134
rect 91222 523898 91404 524134
rect 90804 488454 91404 523898
rect 90804 488218 90986 488454
rect 91222 488218 91404 488454
rect 90804 488134 91404 488218
rect 90804 487898 90986 488134
rect 91222 487898 91404 488134
rect 90804 452454 91404 487898
rect 90804 452218 90986 452454
rect 91222 452218 91404 452454
rect 90804 452134 91404 452218
rect 90804 451898 90986 452134
rect 91222 451898 91404 452134
rect 90804 416454 91404 451898
rect 90804 416218 90986 416454
rect 91222 416218 91404 416454
rect 90804 416134 91404 416218
rect 90804 415898 90986 416134
rect 91222 415898 91404 416134
rect 90804 380454 91404 415898
rect 90804 380218 90986 380454
rect 91222 380218 91404 380454
rect 90804 380134 91404 380218
rect 90804 379898 90986 380134
rect 91222 379898 91404 380134
rect 90804 344454 91404 379898
rect 90804 344218 90986 344454
rect 91222 344218 91404 344454
rect 90804 344134 91404 344218
rect 90804 343898 90986 344134
rect 91222 343898 91404 344134
rect 90804 308454 91404 343898
rect 90804 308218 90986 308454
rect 91222 308218 91404 308454
rect 90804 308134 91404 308218
rect 90804 307898 90986 308134
rect 91222 307898 91404 308134
rect 90804 272454 91404 307898
rect 90804 272218 90986 272454
rect 91222 272218 91404 272454
rect 90804 272134 91404 272218
rect 90804 271898 90986 272134
rect 91222 271898 91404 272134
rect 90804 236454 91404 271898
rect 90804 236218 90986 236454
rect 91222 236218 91404 236454
rect 90804 236134 91404 236218
rect 90804 235898 90986 236134
rect 91222 235898 91404 236134
rect 90804 200454 91404 235898
rect 90804 200218 90986 200454
rect 91222 200218 91404 200454
rect 90804 200134 91404 200218
rect 90804 199898 90986 200134
rect 91222 199898 91404 200134
rect 90804 164454 91404 199898
rect 90804 164218 90986 164454
rect 91222 164218 91404 164454
rect 90804 164134 91404 164218
rect 90804 163898 90986 164134
rect 91222 163898 91404 164134
rect 90804 128454 91404 163898
rect 90804 128218 90986 128454
rect 91222 128218 91404 128454
rect 90804 128134 91404 128218
rect 90804 127898 90986 128134
rect 91222 127898 91404 128134
rect 90804 92454 91404 127898
rect 90804 92218 90986 92454
rect 91222 92218 91404 92454
rect 90804 92134 91404 92218
rect 90804 91898 90986 92134
rect 91222 91898 91404 92134
rect 90804 56454 91404 91898
rect 90804 56218 90986 56454
rect 91222 56218 91404 56454
rect 90804 56134 91404 56218
rect 90804 55898 90986 56134
rect 91222 55898 91404 56134
rect 90804 20454 91404 55898
rect 90804 20218 90986 20454
rect 91222 20218 91404 20454
rect 90804 20134 91404 20218
rect 90804 19898 90986 20134
rect 91222 19898 91404 20134
rect 90804 -1266 91404 19898
rect 90804 -1502 90986 -1266
rect 91222 -1502 91404 -1266
rect 90804 -1586 91404 -1502
rect 90804 -1822 90986 -1586
rect 91222 -1822 91404 -1586
rect 90804 -1844 91404 -1822
rect 94404 672054 95004 707042
rect 94404 671818 94586 672054
rect 94822 671818 95004 672054
rect 94404 671734 95004 671818
rect 94404 671498 94586 671734
rect 94822 671498 95004 671734
rect 94404 636054 95004 671498
rect 94404 635818 94586 636054
rect 94822 635818 95004 636054
rect 94404 635734 95004 635818
rect 94404 635498 94586 635734
rect 94822 635498 95004 635734
rect 94404 600054 95004 635498
rect 94404 599818 94586 600054
rect 94822 599818 95004 600054
rect 94404 599734 95004 599818
rect 94404 599498 94586 599734
rect 94822 599498 95004 599734
rect 94404 564054 95004 599498
rect 94404 563818 94586 564054
rect 94822 563818 95004 564054
rect 94404 563734 95004 563818
rect 94404 563498 94586 563734
rect 94822 563498 95004 563734
rect 94404 528054 95004 563498
rect 94404 527818 94586 528054
rect 94822 527818 95004 528054
rect 94404 527734 95004 527818
rect 94404 527498 94586 527734
rect 94822 527498 95004 527734
rect 94404 492054 95004 527498
rect 94404 491818 94586 492054
rect 94822 491818 95004 492054
rect 94404 491734 95004 491818
rect 94404 491498 94586 491734
rect 94822 491498 95004 491734
rect 94404 456054 95004 491498
rect 94404 455818 94586 456054
rect 94822 455818 95004 456054
rect 94404 455734 95004 455818
rect 94404 455498 94586 455734
rect 94822 455498 95004 455734
rect 94404 420054 95004 455498
rect 94404 419818 94586 420054
rect 94822 419818 95004 420054
rect 94404 419734 95004 419818
rect 94404 419498 94586 419734
rect 94822 419498 95004 419734
rect 94404 384054 95004 419498
rect 94404 383818 94586 384054
rect 94822 383818 95004 384054
rect 94404 383734 95004 383818
rect 94404 383498 94586 383734
rect 94822 383498 95004 383734
rect 94404 348054 95004 383498
rect 94404 347818 94586 348054
rect 94822 347818 95004 348054
rect 94404 347734 95004 347818
rect 94404 347498 94586 347734
rect 94822 347498 95004 347734
rect 94404 312054 95004 347498
rect 94404 311818 94586 312054
rect 94822 311818 95004 312054
rect 94404 311734 95004 311818
rect 94404 311498 94586 311734
rect 94822 311498 95004 311734
rect 94404 276054 95004 311498
rect 94404 275818 94586 276054
rect 94822 275818 95004 276054
rect 94404 275734 95004 275818
rect 94404 275498 94586 275734
rect 94822 275498 95004 275734
rect 94404 240054 95004 275498
rect 94404 239818 94586 240054
rect 94822 239818 95004 240054
rect 94404 239734 95004 239818
rect 94404 239498 94586 239734
rect 94822 239498 95004 239734
rect 94404 204054 95004 239498
rect 94404 203818 94586 204054
rect 94822 203818 95004 204054
rect 94404 203734 95004 203818
rect 94404 203498 94586 203734
rect 94822 203498 95004 203734
rect 94404 168054 95004 203498
rect 94404 167818 94586 168054
rect 94822 167818 95004 168054
rect 94404 167734 95004 167818
rect 94404 167498 94586 167734
rect 94822 167498 95004 167734
rect 94404 132054 95004 167498
rect 94404 131818 94586 132054
rect 94822 131818 95004 132054
rect 94404 131734 95004 131818
rect 94404 131498 94586 131734
rect 94822 131498 95004 131734
rect 94404 96054 95004 131498
rect 94404 95818 94586 96054
rect 94822 95818 95004 96054
rect 94404 95734 95004 95818
rect 94404 95498 94586 95734
rect 94822 95498 95004 95734
rect 94404 60054 95004 95498
rect 94404 59818 94586 60054
rect 94822 59818 95004 60054
rect 94404 59734 95004 59818
rect 94404 59498 94586 59734
rect 94822 59498 95004 59734
rect 94404 24054 95004 59498
rect 94404 23818 94586 24054
rect 94822 23818 95004 24054
rect 94404 23734 95004 23818
rect 94404 23498 94586 23734
rect 94822 23498 95004 23734
rect 94404 -3106 95004 23498
rect 94404 -3342 94586 -3106
rect 94822 -3342 95004 -3106
rect 94404 -3426 95004 -3342
rect 94404 -3662 94586 -3426
rect 94822 -3662 95004 -3426
rect 94404 -3684 95004 -3662
rect 98004 675654 98604 708882
rect 98004 675418 98186 675654
rect 98422 675418 98604 675654
rect 98004 675334 98604 675418
rect 98004 675098 98186 675334
rect 98422 675098 98604 675334
rect 98004 639654 98604 675098
rect 98004 639418 98186 639654
rect 98422 639418 98604 639654
rect 98004 639334 98604 639418
rect 98004 639098 98186 639334
rect 98422 639098 98604 639334
rect 98004 603654 98604 639098
rect 98004 603418 98186 603654
rect 98422 603418 98604 603654
rect 98004 603334 98604 603418
rect 98004 603098 98186 603334
rect 98422 603098 98604 603334
rect 98004 567654 98604 603098
rect 98004 567418 98186 567654
rect 98422 567418 98604 567654
rect 98004 567334 98604 567418
rect 98004 567098 98186 567334
rect 98422 567098 98604 567334
rect 98004 531654 98604 567098
rect 98004 531418 98186 531654
rect 98422 531418 98604 531654
rect 98004 531334 98604 531418
rect 98004 531098 98186 531334
rect 98422 531098 98604 531334
rect 98004 495654 98604 531098
rect 98004 495418 98186 495654
rect 98422 495418 98604 495654
rect 98004 495334 98604 495418
rect 98004 495098 98186 495334
rect 98422 495098 98604 495334
rect 98004 459654 98604 495098
rect 98004 459418 98186 459654
rect 98422 459418 98604 459654
rect 98004 459334 98604 459418
rect 98004 459098 98186 459334
rect 98422 459098 98604 459334
rect 98004 423654 98604 459098
rect 98004 423418 98186 423654
rect 98422 423418 98604 423654
rect 98004 423334 98604 423418
rect 98004 423098 98186 423334
rect 98422 423098 98604 423334
rect 98004 387654 98604 423098
rect 98004 387418 98186 387654
rect 98422 387418 98604 387654
rect 98004 387334 98604 387418
rect 98004 387098 98186 387334
rect 98422 387098 98604 387334
rect 98004 351654 98604 387098
rect 98004 351418 98186 351654
rect 98422 351418 98604 351654
rect 98004 351334 98604 351418
rect 98004 351098 98186 351334
rect 98422 351098 98604 351334
rect 98004 315654 98604 351098
rect 98004 315418 98186 315654
rect 98422 315418 98604 315654
rect 98004 315334 98604 315418
rect 98004 315098 98186 315334
rect 98422 315098 98604 315334
rect 98004 279654 98604 315098
rect 98004 279418 98186 279654
rect 98422 279418 98604 279654
rect 98004 279334 98604 279418
rect 98004 279098 98186 279334
rect 98422 279098 98604 279334
rect 98004 243654 98604 279098
rect 98004 243418 98186 243654
rect 98422 243418 98604 243654
rect 98004 243334 98604 243418
rect 98004 243098 98186 243334
rect 98422 243098 98604 243334
rect 98004 207654 98604 243098
rect 98004 207418 98186 207654
rect 98422 207418 98604 207654
rect 98004 207334 98604 207418
rect 98004 207098 98186 207334
rect 98422 207098 98604 207334
rect 98004 171654 98604 207098
rect 98004 171418 98186 171654
rect 98422 171418 98604 171654
rect 98004 171334 98604 171418
rect 98004 171098 98186 171334
rect 98422 171098 98604 171334
rect 98004 135654 98604 171098
rect 98004 135418 98186 135654
rect 98422 135418 98604 135654
rect 98004 135334 98604 135418
rect 98004 135098 98186 135334
rect 98422 135098 98604 135334
rect 98004 99654 98604 135098
rect 98004 99418 98186 99654
rect 98422 99418 98604 99654
rect 98004 99334 98604 99418
rect 98004 99098 98186 99334
rect 98422 99098 98604 99334
rect 98004 63654 98604 99098
rect 98004 63418 98186 63654
rect 98422 63418 98604 63654
rect 98004 63334 98604 63418
rect 98004 63098 98186 63334
rect 98422 63098 98604 63334
rect 98004 27654 98604 63098
rect 98004 27418 98186 27654
rect 98422 27418 98604 27654
rect 98004 27334 98604 27418
rect 98004 27098 98186 27334
rect 98422 27098 98604 27334
rect 98004 -4946 98604 27098
rect 98004 -5182 98186 -4946
rect 98422 -5182 98604 -4946
rect 98004 -5266 98604 -5182
rect 98004 -5502 98186 -5266
rect 98422 -5502 98604 -5266
rect 98004 -5524 98604 -5502
rect 101604 679254 102204 710722
rect 119604 710358 120204 711300
rect 119604 710122 119786 710358
rect 120022 710122 120204 710358
rect 119604 710038 120204 710122
rect 119604 709802 119786 710038
rect 120022 709802 120204 710038
rect 116004 708518 116604 709460
rect 116004 708282 116186 708518
rect 116422 708282 116604 708518
rect 116004 708198 116604 708282
rect 116004 707962 116186 708198
rect 116422 707962 116604 708198
rect 112404 706678 113004 707620
rect 112404 706442 112586 706678
rect 112822 706442 113004 706678
rect 112404 706358 113004 706442
rect 112404 706122 112586 706358
rect 112822 706122 113004 706358
rect 101604 679018 101786 679254
rect 102022 679018 102204 679254
rect 101604 678934 102204 679018
rect 101604 678698 101786 678934
rect 102022 678698 102204 678934
rect 101604 643254 102204 678698
rect 101604 643018 101786 643254
rect 102022 643018 102204 643254
rect 101604 642934 102204 643018
rect 101604 642698 101786 642934
rect 102022 642698 102204 642934
rect 101604 607254 102204 642698
rect 101604 607018 101786 607254
rect 102022 607018 102204 607254
rect 101604 606934 102204 607018
rect 101604 606698 101786 606934
rect 102022 606698 102204 606934
rect 101604 571254 102204 606698
rect 101604 571018 101786 571254
rect 102022 571018 102204 571254
rect 101604 570934 102204 571018
rect 101604 570698 101786 570934
rect 102022 570698 102204 570934
rect 101604 535254 102204 570698
rect 108804 704838 109404 705780
rect 108804 704602 108986 704838
rect 109222 704602 109404 704838
rect 108804 704518 109404 704602
rect 108804 704282 108986 704518
rect 109222 704282 109404 704518
rect 108804 686454 109404 704282
rect 108804 686218 108986 686454
rect 109222 686218 109404 686454
rect 108804 686134 109404 686218
rect 108804 685898 108986 686134
rect 109222 685898 109404 686134
rect 108804 650454 109404 685898
rect 108804 650218 108986 650454
rect 109222 650218 109404 650454
rect 108804 650134 109404 650218
rect 108804 649898 108986 650134
rect 109222 649898 109404 650134
rect 108804 614454 109404 649898
rect 108804 614218 108986 614454
rect 109222 614218 109404 614454
rect 108804 614134 109404 614218
rect 108804 613898 108986 614134
rect 109222 613898 109404 614134
rect 108804 578454 109404 613898
rect 108804 578218 108986 578454
rect 109222 578218 109404 578454
rect 108804 578134 109404 578218
rect 108804 577898 108986 578134
rect 109222 577898 109404 578134
rect 101604 535018 101786 535254
rect 102022 535018 102204 535254
rect 101604 534934 102204 535018
rect 101604 534698 101786 534934
rect 102022 534698 102204 534934
rect 101604 499254 102204 534698
rect 101604 499018 101786 499254
rect 102022 499018 102204 499254
rect 101604 498934 102204 499018
rect 101604 498698 101786 498934
rect 102022 498698 102204 498934
rect 101604 463254 102204 498698
rect 101604 463018 101786 463254
rect 102022 463018 102204 463254
rect 101604 462934 102204 463018
rect 101604 462698 101786 462934
rect 102022 462698 102204 462934
rect 101604 427254 102204 462698
rect 101604 427018 101786 427254
rect 102022 427018 102204 427254
rect 101604 426934 102204 427018
rect 101604 426698 101786 426934
rect 102022 426698 102204 426934
rect 101604 391254 102204 426698
rect 101604 391018 101786 391254
rect 102022 391018 102204 391254
rect 101604 390934 102204 391018
rect 101604 390698 101786 390934
rect 102022 390698 102204 390934
rect 101604 355254 102204 390698
rect 101604 355018 101786 355254
rect 102022 355018 102204 355254
rect 101604 354934 102204 355018
rect 101604 354698 101786 354934
rect 102022 354698 102204 354934
rect 101604 319254 102204 354698
rect 101604 319018 101786 319254
rect 102022 319018 102204 319254
rect 101604 318934 102204 319018
rect 101604 318698 101786 318934
rect 102022 318698 102204 318934
rect 101604 283254 102204 318698
rect 101604 283018 101786 283254
rect 102022 283018 102204 283254
rect 101604 282934 102204 283018
rect 101604 282698 101786 282934
rect 102022 282698 102204 282934
rect 101604 247254 102204 282698
rect 101604 247018 101786 247254
rect 102022 247018 102204 247254
rect 101604 246934 102204 247018
rect 101604 246698 101786 246934
rect 102022 246698 102204 246934
rect 101604 211254 102204 246698
rect 101604 211018 101786 211254
rect 102022 211018 102204 211254
rect 101604 210934 102204 211018
rect 101604 210698 101786 210934
rect 102022 210698 102204 210934
rect 101604 175254 102204 210698
rect 101604 175018 101786 175254
rect 102022 175018 102204 175254
rect 101604 174934 102204 175018
rect 101604 174698 101786 174934
rect 102022 174698 102204 174934
rect 101604 139254 102204 174698
rect 101604 139018 101786 139254
rect 102022 139018 102204 139254
rect 101604 138934 102204 139018
rect 101604 138698 101786 138934
rect 102022 138698 102204 138934
rect 101604 103254 102204 138698
rect 101604 103018 101786 103254
rect 102022 103018 102204 103254
rect 101604 102934 102204 103018
rect 101604 102698 101786 102934
rect 102022 102698 102204 102934
rect 101604 67254 102204 102698
rect 101604 67018 101786 67254
rect 102022 67018 102204 67254
rect 101604 66934 102204 67018
rect 101604 66698 101786 66934
rect 102022 66698 102204 66934
rect 101604 31254 102204 66698
rect 101604 31018 101786 31254
rect 102022 31018 102204 31254
rect 101604 30934 102204 31018
rect 101604 30698 101786 30934
rect 102022 30698 102204 30934
rect 83604 -6102 83786 -5866
rect 84022 -6102 84204 -5866
rect 83604 -6186 84204 -6102
rect 83604 -6422 83786 -6186
rect 84022 -6422 84204 -6186
rect 83604 -7364 84204 -6422
rect 101604 -6786 102204 30698
rect 108804 542454 109404 577898
rect 112404 690054 113004 706122
rect 112404 689818 112586 690054
rect 112822 689818 113004 690054
rect 112404 689734 113004 689818
rect 112404 689498 112586 689734
rect 112822 689498 113004 689734
rect 112404 654054 113004 689498
rect 112404 653818 112586 654054
rect 112822 653818 113004 654054
rect 112404 653734 113004 653818
rect 112404 653498 112586 653734
rect 112822 653498 113004 653734
rect 112404 618054 113004 653498
rect 112404 617818 112586 618054
rect 112822 617818 113004 618054
rect 112404 617734 113004 617818
rect 112404 617498 112586 617734
rect 112822 617498 113004 617734
rect 112404 582054 113004 617498
rect 112404 581818 112586 582054
rect 112822 581818 113004 582054
rect 112404 581734 113004 581818
rect 112404 581498 112586 581734
rect 112822 581498 113004 581734
rect 108804 542218 108986 542454
rect 109222 542218 109404 542454
rect 108804 542134 109404 542218
rect 108804 541898 108986 542134
rect 109222 541898 109404 542134
rect 108804 506454 109404 541898
rect 108804 506218 108986 506454
rect 109222 506218 109404 506454
rect 108804 506134 109404 506218
rect 108804 505898 108986 506134
rect 109222 505898 109404 506134
rect 108804 470454 109404 505898
rect 108804 470218 108986 470454
rect 109222 470218 109404 470454
rect 108804 470134 109404 470218
rect 108804 469898 108986 470134
rect 109222 469898 109404 470134
rect 108804 434454 109404 469898
rect 108804 434218 108986 434454
rect 109222 434218 109404 434454
rect 108804 434134 109404 434218
rect 108804 433898 108986 434134
rect 109222 433898 109404 434134
rect 108804 398454 109404 433898
rect 108804 398218 108986 398454
rect 109222 398218 109404 398454
rect 108804 398134 109404 398218
rect 108804 397898 108986 398134
rect 109222 397898 109404 398134
rect 108804 362454 109404 397898
rect 108804 362218 108986 362454
rect 109222 362218 109404 362454
rect 108804 362134 109404 362218
rect 108804 361898 108986 362134
rect 109222 361898 109404 362134
rect 108804 326454 109404 361898
rect 108804 326218 108986 326454
rect 109222 326218 109404 326454
rect 108804 326134 109404 326218
rect 108804 325898 108986 326134
rect 109222 325898 109404 326134
rect 108804 290454 109404 325898
rect 108804 290218 108986 290454
rect 109222 290218 109404 290454
rect 108804 290134 109404 290218
rect 108804 289898 108986 290134
rect 109222 289898 109404 290134
rect 108804 254454 109404 289898
rect 108804 254218 108986 254454
rect 109222 254218 109404 254454
rect 108804 254134 109404 254218
rect 108804 253898 108986 254134
rect 109222 253898 109404 254134
rect 108804 218454 109404 253898
rect 108804 218218 108986 218454
rect 109222 218218 109404 218454
rect 108804 218134 109404 218218
rect 108804 217898 108986 218134
rect 109222 217898 109404 218134
rect 108804 182454 109404 217898
rect 108804 182218 108986 182454
rect 109222 182218 109404 182454
rect 108804 182134 109404 182218
rect 108804 181898 108986 182134
rect 109222 181898 109404 182134
rect 108804 146454 109404 181898
rect 108804 146218 108986 146454
rect 109222 146218 109404 146454
rect 108804 146134 109404 146218
rect 108804 145898 108986 146134
rect 109222 145898 109404 146134
rect 108804 110454 109404 145898
rect 108804 110218 108986 110454
rect 109222 110218 109404 110454
rect 108804 110134 109404 110218
rect 108804 109898 108986 110134
rect 109222 109898 109404 110134
rect 108804 74454 109404 109898
rect 108804 74218 108986 74454
rect 109222 74218 109404 74454
rect 108804 74134 109404 74218
rect 108804 73898 108986 74134
rect 109222 73898 109404 74134
rect 108804 38454 109404 73898
rect 108804 38218 108986 38454
rect 109222 38218 109404 38454
rect 108804 38134 109404 38218
rect 108804 37898 108986 38134
rect 109222 37898 109404 38134
rect 108804 2454 109404 37898
rect 108804 2218 108986 2454
rect 109222 2218 109404 2454
rect 108804 2134 109404 2218
rect 108804 1898 108986 2134
rect 109222 1898 109404 2134
rect 108804 -346 109404 1898
rect 108804 -582 108986 -346
rect 109222 -582 109404 -346
rect 108804 -666 109404 -582
rect 108804 -902 108986 -666
rect 109222 -902 109404 -666
rect 108804 -1844 109404 -902
rect 112404 546054 113004 581498
rect 112404 545818 112586 546054
rect 112822 545818 113004 546054
rect 112404 545734 113004 545818
rect 112404 545498 112586 545734
rect 112822 545498 113004 545734
rect 112404 510054 113004 545498
rect 112404 509818 112586 510054
rect 112822 509818 113004 510054
rect 112404 509734 113004 509818
rect 112404 509498 112586 509734
rect 112822 509498 113004 509734
rect 112404 474054 113004 509498
rect 112404 473818 112586 474054
rect 112822 473818 113004 474054
rect 112404 473734 113004 473818
rect 112404 473498 112586 473734
rect 112822 473498 113004 473734
rect 112404 438054 113004 473498
rect 112404 437818 112586 438054
rect 112822 437818 113004 438054
rect 112404 437734 113004 437818
rect 112404 437498 112586 437734
rect 112822 437498 113004 437734
rect 112404 402054 113004 437498
rect 112404 401818 112586 402054
rect 112822 401818 113004 402054
rect 112404 401734 113004 401818
rect 112404 401498 112586 401734
rect 112822 401498 113004 401734
rect 112404 366054 113004 401498
rect 112404 365818 112586 366054
rect 112822 365818 113004 366054
rect 112404 365734 113004 365818
rect 112404 365498 112586 365734
rect 112822 365498 113004 365734
rect 112404 330054 113004 365498
rect 112404 329818 112586 330054
rect 112822 329818 113004 330054
rect 112404 329734 113004 329818
rect 112404 329498 112586 329734
rect 112822 329498 113004 329734
rect 112404 294054 113004 329498
rect 112404 293818 112586 294054
rect 112822 293818 113004 294054
rect 112404 293734 113004 293818
rect 112404 293498 112586 293734
rect 112822 293498 113004 293734
rect 112404 258054 113004 293498
rect 112404 257818 112586 258054
rect 112822 257818 113004 258054
rect 112404 257734 113004 257818
rect 112404 257498 112586 257734
rect 112822 257498 113004 257734
rect 112404 222054 113004 257498
rect 112404 221818 112586 222054
rect 112822 221818 113004 222054
rect 112404 221734 113004 221818
rect 112404 221498 112586 221734
rect 112822 221498 113004 221734
rect 112404 186054 113004 221498
rect 112404 185818 112586 186054
rect 112822 185818 113004 186054
rect 112404 185734 113004 185818
rect 112404 185498 112586 185734
rect 112822 185498 113004 185734
rect 112404 150054 113004 185498
rect 112404 149818 112586 150054
rect 112822 149818 113004 150054
rect 112404 149734 113004 149818
rect 112404 149498 112586 149734
rect 112822 149498 113004 149734
rect 112404 114054 113004 149498
rect 112404 113818 112586 114054
rect 112822 113818 113004 114054
rect 112404 113734 113004 113818
rect 112404 113498 112586 113734
rect 112822 113498 113004 113734
rect 112404 78054 113004 113498
rect 112404 77818 112586 78054
rect 112822 77818 113004 78054
rect 112404 77734 113004 77818
rect 112404 77498 112586 77734
rect 112822 77498 113004 77734
rect 112404 42054 113004 77498
rect 112404 41818 112586 42054
rect 112822 41818 113004 42054
rect 112404 41734 113004 41818
rect 112404 41498 112586 41734
rect 112822 41498 113004 41734
rect 112404 6054 113004 41498
rect 112404 5818 112586 6054
rect 112822 5818 113004 6054
rect 112404 5734 113004 5818
rect 112404 5498 112586 5734
rect 112822 5498 113004 5734
rect 112404 -2186 113004 5498
rect 112404 -2422 112586 -2186
rect 112822 -2422 113004 -2186
rect 112404 -2506 113004 -2422
rect 112404 -2742 112586 -2506
rect 112822 -2742 113004 -2506
rect 112404 -3684 113004 -2742
rect 116004 693654 116604 707962
rect 116004 693418 116186 693654
rect 116422 693418 116604 693654
rect 116004 693334 116604 693418
rect 116004 693098 116186 693334
rect 116422 693098 116604 693334
rect 116004 657654 116604 693098
rect 116004 657418 116186 657654
rect 116422 657418 116604 657654
rect 116004 657334 116604 657418
rect 116004 657098 116186 657334
rect 116422 657098 116604 657334
rect 116004 621654 116604 657098
rect 116004 621418 116186 621654
rect 116422 621418 116604 621654
rect 116004 621334 116604 621418
rect 116004 621098 116186 621334
rect 116422 621098 116604 621334
rect 116004 585654 116604 621098
rect 116004 585418 116186 585654
rect 116422 585418 116604 585654
rect 116004 585334 116604 585418
rect 116004 585098 116186 585334
rect 116422 585098 116604 585334
rect 116004 549654 116604 585098
rect 119604 697254 120204 709802
rect 137604 711278 138204 711300
rect 137604 711042 137786 711278
rect 138022 711042 138204 711278
rect 137604 710958 138204 711042
rect 137604 710722 137786 710958
rect 138022 710722 138204 710958
rect 134004 709438 134604 709460
rect 134004 709202 134186 709438
rect 134422 709202 134604 709438
rect 134004 709118 134604 709202
rect 134004 708882 134186 709118
rect 134422 708882 134604 709118
rect 130404 707598 131004 707620
rect 130404 707362 130586 707598
rect 130822 707362 131004 707598
rect 130404 707278 131004 707362
rect 130404 707042 130586 707278
rect 130822 707042 131004 707278
rect 119604 697018 119786 697254
rect 120022 697018 120204 697254
rect 119604 696934 120204 697018
rect 119604 696698 119786 696934
rect 120022 696698 120204 696934
rect 119604 661254 120204 696698
rect 119604 661018 119786 661254
rect 120022 661018 120204 661254
rect 119604 660934 120204 661018
rect 119604 660698 119786 660934
rect 120022 660698 120204 660934
rect 119604 625254 120204 660698
rect 119604 625018 119786 625254
rect 120022 625018 120204 625254
rect 119604 624934 120204 625018
rect 119604 624698 119786 624934
rect 120022 624698 120204 624934
rect 119604 589254 120204 624698
rect 119604 589018 119786 589254
rect 120022 589018 120204 589254
rect 119604 588934 120204 589018
rect 119604 588698 119786 588934
rect 120022 588698 120204 588934
rect 116004 549418 116186 549654
rect 116422 549418 116604 549654
rect 116004 549334 116604 549418
rect 116004 549098 116186 549334
rect 116422 549098 116604 549334
rect 116004 513654 116604 549098
rect 116004 513418 116186 513654
rect 116422 513418 116604 513654
rect 116004 513334 116604 513418
rect 116004 513098 116186 513334
rect 116422 513098 116604 513334
rect 116004 477654 116604 513098
rect 116004 477418 116186 477654
rect 116422 477418 116604 477654
rect 116004 477334 116604 477418
rect 116004 477098 116186 477334
rect 116422 477098 116604 477334
rect 116004 441654 116604 477098
rect 116004 441418 116186 441654
rect 116422 441418 116604 441654
rect 116004 441334 116604 441418
rect 116004 441098 116186 441334
rect 116422 441098 116604 441334
rect 116004 405654 116604 441098
rect 116004 405418 116186 405654
rect 116422 405418 116604 405654
rect 116004 405334 116604 405418
rect 116004 405098 116186 405334
rect 116422 405098 116604 405334
rect 116004 369654 116604 405098
rect 116004 369418 116186 369654
rect 116422 369418 116604 369654
rect 116004 369334 116604 369418
rect 116004 369098 116186 369334
rect 116422 369098 116604 369334
rect 116004 333654 116604 369098
rect 116004 333418 116186 333654
rect 116422 333418 116604 333654
rect 116004 333334 116604 333418
rect 116004 333098 116186 333334
rect 116422 333098 116604 333334
rect 116004 297654 116604 333098
rect 116004 297418 116186 297654
rect 116422 297418 116604 297654
rect 116004 297334 116604 297418
rect 116004 297098 116186 297334
rect 116422 297098 116604 297334
rect 116004 261654 116604 297098
rect 116004 261418 116186 261654
rect 116422 261418 116604 261654
rect 116004 261334 116604 261418
rect 116004 261098 116186 261334
rect 116422 261098 116604 261334
rect 116004 225654 116604 261098
rect 116004 225418 116186 225654
rect 116422 225418 116604 225654
rect 116004 225334 116604 225418
rect 116004 225098 116186 225334
rect 116422 225098 116604 225334
rect 116004 189654 116604 225098
rect 116004 189418 116186 189654
rect 116422 189418 116604 189654
rect 116004 189334 116604 189418
rect 116004 189098 116186 189334
rect 116422 189098 116604 189334
rect 116004 153654 116604 189098
rect 116004 153418 116186 153654
rect 116422 153418 116604 153654
rect 116004 153334 116604 153418
rect 116004 153098 116186 153334
rect 116422 153098 116604 153334
rect 116004 117654 116604 153098
rect 116004 117418 116186 117654
rect 116422 117418 116604 117654
rect 116004 117334 116604 117418
rect 116004 117098 116186 117334
rect 116422 117098 116604 117334
rect 116004 81654 116604 117098
rect 116004 81418 116186 81654
rect 116422 81418 116604 81654
rect 116004 81334 116604 81418
rect 116004 81098 116186 81334
rect 116422 81098 116604 81334
rect 116004 45654 116604 81098
rect 116004 45418 116186 45654
rect 116422 45418 116604 45654
rect 116004 45334 116604 45418
rect 116004 45098 116186 45334
rect 116422 45098 116604 45334
rect 116004 9654 116604 45098
rect 116004 9418 116186 9654
rect 116422 9418 116604 9654
rect 116004 9334 116604 9418
rect 116004 9098 116186 9334
rect 116422 9098 116604 9334
rect 116004 -4026 116604 9098
rect 116004 -4262 116186 -4026
rect 116422 -4262 116604 -4026
rect 116004 -4346 116604 -4262
rect 116004 -4582 116186 -4346
rect 116422 -4582 116604 -4346
rect 116004 -5524 116604 -4582
rect 119604 553254 120204 588698
rect 126804 705758 127404 705780
rect 126804 705522 126986 705758
rect 127222 705522 127404 705758
rect 126804 705438 127404 705522
rect 126804 705202 126986 705438
rect 127222 705202 127404 705438
rect 126804 668454 127404 705202
rect 126804 668218 126986 668454
rect 127222 668218 127404 668454
rect 126804 668134 127404 668218
rect 126804 667898 126986 668134
rect 127222 667898 127404 668134
rect 126804 632454 127404 667898
rect 126804 632218 126986 632454
rect 127222 632218 127404 632454
rect 126804 632134 127404 632218
rect 126804 631898 126986 632134
rect 127222 631898 127404 632134
rect 126804 596454 127404 631898
rect 126804 596218 126986 596454
rect 127222 596218 127404 596454
rect 126804 596134 127404 596218
rect 126804 595898 126986 596134
rect 127222 595898 127404 596134
rect 120766 561373 120826 562582
rect 120763 561372 120829 561373
rect 120763 561308 120764 561372
rect 120828 561308 120829 561372
rect 120763 561307 120829 561308
rect 119604 553018 119786 553254
rect 120022 553018 120204 553254
rect 119604 552934 120204 553018
rect 119604 552698 119786 552934
rect 120022 552698 120204 552934
rect 119604 517254 120204 552698
rect 119604 517018 119786 517254
rect 120022 517018 120204 517254
rect 119604 516934 120204 517018
rect 119604 516698 119786 516934
rect 120022 516698 120204 516934
rect 119604 481254 120204 516698
rect 119604 481018 119786 481254
rect 120022 481018 120204 481254
rect 119604 480934 120204 481018
rect 119604 480698 119786 480934
rect 120022 480698 120204 480934
rect 119604 445254 120204 480698
rect 119604 445018 119786 445254
rect 120022 445018 120204 445254
rect 119604 444934 120204 445018
rect 119604 444698 119786 444934
rect 120022 444698 120204 444934
rect 119604 409254 120204 444698
rect 119604 409018 119786 409254
rect 120022 409018 120204 409254
rect 119604 408934 120204 409018
rect 119604 408698 119786 408934
rect 120022 408698 120204 408934
rect 119604 373254 120204 408698
rect 119604 373018 119786 373254
rect 120022 373018 120204 373254
rect 119604 372934 120204 373018
rect 119604 372698 119786 372934
rect 120022 372698 120204 372934
rect 119604 337254 120204 372698
rect 119604 337018 119786 337254
rect 120022 337018 120204 337254
rect 119604 336934 120204 337018
rect 119604 336698 119786 336934
rect 120022 336698 120204 336934
rect 119604 301254 120204 336698
rect 119604 301018 119786 301254
rect 120022 301018 120204 301254
rect 119604 300934 120204 301018
rect 119604 300698 119786 300934
rect 120022 300698 120204 300934
rect 119604 265254 120204 300698
rect 119604 265018 119786 265254
rect 120022 265018 120204 265254
rect 119604 264934 120204 265018
rect 119604 264698 119786 264934
rect 120022 264698 120204 264934
rect 119604 229254 120204 264698
rect 119604 229018 119786 229254
rect 120022 229018 120204 229254
rect 119604 228934 120204 229018
rect 119604 228698 119786 228934
rect 120022 228698 120204 228934
rect 119604 193254 120204 228698
rect 119604 193018 119786 193254
rect 120022 193018 120204 193254
rect 119604 192934 120204 193018
rect 119604 192698 119786 192934
rect 120022 192698 120204 192934
rect 119604 157254 120204 192698
rect 119604 157018 119786 157254
rect 120022 157018 120204 157254
rect 119604 156934 120204 157018
rect 119604 156698 119786 156934
rect 120022 156698 120204 156934
rect 119604 121254 120204 156698
rect 119604 121018 119786 121254
rect 120022 121018 120204 121254
rect 119604 120934 120204 121018
rect 119604 120698 119786 120934
rect 120022 120698 120204 120934
rect 119604 85254 120204 120698
rect 119604 85018 119786 85254
rect 120022 85018 120204 85254
rect 119604 84934 120204 85018
rect 119604 84698 119786 84934
rect 120022 84698 120204 84934
rect 119604 49254 120204 84698
rect 119604 49018 119786 49254
rect 120022 49018 120204 49254
rect 119604 48934 120204 49018
rect 119604 48698 119786 48934
rect 120022 48698 120204 48934
rect 119604 13254 120204 48698
rect 119604 13018 119786 13254
rect 120022 13018 120204 13254
rect 119604 12934 120204 13018
rect 119604 12698 119786 12934
rect 120022 12698 120204 12934
rect 101604 -7022 101786 -6786
rect 102022 -7022 102204 -6786
rect 101604 -7106 102204 -7022
rect 101604 -7342 101786 -7106
rect 102022 -7342 102204 -7106
rect 101604 -7364 102204 -7342
rect 119604 -5866 120204 12698
rect 126804 560454 127404 595898
rect 126804 560218 126986 560454
rect 127222 560218 127404 560454
rect 126804 560134 127404 560218
rect 126804 559898 126986 560134
rect 127222 559898 127404 560134
rect 126804 524454 127404 559898
rect 126804 524218 126986 524454
rect 127222 524218 127404 524454
rect 126804 524134 127404 524218
rect 126804 523898 126986 524134
rect 127222 523898 127404 524134
rect 126804 488454 127404 523898
rect 126804 488218 126986 488454
rect 127222 488218 127404 488454
rect 126804 488134 127404 488218
rect 126804 487898 126986 488134
rect 127222 487898 127404 488134
rect 126804 452454 127404 487898
rect 126804 452218 126986 452454
rect 127222 452218 127404 452454
rect 126804 452134 127404 452218
rect 126804 451898 126986 452134
rect 127222 451898 127404 452134
rect 126804 416454 127404 451898
rect 126804 416218 126986 416454
rect 127222 416218 127404 416454
rect 126804 416134 127404 416218
rect 126804 415898 126986 416134
rect 127222 415898 127404 416134
rect 126804 380454 127404 415898
rect 126804 380218 126986 380454
rect 127222 380218 127404 380454
rect 126804 380134 127404 380218
rect 126804 379898 126986 380134
rect 127222 379898 127404 380134
rect 126804 344454 127404 379898
rect 126804 344218 126986 344454
rect 127222 344218 127404 344454
rect 126804 344134 127404 344218
rect 126804 343898 126986 344134
rect 127222 343898 127404 344134
rect 126804 308454 127404 343898
rect 126804 308218 126986 308454
rect 127222 308218 127404 308454
rect 126804 308134 127404 308218
rect 126804 307898 126986 308134
rect 127222 307898 127404 308134
rect 126804 272454 127404 307898
rect 126804 272218 126986 272454
rect 127222 272218 127404 272454
rect 126804 272134 127404 272218
rect 126804 271898 126986 272134
rect 127222 271898 127404 272134
rect 126804 236454 127404 271898
rect 126804 236218 126986 236454
rect 127222 236218 127404 236454
rect 126804 236134 127404 236218
rect 126804 235898 126986 236134
rect 127222 235898 127404 236134
rect 126804 200454 127404 235898
rect 126804 200218 126986 200454
rect 127222 200218 127404 200454
rect 126804 200134 127404 200218
rect 126804 199898 126986 200134
rect 127222 199898 127404 200134
rect 126804 164454 127404 199898
rect 126804 164218 126986 164454
rect 127222 164218 127404 164454
rect 126804 164134 127404 164218
rect 126804 163898 126986 164134
rect 127222 163898 127404 164134
rect 126804 128454 127404 163898
rect 126804 128218 126986 128454
rect 127222 128218 127404 128454
rect 126804 128134 127404 128218
rect 126804 127898 126986 128134
rect 127222 127898 127404 128134
rect 126804 92454 127404 127898
rect 126804 92218 126986 92454
rect 127222 92218 127404 92454
rect 126804 92134 127404 92218
rect 126804 91898 126986 92134
rect 127222 91898 127404 92134
rect 126804 56454 127404 91898
rect 126804 56218 126986 56454
rect 127222 56218 127404 56454
rect 126804 56134 127404 56218
rect 126804 55898 126986 56134
rect 127222 55898 127404 56134
rect 126804 20454 127404 55898
rect 126804 20218 126986 20454
rect 127222 20218 127404 20454
rect 126804 20134 127404 20218
rect 126804 19898 126986 20134
rect 127222 19898 127404 20134
rect 126804 -1266 127404 19898
rect 126804 -1502 126986 -1266
rect 127222 -1502 127404 -1266
rect 126804 -1586 127404 -1502
rect 126804 -1822 126986 -1586
rect 127222 -1822 127404 -1586
rect 126804 -1844 127404 -1822
rect 130404 672054 131004 707042
rect 130404 671818 130586 672054
rect 130822 671818 131004 672054
rect 130404 671734 131004 671818
rect 130404 671498 130586 671734
rect 130822 671498 131004 671734
rect 130404 636054 131004 671498
rect 130404 635818 130586 636054
rect 130822 635818 131004 636054
rect 130404 635734 131004 635818
rect 130404 635498 130586 635734
rect 130822 635498 131004 635734
rect 130404 600054 131004 635498
rect 130404 599818 130586 600054
rect 130822 599818 131004 600054
rect 130404 599734 131004 599818
rect 130404 599498 130586 599734
rect 130822 599498 131004 599734
rect 130404 564054 131004 599498
rect 130404 563818 130586 564054
rect 130822 563818 131004 564054
rect 130404 563734 131004 563818
rect 130404 563498 130586 563734
rect 130822 563498 131004 563734
rect 130404 528054 131004 563498
rect 130404 527818 130586 528054
rect 130822 527818 131004 528054
rect 130404 527734 131004 527818
rect 130404 527498 130586 527734
rect 130822 527498 131004 527734
rect 130404 492054 131004 527498
rect 130404 491818 130586 492054
rect 130822 491818 131004 492054
rect 130404 491734 131004 491818
rect 130404 491498 130586 491734
rect 130822 491498 131004 491734
rect 130404 456054 131004 491498
rect 130404 455818 130586 456054
rect 130822 455818 131004 456054
rect 130404 455734 131004 455818
rect 130404 455498 130586 455734
rect 130822 455498 131004 455734
rect 130404 420054 131004 455498
rect 130404 419818 130586 420054
rect 130822 419818 131004 420054
rect 130404 419734 131004 419818
rect 130404 419498 130586 419734
rect 130822 419498 131004 419734
rect 130404 384054 131004 419498
rect 130404 383818 130586 384054
rect 130822 383818 131004 384054
rect 130404 383734 131004 383818
rect 130404 383498 130586 383734
rect 130822 383498 131004 383734
rect 130404 348054 131004 383498
rect 130404 347818 130586 348054
rect 130822 347818 131004 348054
rect 130404 347734 131004 347818
rect 130404 347498 130586 347734
rect 130822 347498 131004 347734
rect 130404 312054 131004 347498
rect 130404 311818 130586 312054
rect 130822 311818 131004 312054
rect 130404 311734 131004 311818
rect 130404 311498 130586 311734
rect 130822 311498 131004 311734
rect 130404 276054 131004 311498
rect 130404 275818 130586 276054
rect 130822 275818 131004 276054
rect 130404 275734 131004 275818
rect 130404 275498 130586 275734
rect 130822 275498 131004 275734
rect 130404 240054 131004 275498
rect 130404 239818 130586 240054
rect 130822 239818 131004 240054
rect 130404 239734 131004 239818
rect 130404 239498 130586 239734
rect 130822 239498 131004 239734
rect 130404 204054 131004 239498
rect 130404 203818 130586 204054
rect 130822 203818 131004 204054
rect 130404 203734 131004 203818
rect 130404 203498 130586 203734
rect 130822 203498 131004 203734
rect 130404 168054 131004 203498
rect 130404 167818 130586 168054
rect 130822 167818 131004 168054
rect 130404 167734 131004 167818
rect 130404 167498 130586 167734
rect 130822 167498 131004 167734
rect 130404 132054 131004 167498
rect 130404 131818 130586 132054
rect 130822 131818 131004 132054
rect 130404 131734 131004 131818
rect 130404 131498 130586 131734
rect 130822 131498 131004 131734
rect 130404 96054 131004 131498
rect 130404 95818 130586 96054
rect 130822 95818 131004 96054
rect 130404 95734 131004 95818
rect 130404 95498 130586 95734
rect 130822 95498 131004 95734
rect 130404 60054 131004 95498
rect 130404 59818 130586 60054
rect 130822 59818 131004 60054
rect 130404 59734 131004 59818
rect 130404 59498 130586 59734
rect 130822 59498 131004 59734
rect 130404 24054 131004 59498
rect 130404 23818 130586 24054
rect 130822 23818 131004 24054
rect 130404 23734 131004 23818
rect 130404 23498 130586 23734
rect 130822 23498 131004 23734
rect 130404 -3106 131004 23498
rect 130404 -3342 130586 -3106
rect 130822 -3342 131004 -3106
rect 130404 -3426 131004 -3342
rect 130404 -3662 130586 -3426
rect 130822 -3662 131004 -3426
rect 130404 -3684 131004 -3662
rect 134004 675654 134604 708882
rect 134004 675418 134186 675654
rect 134422 675418 134604 675654
rect 134004 675334 134604 675418
rect 134004 675098 134186 675334
rect 134422 675098 134604 675334
rect 134004 639654 134604 675098
rect 134004 639418 134186 639654
rect 134422 639418 134604 639654
rect 134004 639334 134604 639418
rect 134004 639098 134186 639334
rect 134422 639098 134604 639334
rect 134004 603654 134604 639098
rect 134004 603418 134186 603654
rect 134422 603418 134604 603654
rect 134004 603334 134604 603418
rect 134004 603098 134186 603334
rect 134422 603098 134604 603334
rect 134004 567654 134604 603098
rect 134004 567418 134186 567654
rect 134422 567418 134604 567654
rect 134004 567334 134604 567418
rect 134004 567098 134186 567334
rect 134422 567098 134604 567334
rect 134004 531654 134604 567098
rect 137604 679254 138204 710722
rect 155604 710358 156204 711300
rect 155604 710122 155786 710358
rect 156022 710122 156204 710358
rect 155604 710038 156204 710122
rect 155604 709802 155786 710038
rect 156022 709802 156204 710038
rect 152004 708518 152604 709460
rect 152004 708282 152186 708518
rect 152422 708282 152604 708518
rect 152004 708198 152604 708282
rect 152004 707962 152186 708198
rect 152422 707962 152604 708198
rect 148404 706678 149004 707620
rect 148404 706442 148586 706678
rect 148822 706442 149004 706678
rect 148404 706358 149004 706442
rect 148404 706122 148586 706358
rect 148822 706122 149004 706358
rect 137604 679018 137786 679254
rect 138022 679018 138204 679254
rect 137604 678934 138204 679018
rect 137604 678698 137786 678934
rect 138022 678698 138204 678934
rect 137604 643254 138204 678698
rect 137604 643018 137786 643254
rect 138022 643018 138204 643254
rect 137604 642934 138204 643018
rect 137604 642698 137786 642934
rect 138022 642698 138204 642934
rect 137604 607254 138204 642698
rect 137604 607018 137786 607254
rect 138022 607018 138204 607254
rect 137604 606934 138204 607018
rect 137604 606698 137786 606934
rect 138022 606698 138204 606934
rect 137604 571254 138204 606698
rect 137604 571018 137786 571254
rect 138022 571018 138204 571254
rect 137604 570934 138204 571018
rect 137604 570698 137786 570934
rect 138022 570698 138204 570934
rect 135115 562732 135181 562733
rect 135115 562668 135116 562732
rect 135180 562668 135181 562732
rect 135115 562667 135181 562668
rect 135118 561458 135178 562667
rect 134004 531418 134186 531654
rect 134422 531418 134604 531654
rect 134004 531334 134604 531418
rect 134004 531098 134186 531334
rect 134422 531098 134604 531334
rect 134004 495654 134604 531098
rect 134004 495418 134186 495654
rect 134422 495418 134604 495654
rect 134004 495334 134604 495418
rect 134004 495098 134186 495334
rect 134422 495098 134604 495334
rect 134004 459654 134604 495098
rect 134004 459418 134186 459654
rect 134422 459418 134604 459654
rect 134004 459334 134604 459418
rect 134004 459098 134186 459334
rect 134422 459098 134604 459334
rect 134004 423654 134604 459098
rect 134004 423418 134186 423654
rect 134422 423418 134604 423654
rect 134004 423334 134604 423418
rect 134004 423098 134186 423334
rect 134422 423098 134604 423334
rect 134004 387654 134604 423098
rect 134004 387418 134186 387654
rect 134422 387418 134604 387654
rect 134004 387334 134604 387418
rect 134004 387098 134186 387334
rect 134422 387098 134604 387334
rect 134004 351654 134604 387098
rect 134004 351418 134186 351654
rect 134422 351418 134604 351654
rect 134004 351334 134604 351418
rect 134004 351098 134186 351334
rect 134422 351098 134604 351334
rect 134004 315654 134604 351098
rect 134004 315418 134186 315654
rect 134422 315418 134604 315654
rect 134004 315334 134604 315418
rect 134004 315098 134186 315334
rect 134422 315098 134604 315334
rect 134004 279654 134604 315098
rect 134004 279418 134186 279654
rect 134422 279418 134604 279654
rect 134004 279334 134604 279418
rect 134004 279098 134186 279334
rect 134422 279098 134604 279334
rect 134004 243654 134604 279098
rect 134004 243418 134186 243654
rect 134422 243418 134604 243654
rect 134004 243334 134604 243418
rect 134004 243098 134186 243334
rect 134422 243098 134604 243334
rect 134004 207654 134604 243098
rect 134004 207418 134186 207654
rect 134422 207418 134604 207654
rect 134004 207334 134604 207418
rect 134004 207098 134186 207334
rect 134422 207098 134604 207334
rect 134004 171654 134604 207098
rect 134004 171418 134186 171654
rect 134422 171418 134604 171654
rect 134004 171334 134604 171418
rect 134004 171098 134186 171334
rect 134422 171098 134604 171334
rect 134004 135654 134604 171098
rect 134004 135418 134186 135654
rect 134422 135418 134604 135654
rect 134004 135334 134604 135418
rect 134004 135098 134186 135334
rect 134422 135098 134604 135334
rect 134004 99654 134604 135098
rect 134004 99418 134186 99654
rect 134422 99418 134604 99654
rect 134004 99334 134604 99418
rect 134004 99098 134186 99334
rect 134422 99098 134604 99334
rect 134004 63654 134604 99098
rect 134004 63418 134186 63654
rect 134422 63418 134604 63654
rect 134004 63334 134604 63418
rect 134004 63098 134186 63334
rect 134422 63098 134604 63334
rect 134004 27654 134604 63098
rect 134004 27418 134186 27654
rect 134422 27418 134604 27654
rect 134004 27334 134604 27418
rect 134004 27098 134186 27334
rect 134422 27098 134604 27334
rect 134004 -4946 134604 27098
rect 134004 -5182 134186 -4946
rect 134422 -5182 134604 -4946
rect 134004 -5266 134604 -5182
rect 134004 -5502 134186 -5266
rect 134422 -5502 134604 -5266
rect 134004 -5524 134604 -5502
rect 137604 535254 138204 570698
rect 144804 704838 145404 705780
rect 144804 704602 144986 704838
rect 145222 704602 145404 704838
rect 144804 704518 145404 704602
rect 144804 704282 144986 704518
rect 145222 704282 145404 704518
rect 144804 686454 145404 704282
rect 144804 686218 144986 686454
rect 145222 686218 145404 686454
rect 144804 686134 145404 686218
rect 144804 685898 144986 686134
rect 145222 685898 145404 686134
rect 144804 650454 145404 685898
rect 144804 650218 144986 650454
rect 145222 650218 145404 650454
rect 144804 650134 145404 650218
rect 144804 649898 144986 650134
rect 145222 649898 145404 650134
rect 144804 614454 145404 649898
rect 144804 614218 144986 614454
rect 145222 614218 145404 614454
rect 144804 614134 145404 614218
rect 144804 613898 144986 614134
rect 145222 613898 145404 614134
rect 144804 578454 145404 613898
rect 144804 578218 144986 578454
rect 145222 578218 145404 578454
rect 144804 578134 145404 578218
rect 144804 577898 144986 578134
rect 145222 577898 145404 578134
rect 140086 561373 140146 562582
rect 140083 561372 140149 561373
rect 140083 561308 140084 561372
rect 140148 561308 140149 561372
rect 140083 561307 140149 561308
rect 137604 535018 137786 535254
rect 138022 535018 138204 535254
rect 137604 534934 138204 535018
rect 137604 534698 137786 534934
rect 138022 534698 138204 534934
rect 137604 499254 138204 534698
rect 137604 499018 137786 499254
rect 138022 499018 138204 499254
rect 137604 498934 138204 499018
rect 137604 498698 137786 498934
rect 138022 498698 138204 498934
rect 137604 463254 138204 498698
rect 137604 463018 137786 463254
rect 138022 463018 138204 463254
rect 137604 462934 138204 463018
rect 137604 462698 137786 462934
rect 138022 462698 138204 462934
rect 137604 427254 138204 462698
rect 137604 427018 137786 427254
rect 138022 427018 138204 427254
rect 137604 426934 138204 427018
rect 137604 426698 137786 426934
rect 138022 426698 138204 426934
rect 137604 391254 138204 426698
rect 137604 391018 137786 391254
rect 138022 391018 138204 391254
rect 137604 390934 138204 391018
rect 137604 390698 137786 390934
rect 138022 390698 138204 390934
rect 137604 355254 138204 390698
rect 137604 355018 137786 355254
rect 138022 355018 138204 355254
rect 137604 354934 138204 355018
rect 137604 354698 137786 354934
rect 138022 354698 138204 354934
rect 137604 319254 138204 354698
rect 137604 319018 137786 319254
rect 138022 319018 138204 319254
rect 137604 318934 138204 319018
rect 137604 318698 137786 318934
rect 138022 318698 138204 318934
rect 137604 283254 138204 318698
rect 137604 283018 137786 283254
rect 138022 283018 138204 283254
rect 137604 282934 138204 283018
rect 137604 282698 137786 282934
rect 138022 282698 138204 282934
rect 137604 247254 138204 282698
rect 137604 247018 137786 247254
rect 138022 247018 138204 247254
rect 137604 246934 138204 247018
rect 137604 246698 137786 246934
rect 138022 246698 138204 246934
rect 137604 211254 138204 246698
rect 137604 211018 137786 211254
rect 138022 211018 138204 211254
rect 137604 210934 138204 211018
rect 137604 210698 137786 210934
rect 138022 210698 138204 210934
rect 137604 175254 138204 210698
rect 137604 175018 137786 175254
rect 138022 175018 138204 175254
rect 137604 174934 138204 175018
rect 137604 174698 137786 174934
rect 138022 174698 138204 174934
rect 137604 139254 138204 174698
rect 137604 139018 137786 139254
rect 138022 139018 138204 139254
rect 137604 138934 138204 139018
rect 137604 138698 137786 138934
rect 138022 138698 138204 138934
rect 137604 103254 138204 138698
rect 137604 103018 137786 103254
rect 138022 103018 138204 103254
rect 137604 102934 138204 103018
rect 137604 102698 137786 102934
rect 138022 102698 138204 102934
rect 137604 67254 138204 102698
rect 137604 67018 137786 67254
rect 138022 67018 138204 67254
rect 137604 66934 138204 67018
rect 137604 66698 137786 66934
rect 138022 66698 138204 66934
rect 137604 31254 138204 66698
rect 137604 31018 137786 31254
rect 138022 31018 138204 31254
rect 137604 30934 138204 31018
rect 137604 30698 137786 30934
rect 138022 30698 138204 30934
rect 119604 -6102 119786 -5866
rect 120022 -6102 120204 -5866
rect 119604 -6186 120204 -6102
rect 119604 -6422 119786 -6186
rect 120022 -6422 120204 -6186
rect 119604 -7364 120204 -6422
rect 137604 -6786 138204 30698
rect 144804 542454 145404 577898
rect 148404 690054 149004 706122
rect 148404 689818 148586 690054
rect 148822 689818 149004 690054
rect 148404 689734 149004 689818
rect 148404 689498 148586 689734
rect 148822 689498 149004 689734
rect 148404 654054 149004 689498
rect 148404 653818 148586 654054
rect 148822 653818 149004 654054
rect 148404 653734 149004 653818
rect 148404 653498 148586 653734
rect 148822 653498 149004 653734
rect 148404 618054 149004 653498
rect 148404 617818 148586 618054
rect 148822 617818 149004 618054
rect 148404 617734 149004 617818
rect 148404 617498 148586 617734
rect 148822 617498 149004 617734
rect 148404 582054 149004 617498
rect 148404 581818 148586 582054
rect 148822 581818 149004 582054
rect 148404 581734 149004 581818
rect 148404 581498 148586 581734
rect 148822 581498 149004 581734
rect 144804 542218 144986 542454
rect 145222 542218 145404 542454
rect 144804 542134 145404 542218
rect 144804 541898 144986 542134
rect 145222 541898 145404 542134
rect 144804 506454 145404 541898
rect 144804 506218 144986 506454
rect 145222 506218 145404 506454
rect 144804 506134 145404 506218
rect 144804 505898 144986 506134
rect 145222 505898 145404 506134
rect 144804 470454 145404 505898
rect 144804 470218 144986 470454
rect 145222 470218 145404 470454
rect 144804 470134 145404 470218
rect 144804 469898 144986 470134
rect 145222 469898 145404 470134
rect 144804 434454 145404 469898
rect 144804 434218 144986 434454
rect 145222 434218 145404 434454
rect 144804 434134 145404 434218
rect 144804 433898 144986 434134
rect 145222 433898 145404 434134
rect 144804 398454 145404 433898
rect 144804 398218 144986 398454
rect 145222 398218 145404 398454
rect 144804 398134 145404 398218
rect 144804 397898 144986 398134
rect 145222 397898 145404 398134
rect 144804 362454 145404 397898
rect 144804 362218 144986 362454
rect 145222 362218 145404 362454
rect 144804 362134 145404 362218
rect 144804 361898 144986 362134
rect 145222 361898 145404 362134
rect 144804 326454 145404 361898
rect 144804 326218 144986 326454
rect 145222 326218 145404 326454
rect 144804 326134 145404 326218
rect 144804 325898 144986 326134
rect 145222 325898 145404 326134
rect 144804 290454 145404 325898
rect 144804 290218 144986 290454
rect 145222 290218 145404 290454
rect 144804 290134 145404 290218
rect 144804 289898 144986 290134
rect 145222 289898 145404 290134
rect 144804 254454 145404 289898
rect 144804 254218 144986 254454
rect 145222 254218 145404 254454
rect 144804 254134 145404 254218
rect 144804 253898 144986 254134
rect 145222 253898 145404 254134
rect 144804 218454 145404 253898
rect 144804 218218 144986 218454
rect 145222 218218 145404 218454
rect 144804 218134 145404 218218
rect 144804 217898 144986 218134
rect 145222 217898 145404 218134
rect 144804 182454 145404 217898
rect 144804 182218 144986 182454
rect 145222 182218 145404 182454
rect 144804 182134 145404 182218
rect 144804 181898 144986 182134
rect 145222 181898 145404 182134
rect 144804 146454 145404 181898
rect 144804 146218 144986 146454
rect 145222 146218 145404 146454
rect 144804 146134 145404 146218
rect 144804 145898 144986 146134
rect 145222 145898 145404 146134
rect 144804 110454 145404 145898
rect 144804 110218 144986 110454
rect 145222 110218 145404 110454
rect 144804 110134 145404 110218
rect 144804 109898 144986 110134
rect 145222 109898 145404 110134
rect 144804 74454 145404 109898
rect 144804 74218 144986 74454
rect 145222 74218 145404 74454
rect 144804 74134 145404 74218
rect 144804 73898 144986 74134
rect 145222 73898 145404 74134
rect 144804 38454 145404 73898
rect 144804 38218 144986 38454
rect 145222 38218 145404 38454
rect 144804 38134 145404 38218
rect 144804 37898 144986 38134
rect 145222 37898 145404 38134
rect 144804 2454 145404 37898
rect 144804 2218 144986 2454
rect 145222 2218 145404 2454
rect 144804 2134 145404 2218
rect 144804 1898 144986 2134
rect 145222 1898 145404 2134
rect 144804 -346 145404 1898
rect 144804 -582 144986 -346
rect 145222 -582 145404 -346
rect 144804 -666 145404 -582
rect 144804 -902 144986 -666
rect 145222 -902 145404 -666
rect 144804 -1844 145404 -902
rect 148404 546054 149004 581498
rect 148404 545818 148586 546054
rect 148822 545818 149004 546054
rect 148404 545734 149004 545818
rect 148404 545498 148586 545734
rect 148822 545498 149004 545734
rect 148404 510054 149004 545498
rect 148404 509818 148586 510054
rect 148822 509818 149004 510054
rect 148404 509734 149004 509818
rect 148404 509498 148586 509734
rect 148822 509498 149004 509734
rect 148404 474054 149004 509498
rect 148404 473818 148586 474054
rect 148822 473818 149004 474054
rect 148404 473734 149004 473818
rect 148404 473498 148586 473734
rect 148822 473498 149004 473734
rect 148404 438054 149004 473498
rect 148404 437818 148586 438054
rect 148822 437818 149004 438054
rect 148404 437734 149004 437818
rect 148404 437498 148586 437734
rect 148822 437498 149004 437734
rect 148404 402054 149004 437498
rect 148404 401818 148586 402054
rect 148822 401818 149004 402054
rect 148404 401734 149004 401818
rect 148404 401498 148586 401734
rect 148822 401498 149004 401734
rect 148404 366054 149004 401498
rect 148404 365818 148586 366054
rect 148822 365818 149004 366054
rect 148404 365734 149004 365818
rect 148404 365498 148586 365734
rect 148822 365498 149004 365734
rect 148404 330054 149004 365498
rect 148404 329818 148586 330054
rect 148822 329818 149004 330054
rect 148404 329734 149004 329818
rect 148404 329498 148586 329734
rect 148822 329498 149004 329734
rect 148404 294054 149004 329498
rect 148404 293818 148586 294054
rect 148822 293818 149004 294054
rect 148404 293734 149004 293818
rect 148404 293498 148586 293734
rect 148822 293498 149004 293734
rect 148404 258054 149004 293498
rect 148404 257818 148586 258054
rect 148822 257818 149004 258054
rect 148404 257734 149004 257818
rect 148404 257498 148586 257734
rect 148822 257498 149004 257734
rect 148404 222054 149004 257498
rect 148404 221818 148586 222054
rect 148822 221818 149004 222054
rect 148404 221734 149004 221818
rect 148404 221498 148586 221734
rect 148822 221498 149004 221734
rect 148404 186054 149004 221498
rect 148404 185818 148586 186054
rect 148822 185818 149004 186054
rect 148404 185734 149004 185818
rect 148404 185498 148586 185734
rect 148822 185498 149004 185734
rect 148404 150054 149004 185498
rect 148404 149818 148586 150054
rect 148822 149818 149004 150054
rect 148404 149734 149004 149818
rect 148404 149498 148586 149734
rect 148822 149498 149004 149734
rect 148404 114054 149004 149498
rect 148404 113818 148586 114054
rect 148822 113818 149004 114054
rect 148404 113734 149004 113818
rect 148404 113498 148586 113734
rect 148822 113498 149004 113734
rect 148404 78054 149004 113498
rect 148404 77818 148586 78054
rect 148822 77818 149004 78054
rect 148404 77734 149004 77818
rect 148404 77498 148586 77734
rect 148822 77498 149004 77734
rect 148404 42054 149004 77498
rect 148404 41818 148586 42054
rect 148822 41818 149004 42054
rect 148404 41734 149004 41818
rect 148404 41498 148586 41734
rect 148822 41498 149004 41734
rect 148404 6054 149004 41498
rect 148404 5818 148586 6054
rect 148822 5818 149004 6054
rect 148404 5734 149004 5818
rect 148404 5498 148586 5734
rect 148822 5498 149004 5734
rect 148404 -2186 149004 5498
rect 148404 -2422 148586 -2186
rect 148822 -2422 149004 -2186
rect 148404 -2506 149004 -2422
rect 148404 -2742 148586 -2506
rect 148822 -2742 149004 -2506
rect 148404 -3684 149004 -2742
rect 152004 693654 152604 707962
rect 152004 693418 152186 693654
rect 152422 693418 152604 693654
rect 152004 693334 152604 693418
rect 152004 693098 152186 693334
rect 152422 693098 152604 693334
rect 152004 657654 152604 693098
rect 152004 657418 152186 657654
rect 152422 657418 152604 657654
rect 152004 657334 152604 657418
rect 152004 657098 152186 657334
rect 152422 657098 152604 657334
rect 152004 621654 152604 657098
rect 152004 621418 152186 621654
rect 152422 621418 152604 621654
rect 152004 621334 152604 621418
rect 152004 621098 152186 621334
rect 152422 621098 152604 621334
rect 152004 585654 152604 621098
rect 152004 585418 152186 585654
rect 152422 585418 152604 585654
rect 152004 585334 152604 585418
rect 152004 585098 152186 585334
rect 152422 585098 152604 585334
rect 152004 549654 152604 585098
rect 155604 697254 156204 709802
rect 173604 711278 174204 711300
rect 173604 711042 173786 711278
rect 174022 711042 174204 711278
rect 173604 710958 174204 711042
rect 173604 710722 173786 710958
rect 174022 710722 174204 710958
rect 170004 709438 170604 709460
rect 170004 709202 170186 709438
rect 170422 709202 170604 709438
rect 170004 709118 170604 709202
rect 170004 708882 170186 709118
rect 170422 708882 170604 709118
rect 166404 707598 167004 707620
rect 166404 707362 166586 707598
rect 166822 707362 167004 707598
rect 166404 707278 167004 707362
rect 166404 707042 166586 707278
rect 166822 707042 167004 707278
rect 155604 697018 155786 697254
rect 156022 697018 156204 697254
rect 155604 696934 156204 697018
rect 155604 696698 155786 696934
rect 156022 696698 156204 696934
rect 155604 661254 156204 696698
rect 155604 661018 155786 661254
rect 156022 661018 156204 661254
rect 155604 660934 156204 661018
rect 155604 660698 155786 660934
rect 156022 660698 156204 660934
rect 155604 625254 156204 660698
rect 155604 625018 155786 625254
rect 156022 625018 156204 625254
rect 155604 624934 156204 625018
rect 155604 624698 155786 624934
rect 156022 624698 156204 624934
rect 155604 589254 156204 624698
rect 155604 589018 155786 589254
rect 156022 589018 156204 589254
rect 155604 588934 156204 589018
rect 155604 588698 155786 588934
rect 156022 588698 156204 588934
rect 152004 549418 152186 549654
rect 152422 549418 152604 549654
rect 152004 549334 152604 549418
rect 152004 549098 152186 549334
rect 152422 549098 152604 549334
rect 152004 513654 152604 549098
rect 152004 513418 152186 513654
rect 152422 513418 152604 513654
rect 152004 513334 152604 513418
rect 152004 513098 152186 513334
rect 152422 513098 152604 513334
rect 152004 477654 152604 513098
rect 152004 477418 152186 477654
rect 152422 477418 152604 477654
rect 152004 477334 152604 477418
rect 152004 477098 152186 477334
rect 152422 477098 152604 477334
rect 152004 441654 152604 477098
rect 152004 441418 152186 441654
rect 152422 441418 152604 441654
rect 152004 441334 152604 441418
rect 152004 441098 152186 441334
rect 152422 441098 152604 441334
rect 152004 405654 152604 441098
rect 152004 405418 152186 405654
rect 152422 405418 152604 405654
rect 152004 405334 152604 405418
rect 152004 405098 152186 405334
rect 152422 405098 152604 405334
rect 152004 369654 152604 405098
rect 152004 369418 152186 369654
rect 152422 369418 152604 369654
rect 152004 369334 152604 369418
rect 152004 369098 152186 369334
rect 152422 369098 152604 369334
rect 152004 333654 152604 369098
rect 152004 333418 152186 333654
rect 152422 333418 152604 333654
rect 152004 333334 152604 333418
rect 152004 333098 152186 333334
rect 152422 333098 152604 333334
rect 152004 297654 152604 333098
rect 152004 297418 152186 297654
rect 152422 297418 152604 297654
rect 152004 297334 152604 297418
rect 152004 297098 152186 297334
rect 152422 297098 152604 297334
rect 152004 261654 152604 297098
rect 152004 261418 152186 261654
rect 152422 261418 152604 261654
rect 152004 261334 152604 261418
rect 152004 261098 152186 261334
rect 152422 261098 152604 261334
rect 152004 225654 152604 261098
rect 152004 225418 152186 225654
rect 152422 225418 152604 225654
rect 152004 225334 152604 225418
rect 152004 225098 152186 225334
rect 152422 225098 152604 225334
rect 152004 189654 152604 225098
rect 152004 189418 152186 189654
rect 152422 189418 152604 189654
rect 152004 189334 152604 189418
rect 152004 189098 152186 189334
rect 152422 189098 152604 189334
rect 152004 153654 152604 189098
rect 152004 153418 152186 153654
rect 152422 153418 152604 153654
rect 152004 153334 152604 153418
rect 152004 153098 152186 153334
rect 152422 153098 152604 153334
rect 152004 117654 152604 153098
rect 152004 117418 152186 117654
rect 152422 117418 152604 117654
rect 152004 117334 152604 117418
rect 152004 117098 152186 117334
rect 152422 117098 152604 117334
rect 152004 81654 152604 117098
rect 152004 81418 152186 81654
rect 152422 81418 152604 81654
rect 152004 81334 152604 81418
rect 152004 81098 152186 81334
rect 152422 81098 152604 81334
rect 152004 45654 152604 81098
rect 152004 45418 152186 45654
rect 152422 45418 152604 45654
rect 152004 45334 152604 45418
rect 152004 45098 152186 45334
rect 152422 45098 152604 45334
rect 152004 9654 152604 45098
rect 152004 9418 152186 9654
rect 152422 9418 152604 9654
rect 152004 9334 152604 9418
rect 152004 9098 152186 9334
rect 152422 9098 152604 9334
rect 152004 -4026 152604 9098
rect 152004 -4262 152186 -4026
rect 152422 -4262 152604 -4026
rect 152004 -4346 152604 -4262
rect 152004 -4582 152186 -4346
rect 152422 -4582 152604 -4346
rect 152004 -5524 152604 -4582
rect 155604 553254 156204 588698
rect 162804 705758 163404 705780
rect 162804 705522 162986 705758
rect 163222 705522 163404 705758
rect 162804 705438 163404 705522
rect 162804 705202 162986 705438
rect 163222 705202 163404 705438
rect 162804 668454 163404 705202
rect 162804 668218 162986 668454
rect 163222 668218 163404 668454
rect 162804 668134 163404 668218
rect 162804 667898 162986 668134
rect 163222 667898 163404 668134
rect 162804 632454 163404 667898
rect 162804 632218 162986 632454
rect 163222 632218 163404 632454
rect 162804 632134 163404 632218
rect 162804 631898 162986 632134
rect 163222 631898 163404 632134
rect 162804 596454 163404 631898
rect 162804 596218 162986 596454
rect 163222 596218 163404 596454
rect 162804 596134 163404 596218
rect 162804 595898 162986 596134
rect 163222 595898 163404 596134
rect 159406 561373 159466 562582
rect 159403 561372 159469 561373
rect 159403 561308 159404 561372
rect 159468 561308 159469 561372
rect 159403 561307 159469 561308
rect 155604 553018 155786 553254
rect 156022 553018 156204 553254
rect 155604 552934 156204 553018
rect 155604 552698 155786 552934
rect 156022 552698 156204 552934
rect 155604 517254 156204 552698
rect 155604 517018 155786 517254
rect 156022 517018 156204 517254
rect 155604 516934 156204 517018
rect 155604 516698 155786 516934
rect 156022 516698 156204 516934
rect 155604 481254 156204 516698
rect 155604 481018 155786 481254
rect 156022 481018 156204 481254
rect 155604 480934 156204 481018
rect 155604 480698 155786 480934
rect 156022 480698 156204 480934
rect 155604 445254 156204 480698
rect 155604 445018 155786 445254
rect 156022 445018 156204 445254
rect 155604 444934 156204 445018
rect 155604 444698 155786 444934
rect 156022 444698 156204 444934
rect 155604 409254 156204 444698
rect 155604 409018 155786 409254
rect 156022 409018 156204 409254
rect 155604 408934 156204 409018
rect 155604 408698 155786 408934
rect 156022 408698 156204 408934
rect 155604 373254 156204 408698
rect 155604 373018 155786 373254
rect 156022 373018 156204 373254
rect 155604 372934 156204 373018
rect 155604 372698 155786 372934
rect 156022 372698 156204 372934
rect 155604 337254 156204 372698
rect 155604 337018 155786 337254
rect 156022 337018 156204 337254
rect 155604 336934 156204 337018
rect 155604 336698 155786 336934
rect 156022 336698 156204 336934
rect 155604 301254 156204 336698
rect 155604 301018 155786 301254
rect 156022 301018 156204 301254
rect 155604 300934 156204 301018
rect 155604 300698 155786 300934
rect 156022 300698 156204 300934
rect 155604 265254 156204 300698
rect 155604 265018 155786 265254
rect 156022 265018 156204 265254
rect 155604 264934 156204 265018
rect 155604 264698 155786 264934
rect 156022 264698 156204 264934
rect 155604 229254 156204 264698
rect 155604 229018 155786 229254
rect 156022 229018 156204 229254
rect 155604 228934 156204 229018
rect 155604 228698 155786 228934
rect 156022 228698 156204 228934
rect 155604 193254 156204 228698
rect 155604 193018 155786 193254
rect 156022 193018 156204 193254
rect 155604 192934 156204 193018
rect 155604 192698 155786 192934
rect 156022 192698 156204 192934
rect 155604 157254 156204 192698
rect 155604 157018 155786 157254
rect 156022 157018 156204 157254
rect 155604 156934 156204 157018
rect 155604 156698 155786 156934
rect 156022 156698 156204 156934
rect 155604 121254 156204 156698
rect 155604 121018 155786 121254
rect 156022 121018 156204 121254
rect 155604 120934 156204 121018
rect 155604 120698 155786 120934
rect 156022 120698 156204 120934
rect 155604 85254 156204 120698
rect 155604 85018 155786 85254
rect 156022 85018 156204 85254
rect 155604 84934 156204 85018
rect 155604 84698 155786 84934
rect 156022 84698 156204 84934
rect 155604 49254 156204 84698
rect 155604 49018 155786 49254
rect 156022 49018 156204 49254
rect 155604 48934 156204 49018
rect 155604 48698 155786 48934
rect 156022 48698 156204 48934
rect 155604 13254 156204 48698
rect 155604 13018 155786 13254
rect 156022 13018 156204 13254
rect 155604 12934 156204 13018
rect 155604 12698 155786 12934
rect 156022 12698 156204 12934
rect 137604 -7022 137786 -6786
rect 138022 -7022 138204 -6786
rect 137604 -7106 138204 -7022
rect 137604 -7342 137786 -7106
rect 138022 -7342 138204 -7106
rect 137604 -7364 138204 -7342
rect 155604 -5866 156204 12698
rect 162804 560454 163404 595898
rect 166404 672054 167004 707042
rect 166404 671818 166586 672054
rect 166822 671818 167004 672054
rect 166404 671734 167004 671818
rect 166404 671498 166586 671734
rect 166822 671498 167004 671734
rect 166404 636054 167004 671498
rect 166404 635818 166586 636054
rect 166822 635818 167004 636054
rect 166404 635734 167004 635818
rect 166404 635498 166586 635734
rect 166822 635498 167004 635734
rect 166404 600054 167004 635498
rect 166404 599818 166586 600054
rect 166822 599818 167004 600054
rect 166404 599734 167004 599818
rect 166404 599498 166586 599734
rect 166822 599498 167004 599734
rect 166404 564054 167004 599498
rect 166404 563818 166586 564054
rect 166822 563818 167004 564054
rect 166404 563734 167004 563818
rect 166404 563498 166586 563734
rect 166822 563498 167004 563734
rect 162804 560218 162986 560454
rect 163222 560218 163404 560454
rect 162804 560134 163404 560218
rect 162804 559898 162986 560134
rect 163222 559898 163404 560134
rect 162804 524454 163404 559898
rect 162804 524218 162986 524454
rect 163222 524218 163404 524454
rect 162804 524134 163404 524218
rect 162804 523898 162986 524134
rect 163222 523898 163404 524134
rect 162804 488454 163404 523898
rect 162804 488218 162986 488454
rect 163222 488218 163404 488454
rect 162804 488134 163404 488218
rect 162804 487898 162986 488134
rect 163222 487898 163404 488134
rect 162804 452454 163404 487898
rect 162804 452218 162986 452454
rect 163222 452218 163404 452454
rect 162804 452134 163404 452218
rect 162804 451898 162986 452134
rect 163222 451898 163404 452134
rect 162804 416454 163404 451898
rect 162804 416218 162986 416454
rect 163222 416218 163404 416454
rect 162804 416134 163404 416218
rect 162804 415898 162986 416134
rect 163222 415898 163404 416134
rect 162804 380454 163404 415898
rect 162804 380218 162986 380454
rect 163222 380218 163404 380454
rect 162804 380134 163404 380218
rect 162804 379898 162986 380134
rect 163222 379898 163404 380134
rect 162804 344454 163404 379898
rect 162804 344218 162986 344454
rect 163222 344218 163404 344454
rect 162804 344134 163404 344218
rect 162804 343898 162986 344134
rect 163222 343898 163404 344134
rect 162804 308454 163404 343898
rect 162804 308218 162986 308454
rect 163222 308218 163404 308454
rect 162804 308134 163404 308218
rect 162804 307898 162986 308134
rect 163222 307898 163404 308134
rect 162804 272454 163404 307898
rect 162804 272218 162986 272454
rect 163222 272218 163404 272454
rect 162804 272134 163404 272218
rect 162804 271898 162986 272134
rect 163222 271898 163404 272134
rect 162804 236454 163404 271898
rect 162804 236218 162986 236454
rect 163222 236218 163404 236454
rect 162804 236134 163404 236218
rect 162804 235898 162986 236134
rect 163222 235898 163404 236134
rect 162804 200454 163404 235898
rect 162804 200218 162986 200454
rect 163222 200218 163404 200454
rect 162804 200134 163404 200218
rect 162804 199898 162986 200134
rect 163222 199898 163404 200134
rect 162804 164454 163404 199898
rect 162804 164218 162986 164454
rect 163222 164218 163404 164454
rect 162804 164134 163404 164218
rect 162804 163898 162986 164134
rect 163222 163898 163404 164134
rect 162804 128454 163404 163898
rect 162804 128218 162986 128454
rect 163222 128218 163404 128454
rect 162804 128134 163404 128218
rect 162804 127898 162986 128134
rect 163222 127898 163404 128134
rect 162804 92454 163404 127898
rect 162804 92218 162986 92454
rect 163222 92218 163404 92454
rect 162804 92134 163404 92218
rect 162804 91898 162986 92134
rect 163222 91898 163404 92134
rect 162804 56454 163404 91898
rect 162804 56218 162986 56454
rect 163222 56218 163404 56454
rect 162804 56134 163404 56218
rect 162804 55898 162986 56134
rect 163222 55898 163404 56134
rect 162804 20454 163404 55898
rect 162804 20218 162986 20454
rect 163222 20218 163404 20454
rect 162804 20134 163404 20218
rect 162804 19898 162986 20134
rect 163222 19898 163404 20134
rect 162804 -1266 163404 19898
rect 162804 -1502 162986 -1266
rect 163222 -1502 163404 -1266
rect 162804 -1586 163404 -1502
rect 162804 -1822 162986 -1586
rect 163222 -1822 163404 -1586
rect 162804 -1844 163404 -1822
rect 166404 528054 167004 563498
rect 170004 675654 170604 708882
rect 170004 675418 170186 675654
rect 170422 675418 170604 675654
rect 170004 675334 170604 675418
rect 170004 675098 170186 675334
rect 170422 675098 170604 675334
rect 170004 639654 170604 675098
rect 170004 639418 170186 639654
rect 170422 639418 170604 639654
rect 170004 639334 170604 639418
rect 170004 639098 170186 639334
rect 170422 639098 170604 639334
rect 170004 603654 170604 639098
rect 170004 603418 170186 603654
rect 170422 603418 170604 603654
rect 170004 603334 170604 603418
rect 170004 603098 170186 603334
rect 170422 603098 170604 603334
rect 170004 567654 170604 603098
rect 170004 567418 170186 567654
rect 170422 567418 170604 567654
rect 170004 567334 170604 567418
rect 170004 567098 170186 567334
rect 170422 567098 170604 567334
rect 166404 527818 166586 528054
rect 166822 527818 167004 528054
rect 166404 527734 167004 527818
rect 166404 527498 166586 527734
rect 166822 527498 167004 527734
rect 166404 492054 167004 527498
rect 166404 491818 166586 492054
rect 166822 491818 167004 492054
rect 166404 491734 167004 491818
rect 166404 491498 166586 491734
rect 166822 491498 167004 491734
rect 166404 456054 167004 491498
rect 166404 455818 166586 456054
rect 166822 455818 167004 456054
rect 166404 455734 167004 455818
rect 166404 455498 166586 455734
rect 166822 455498 167004 455734
rect 166404 420054 167004 455498
rect 166404 419818 166586 420054
rect 166822 419818 167004 420054
rect 166404 419734 167004 419818
rect 166404 419498 166586 419734
rect 166822 419498 167004 419734
rect 166404 384054 167004 419498
rect 166404 383818 166586 384054
rect 166822 383818 167004 384054
rect 166404 383734 167004 383818
rect 166404 383498 166586 383734
rect 166822 383498 167004 383734
rect 166404 348054 167004 383498
rect 166404 347818 166586 348054
rect 166822 347818 167004 348054
rect 166404 347734 167004 347818
rect 166404 347498 166586 347734
rect 166822 347498 167004 347734
rect 166404 312054 167004 347498
rect 166404 311818 166586 312054
rect 166822 311818 167004 312054
rect 166404 311734 167004 311818
rect 166404 311498 166586 311734
rect 166822 311498 167004 311734
rect 166404 276054 167004 311498
rect 166404 275818 166586 276054
rect 166822 275818 167004 276054
rect 166404 275734 167004 275818
rect 166404 275498 166586 275734
rect 166822 275498 167004 275734
rect 166404 240054 167004 275498
rect 166404 239818 166586 240054
rect 166822 239818 167004 240054
rect 166404 239734 167004 239818
rect 166404 239498 166586 239734
rect 166822 239498 167004 239734
rect 166404 204054 167004 239498
rect 166404 203818 166586 204054
rect 166822 203818 167004 204054
rect 166404 203734 167004 203818
rect 166404 203498 166586 203734
rect 166822 203498 167004 203734
rect 166404 168054 167004 203498
rect 166404 167818 166586 168054
rect 166822 167818 167004 168054
rect 166404 167734 167004 167818
rect 166404 167498 166586 167734
rect 166822 167498 167004 167734
rect 166404 132054 167004 167498
rect 166404 131818 166586 132054
rect 166822 131818 167004 132054
rect 166404 131734 167004 131818
rect 166404 131498 166586 131734
rect 166822 131498 167004 131734
rect 166404 96054 167004 131498
rect 166404 95818 166586 96054
rect 166822 95818 167004 96054
rect 166404 95734 167004 95818
rect 166404 95498 166586 95734
rect 166822 95498 167004 95734
rect 166404 60054 167004 95498
rect 166404 59818 166586 60054
rect 166822 59818 167004 60054
rect 166404 59734 167004 59818
rect 166404 59498 166586 59734
rect 166822 59498 167004 59734
rect 166404 24054 167004 59498
rect 166404 23818 166586 24054
rect 166822 23818 167004 24054
rect 166404 23734 167004 23818
rect 166404 23498 166586 23734
rect 166822 23498 167004 23734
rect 166404 -3106 167004 23498
rect 166404 -3342 166586 -3106
rect 166822 -3342 167004 -3106
rect 166404 -3426 167004 -3342
rect 166404 -3662 166586 -3426
rect 166822 -3662 167004 -3426
rect 166404 -3684 167004 -3662
rect 170004 531654 170604 567098
rect 170004 531418 170186 531654
rect 170422 531418 170604 531654
rect 170004 531334 170604 531418
rect 170004 531098 170186 531334
rect 170422 531098 170604 531334
rect 170004 495654 170604 531098
rect 170004 495418 170186 495654
rect 170422 495418 170604 495654
rect 170004 495334 170604 495418
rect 170004 495098 170186 495334
rect 170422 495098 170604 495334
rect 170004 459654 170604 495098
rect 170004 459418 170186 459654
rect 170422 459418 170604 459654
rect 170004 459334 170604 459418
rect 170004 459098 170186 459334
rect 170422 459098 170604 459334
rect 170004 423654 170604 459098
rect 170004 423418 170186 423654
rect 170422 423418 170604 423654
rect 170004 423334 170604 423418
rect 170004 423098 170186 423334
rect 170422 423098 170604 423334
rect 170004 387654 170604 423098
rect 170004 387418 170186 387654
rect 170422 387418 170604 387654
rect 170004 387334 170604 387418
rect 170004 387098 170186 387334
rect 170422 387098 170604 387334
rect 170004 351654 170604 387098
rect 170004 351418 170186 351654
rect 170422 351418 170604 351654
rect 170004 351334 170604 351418
rect 170004 351098 170186 351334
rect 170422 351098 170604 351334
rect 170004 315654 170604 351098
rect 170004 315418 170186 315654
rect 170422 315418 170604 315654
rect 170004 315334 170604 315418
rect 170004 315098 170186 315334
rect 170422 315098 170604 315334
rect 170004 279654 170604 315098
rect 170004 279418 170186 279654
rect 170422 279418 170604 279654
rect 170004 279334 170604 279418
rect 170004 279098 170186 279334
rect 170422 279098 170604 279334
rect 170004 243654 170604 279098
rect 170004 243418 170186 243654
rect 170422 243418 170604 243654
rect 170004 243334 170604 243418
rect 170004 243098 170186 243334
rect 170422 243098 170604 243334
rect 170004 207654 170604 243098
rect 170004 207418 170186 207654
rect 170422 207418 170604 207654
rect 170004 207334 170604 207418
rect 170004 207098 170186 207334
rect 170422 207098 170604 207334
rect 170004 171654 170604 207098
rect 170004 171418 170186 171654
rect 170422 171418 170604 171654
rect 170004 171334 170604 171418
rect 170004 171098 170186 171334
rect 170422 171098 170604 171334
rect 170004 135654 170604 171098
rect 170004 135418 170186 135654
rect 170422 135418 170604 135654
rect 170004 135334 170604 135418
rect 170004 135098 170186 135334
rect 170422 135098 170604 135334
rect 170004 99654 170604 135098
rect 170004 99418 170186 99654
rect 170422 99418 170604 99654
rect 170004 99334 170604 99418
rect 170004 99098 170186 99334
rect 170422 99098 170604 99334
rect 170004 63654 170604 99098
rect 170004 63418 170186 63654
rect 170422 63418 170604 63654
rect 170004 63334 170604 63418
rect 170004 63098 170186 63334
rect 170422 63098 170604 63334
rect 170004 27654 170604 63098
rect 170004 27418 170186 27654
rect 170422 27418 170604 27654
rect 170004 27334 170604 27418
rect 170004 27098 170186 27334
rect 170422 27098 170604 27334
rect 170004 -4946 170604 27098
rect 170004 -5182 170186 -4946
rect 170422 -5182 170604 -4946
rect 170004 -5266 170604 -5182
rect 170004 -5502 170186 -5266
rect 170422 -5502 170604 -5266
rect 170004 -5524 170604 -5502
rect 173604 679254 174204 710722
rect 191604 710358 192204 711300
rect 191604 710122 191786 710358
rect 192022 710122 192204 710358
rect 191604 710038 192204 710122
rect 191604 709802 191786 710038
rect 192022 709802 192204 710038
rect 188004 708518 188604 709460
rect 188004 708282 188186 708518
rect 188422 708282 188604 708518
rect 188004 708198 188604 708282
rect 188004 707962 188186 708198
rect 188422 707962 188604 708198
rect 184404 706678 185004 707620
rect 184404 706442 184586 706678
rect 184822 706442 185004 706678
rect 184404 706358 185004 706442
rect 184404 706122 184586 706358
rect 184822 706122 185004 706358
rect 173604 679018 173786 679254
rect 174022 679018 174204 679254
rect 173604 678934 174204 679018
rect 173604 678698 173786 678934
rect 174022 678698 174204 678934
rect 173604 643254 174204 678698
rect 173604 643018 173786 643254
rect 174022 643018 174204 643254
rect 173604 642934 174204 643018
rect 173604 642698 173786 642934
rect 174022 642698 174204 642934
rect 173604 607254 174204 642698
rect 173604 607018 173786 607254
rect 174022 607018 174204 607254
rect 173604 606934 174204 607018
rect 173604 606698 173786 606934
rect 174022 606698 174204 606934
rect 173604 571254 174204 606698
rect 173604 571018 173786 571254
rect 174022 571018 174204 571254
rect 173604 570934 174204 571018
rect 173604 570698 173786 570934
rect 174022 570698 174204 570934
rect 173604 535254 174204 570698
rect 180804 704838 181404 705780
rect 180804 704602 180986 704838
rect 181222 704602 181404 704838
rect 180804 704518 181404 704602
rect 180804 704282 180986 704518
rect 181222 704282 181404 704518
rect 180804 686454 181404 704282
rect 180804 686218 180986 686454
rect 181222 686218 181404 686454
rect 180804 686134 181404 686218
rect 180804 685898 180986 686134
rect 181222 685898 181404 686134
rect 180804 650454 181404 685898
rect 180804 650218 180986 650454
rect 181222 650218 181404 650454
rect 180804 650134 181404 650218
rect 180804 649898 180986 650134
rect 181222 649898 181404 650134
rect 180804 614454 181404 649898
rect 180804 614218 180986 614454
rect 181222 614218 181404 614454
rect 180804 614134 181404 614218
rect 180804 613898 180986 614134
rect 181222 613898 181404 614134
rect 180804 578454 181404 613898
rect 180804 578218 180986 578454
rect 181222 578218 181404 578454
rect 180804 578134 181404 578218
rect 180804 577898 180986 578134
rect 181222 577898 181404 578134
rect 178726 561373 178786 562582
rect 178723 561372 178789 561373
rect 178723 561308 178724 561372
rect 178788 561308 178789 561372
rect 178723 561307 178789 561308
rect 173604 535018 173786 535254
rect 174022 535018 174204 535254
rect 173604 534934 174204 535018
rect 173604 534698 173786 534934
rect 174022 534698 174204 534934
rect 173604 499254 174204 534698
rect 173604 499018 173786 499254
rect 174022 499018 174204 499254
rect 173604 498934 174204 499018
rect 173604 498698 173786 498934
rect 174022 498698 174204 498934
rect 173604 463254 174204 498698
rect 173604 463018 173786 463254
rect 174022 463018 174204 463254
rect 173604 462934 174204 463018
rect 173604 462698 173786 462934
rect 174022 462698 174204 462934
rect 173604 427254 174204 462698
rect 173604 427018 173786 427254
rect 174022 427018 174204 427254
rect 173604 426934 174204 427018
rect 173604 426698 173786 426934
rect 174022 426698 174204 426934
rect 173604 391254 174204 426698
rect 173604 391018 173786 391254
rect 174022 391018 174204 391254
rect 173604 390934 174204 391018
rect 173604 390698 173786 390934
rect 174022 390698 174204 390934
rect 173604 355254 174204 390698
rect 173604 355018 173786 355254
rect 174022 355018 174204 355254
rect 173604 354934 174204 355018
rect 173604 354698 173786 354934
rect 174022 354698 174204 354934
rect 173604 319254 174204 354698
rect 173604 319018 173786 319254
rect 174022 319018 174204 319254
rect 173604 318934 174204 319018
rect 173604 318698 173786 318934
rect 174022 318698 174204 318934
rect 173604 283254 174204 318698
rect 173604 283018 173786 283254
rect 174022 283018 174204 283254
rect 173604 282934 174204 283018
rect 173604 282698 173786 282934
rect 174022 282698 174204 282934
rect 173604 247254 174204 282698
rect 173604 247018 173786 247254
rect 174022 247018 174204 247254
rect 173604 246934 174204 247018
rect 173604 246698 173786 246934
rect 174022 246698 174204 246934
rect 173604 211254 174204 246698
rect 173604 211018 173786 211254
rect 174022 211018 174204 211254
rect 173604 210934 174204 211018
rect 173604 210698 173786 210934
rect 174022 210698 174204 210934
rect 173604 175254 174204 210698
rect 173604 175018 173786 175254
rect 174022 175018 174204 175254
rect 173604 174934 174204 175018
rect 173604 174698 173786 174934
rect 174022 174698 174204 174934
rect 173604 139254 174204 174698
rect 173604 139018 173786 139254
rect 174022 139018 174204 139254
rect 173604 138934 174204 139018
rect 173604 138698 173786 138934
rect 174022 138698 174204 138934
rect 173604 103254 174204 138698
rect 173604 103018 173786 103254
rect 174022 103018 174204 103254
rect 173604 102934 174204 103018
rect 173604 102698 173786 102934
rect 174022 102698 174204 102934
rect 173604 67254 174204 102698
rect 173604 67018 173786 67254
rect 174022 67018 174204 67254
rect 173604 66934 174204 67018
rect 173604 66698 173786 66934
rect 174022 66698 174204 66934
rect 173604 31254 174204 66698
rect 173604 31018 173786 31254
rect 174022 31018 174204 31254
rect 173604 30934 174204 31018
rect 173604 30698 173786 30934
rect 174022 30698 174204 30934
rect 155604 -6102 155786 -5866
rect 156022 -6102 156204 -5866
rect 155604 -6186 156204 -6102
rect 155604 -6422 155786 -6186
rect 156022 -6422 156204 -6186
rect 155604 -7364 156204 -6422
rect 173604 -6786 174204 30698
rect 180804 542454 181404 577898
rect 184404 690054 185004 706122
rect 184404 689818 184586 690054
rect 184822 689818 185004 690054
rect 184404 689734 185004 689818
rect 184404 689498 184586 689734
rect 184822 689498 185004 689734
rect 184404 654054 185004 689498
rect 184404 653818 184586 654054
rect 184822 653818 185004 654054
rect 184404 653734 185004 653818
rect 184404 653498 184586 653734
rect 184822 653498 185004 653734
rect 184404 618054 185004 653498
rect 184404 617818 184586 618054
rect 184822 617818 185004 618054
rect 184404 617734 185004 617818
rect 184404 617498 184586 617734
rect 184822 617498 185004 617734
rect 184404 582054 185004 617498
rect 184404 581818 184586 582054
rect 184822 581818 185004 582054
rect 184404 581734 185004 581818
rect 184404 581498 184586 581734
rect 184822 581498 185004 581734
rect 180804 542218 180986 542454
rect 181222 542218 181404 542454
rect 180804 542134 181404 542218
rect 180804 541898 180986 542134
rect 181222 541898 181404 542134
rect 180804 506454 181404 541898
rect 180804 506218 180986 506454
rect 181222 506218 181404 506454
rect 180804 506134 181404 506218
rect 180804 505898 180986 506134
rect 181222 505898 181404 506134
rect 180804 470454 181404 505898
rect 180804 470218 180986 470454
rect 181222 470218 181404 470454
rect 180804 470134 181404 470218
rect 180804 469898 180986 470134
rect 181222 469898 181404 470134
rect 180804 434454 181404 469898
rect 180804 434218 180986 434454
rect 181222 434218 181404 434454
rect 180804 434134 181404 434218
rect 180804 433898 180986 434134
rect 181222 433898 181404 434134
rect 180804 398454 181404 433898
rect 180804 398218 180986 398454
rect 181222 398218 181404 398454
rect 180804 398134 181404 398218
rect 180804 397898 180986 398134
rect 181222 397898 181404 398134
rect 180804 362454 181404 397898
rect 180804 362218 180986 362454
rect 181222 362218 181404 362454
rect 180804 362134 181404 362218
rect 180804 361898 180986 362134
rect 181222 361898 181404 362134
rect 180804 326454 181404 361898
rect 180804 326218 180986 326454
rect 181222 326218 181404 326454
rect 180804 326134 181404 326218
rect 180804 325898 180986 326134
rect 181222 325898 181404 326134
rect 180804 290454 181404 325898
rect 180804 290218 180986 290454
rect 181222 290218 181404 290454
rect 180804 290134 181404 290218
rect 180804 289898 180986 290134
rect 181222 289898 181404 290134
rect 180804 254454 181404 289898
rect 180804 254218 180986 254454
rect 181222 254218 181404 254454
rect 180804 254134 181404 254218
rect 180804 253898 180986 254134
rect 181222 253898 181404 254134
rect 180804 218454 181404 253898
rect 180804 218218 180986 218454
rect 181222 218218 181404 218454
rect 180804 218134 181404 218218
rect 180804 217898 180986 218134
rect 181222 217898 181404 218134
rect 180804 182454 181404 217898
rect 180804 182218 180986 182454
rect 181222 182218 181404 182454
rect 180804 182134 181404 182218
rect 180804 181898 180986 182134
rect 181222 181898 181404 182134
rect 180804 146454 181404 181898
rect 180804 146218 180986 146454
rect 181222 146218 181404 146454
rect 180804 146134 181404 146218
rect 180804 145898 180986 146134
rect 181222 145898 181404 146134
rect 180804 110454 181404 145898
rect 180804 110218 180986 110454
rect 181222 110218 181404 110454
rect 180804 110134 181404 110218
rect 180804 109898 180986 110134
rect 181222 109898 181404 110134
rect 180804 74454 181404 109898
rect 180804 74218 180986 74454
rect 181222 74218 181404 74454
rect 180804 74134 181404 74218
rect 180804 73898 180986 74134
rect 181222 73898 181404 74134
rect 180804 38454 181404 73898
rect 180804 38218 180986 38454
rect 181222 38218 181404 38454
rect 180804 38134 181404 38218
rect 180804 37898 180986 38134
rect 181222 37898 181404 38134
rect 180804 2454 181404 37898
rect 180804 2218 180986 2454
rect 181222 2218 181404 2454
rect 180804 2134 181404 2218
rect 180804 1898 180986 2134
rect 181222 1898 181404 2134
rect 180804 -346 181404 1898
rect 180804 -582 180986 -346
rect 181222 -582 181404 -346
rect 180804 -666 181404 -582
rect 180804 -902 180986 -666
rect 181222 -902 181404 -666
rect 180804 -1844 181404 -902
rect 184404 546054 185004 581498
rect 184404 545818 184586 546054
rect 184822 545818 185004 546054
rect 184404 545734 185004 545818
rect 184404 545498 184586 545734
rect 184822 545498 185004 545734
rect 184404 510054 185004 545498
rect 184404 509818 184586 510054
rect 184822 509818 185004 510054
rect 184404 509734 185004 509818
rect 184404 509498 184586 509734
rect 184822 509498 185004 509734
rect 184404 474054 185004 509498
rect 184404 473818 184586 474054
rect 184822 473818 185004 474054
rect 184404 473734 185004 473818
rect 184404 473498 184586 473734
rect 184822 473498 185004 473734
rect 184404 438054 185004 473498
rect 184404 437818 184586 438054
rect 184822 437818 185004 438054
rect 184404 437734 185004 437818
rect 184404 437498 184586 437734
rect 184822 437498 185004 437734
rect 184404 402054 185004 437498
rect 184404 401818 184586 402054
rect 184822 401818 185004 402054
rect 184404 401734 185004 401818
rect 184404 401498 184586 401734
rect 184822 401498 185004 401734
rect 184404 366054 185004 401498
rect 184404 365818 184586 366054
rect 184822 365818 185004 366054
rect 184404 365734 185004 365818
rect 184404 365498 184586 365734
rect 184822 365498 185004 365734
rect 184404 330054 185004 365498
rect 184404 329818 184586 330054
rect 184822 329818 185004 330054
rect 184404 329734 185004 329818
rect 184404 329498 184586 329734
rect 184822 329498 185004 329734
rect 184404 294054 185004 329498
rect 184404 293818 184586 294054
rect 184822 293818 185004 294054
rect 184404 293734 185004 293818
rect 184404 293498 184586 293734
rect 184822 293498 185004 293734
rect 184404 258054 185004 293498
rect 184404 257818 184586 258054
rect 184822 257818 185004 258054
rect 184404 257734 185004 257818
rect 184404 257498 184586 257734
rect 184822 257498 185004 257734
rect 184404 222054 185004 257498
rect 184404 221818 184586 222054
rect 184822 221818 185004 222054
rect 184404 221734 185004 221818
rect 184404 221498 184586 221734
rect 184822 221498 185004 221734
rect 184404 186054 185004 221498
rect 184404 185818 184586 186054
rect 184822 185818 185004 186054
rect 184404 185734 185004 185818
rect 184404 185498 184586 185734
rect 184822 185498 185004 185734
rect 184404 150054 185004 185498
rect 184404 149818 184586 150054
rect 184822 149818 185004 150054
rect 184404 149734 185004 149818
rect 184404 149498 184586 149734
rect 184822 149498 185004 149734
rect 184404 114054 185004 149498
rect 184404 113818 184586 114054
rect 184822 113818 185004 114054
rect 184404 113734 185004 113818
rect 184404 113498 184586 113734
rect 184822 113498 185004 113734
rect 184404 78054 185004 113498
rect 184404 77818 184586 78054
rect 184822 77818 185004 78054
rect 184404 77734 185004 77818
rect 184404 77498 184586 77734
rect 184822 77498 185004 77734
rect 184404 42054 185004 77498
rect 184404 41818 184586 42054
rect 184822 41818 185004 42054
rect 184404 41734 185004 41818
rect 184404 41498 184586 41734
rect 184822 41498 185004 41734
rect 184404 6054 185004 41498
rect 184404 5818 184586 6054
rect 184822 5818 185004 6054
rect 184404 5734 185004 5818
rect 184404 5498 184586 5734
rect 184822 5498 185004 5734
rect 184404 -2186 185004 5498
rect 184404 -2422 184586 -2186
rect 184822 -2422 185004 -2186
rect 184404 -2506 185004 -2422
rect 184404 -2742 184586 -2506
rect 184822 -2742 185004 -2506
rect 184404 -3684 185004 -2742
rect 188004 693654 188604 707962
rect 188004 693418 188186 693654
rect 188422 693418 188604 693654
rect 188004 693334 188604 693418
rect 188004 693098 188186 693334
rect 188422 693098 188604 693334
rect 188004 657654 188604 693098
rect 188004 657418 188186 657654
rect 188422 657418 188604 657654
rect 188004 657334 188604 657418
rect 188004 657098 188186 657334
rect 188422 657098 188604 657334
rect 188004 621654 188604 657098
rect 188004 621418 188186 621654
rect 188422 621418 188604 621654
rect 188004 621334 188604 621418
rect 188004 621098 188186 621334
rect 188422 621098 188604 621334
rect 188004 585654 188604 621098
rect 188004 585418 188186 585654
rect 188422 585418 188604 585654
rect 188004 585334 188604 585418
rect 188004 585098 188186 585334
rect 188422 585098 188604 585334
rect 188004 549654 188604 585098
rect 188004 549418 188186 549654
rect 188422 549418 188604 549654
rect 188004 549334 188604 549418
rect 188004 549098 188186 549334
rect 188422 549098 188604 549334
rect 188004 513654 188604 549098
rect 188004 513418 188186 513654
rect 188422 513418 188604 513654
rect 188004 513334 188604 513418
rect 188004 513098 188186 513334
rect 188422 513098 188604 513334
rect 188004 477654 188604 513098
rect 188004 477418 188186 477654
rect 188422 477418 188604 477654
rect 188004 477334 188604 477418
rect 188004 477098 188186 477334
rect 188422 477098 188604 477334
rect 188004 441654 188604 477098
rect 188004 441418 188186 441654
rect 188422 441418 188604 441654
rect 188004 441334 188604 441418
rect 188004 441098 188186 441334
rect 188422 441098 188604 441334
rect 188004 405654 188604 441098
rect 188004 405418 188186 405654
rect 188422 405418 188604 405654
rect 188004 405334 188604 405418
rect 188004 405098 188186 405334
rect 188422 405098 188604 405334
rect 188004 369654 188604 405098
rect 188004 369418 188186 369654
rect 188422 369418 188604 369654
rect 188004 369334 188604 369418
rect 188004 369098 188186 369334
rect 188422 369098 188604 369334
rect 188004 333654 188604 369098
rect 188004 333418 188186 333654
rect 188422 333418 188604 333654
rect 188004 333334 188604 333418
rect 188004 333098 188186 333334
rect 188422 333098 188604 333334
rect 188004 297654 188604 333098
rect 188004 297418 188186 297654
rect 188422 297418 188604 297654
rect 188004 297334 188604 297418
rect 188004 297098 188186 297334
rect 188422 297098 188604 297334
rect 188004 261654 188604 297098
rect 188004 261418 188186 261654
rect 188422 261418 188604 261654
rect 188004 261334 188604 261418
rect 188004 261098 188186 261334
rect 188422 261098 188604 261334
rect 188004 225654 188604 261098
rect 188004 225418 188186 225654
rect 188422 225418 188604 225654
rect 188004 225334 188604 225418
rect 188004 225098 188186 225334
rect 188422 225098 188604 225334
rect 188004 189654 188604 225098
rect 188004 189418 188186 189654
rect 188422 189418 188604 189654
rect 188004 189334 188604 189418
rect 188004 189098 188186 189334
rect 188422 189098 188604 189334
rect 188004 153654 188604 189098
rect 188004 153418 188186 153654
rect 188422 153418 188604 153654
rect 188004 153334 188604 153418
rect 188004 153098 188186 153334
rect 188422 153098 188604 153334
rect 188004 117654 188604 153098
rect 188004 117418 188186 117654
rect 188422 117418 188604 117654
rect 188004 117334 188604 117418
rect 188004 117098 188186 117334
rect 188422 117098 188604 117334
rect 188004 81654 188604 117098
rect 188004 81418 188186 81654
rect 188422 81418 188604 81654
rect 188004 81334 188604 81418
rect 188004 81098 188186 81334
rect 188422 81098 188604 81334
rect 188004 45654 188604 81098
rect 188004 45418 188186 45654
rect 188422 45418 188604 45654
rect 188004 45334 188604 45418
rect 188004 45098 188186 45334
rect 188422 45098 188604 45334
rect 188004 9654 188604 45098
rect 188004 9418 188186 9654
rect 188422 9418 188604 9654
rect 188004 9334 188604 9418
rect 188004 9098 188186 9334
rect 188422 9098 188604 9334
rect 188004 -4026 188604 9098
rect 188004 -4262 188186 -4026
rect 188422 -4262 188604 -4026
rect 188004 -4346 188604 -4262
rect 188004 -4582 188186 -4346
rect 188422 -4582 188604 -4346
rect 188004 -5524 188604 -4582
rect 191604 697254 192204 709802
rect 209604 711278 210204 711300
rect 209604 711042 209786 711278
rect 210022 711042 210204 711278
rect 209604 710958 210204 711042
rect 209604 710722 209786 710958
rect 210022 710722 210204 710958
rect 206004 709438 206604 709460
rect 206004 709202 206186 709438
rect 206422 709202 206604 709438
rect 206004 709118 206604 709202
rect 206004 708882 206186 709118
rect 206422 708882 206604 709118
rect 202404 707598 203004 707620
rect 202404 707362 202586 707598
rect 202822 707362 203004 707598
rect 202404 707278 203004 707362
rect 202404 707042 202586 707278
rect 202822 707042 203004 707278
rect 191604 697018 191786 697254
rect 192022 697018 192204 697254
rect 191604 696934 192204 697018
rect 191604 696698 191786 696934
rect 192022 696698 192204 696934
rect 191604 661254 192204 696698
rect 191604 661018 191786 661254
rect 192022 661018 192204 661254
rect 191604 660934 192204 661018
rect 191604 660698 191786 660934
rect 192022 660698 192204 660934
rect 191604 625254 192204 660698
rect 191604 625018 191786 625254
rect 192022 625018 192204 625254
rect 191604 624934 192204 625018
rect 191604 624698 191786 624934
rect 192022 624698 192204 624934
rect 191604 589254 192204 624698
rect 191604 589018 191786 589254
rect 192022 589018 192204 589254
rect 191604 588934 192204 589018
rect 191604 588698 191786 588934
rect 192022 588698 192204 588934
rect 191604 553254 192204 588698
rect 198804 705758 199404 705780
rect 198804 705522 198986 705758
rect 199222 705522 199404 705758
rect 198804 705438 199404 705522
rect 198804 705202 198986 705438
rect 199222 705202 199404 705438
rect 198804 668454 199404 705202
rect 198804 668218 198986 668454
rect 199222 668218 199404 668454
rect 198804 668134 199404 668218
rect 198804 667898 198986 668134
rect 199222 667898 199404 668134
rect 198804 632454 199404 667898
rect 198804 632218 198986 632454
rect 199222 632218 199404 632454
rect 198804 632134 199404 632218
rect 198804 631898 198986 632134
rect 199222 631898 199404 632134
rect 198804 596454 199404 631898
rect 198804 596218 198986 596454
rect 199222 596218 199404 596454
rect 198804 596134 199404 596218
rect 198804 595898 198986 596134
rect 199222 595898 199404 596134
rect 193075 562732 193141 562733
rect 193075 562668 193076 562732
rect 193140 562668 193141 562732
rect 193075 562667 193141 562668
rect 193078 561458 193138 562667
rect 196758 561373 196818 562582
rect 196755 561372 196821 561373
rect 196755 561308 196756 561372
rect 196820 561308 196821 561372
rect 196755 561307 196821 561308
rect 191604 553018 191786 553254
rect 192022 553018 192204 553254
rect 191604 552934 192204 553018
rect 191604 552698 191786 552934
rect 192022 552698 192204 552934
rect 191604 517254 192204 552698
rect 191604 517018 191786 517254
rect 192022 517018 192204 517254
rect 191604 516934 192204 517018
rect 191604 516698 191786 516934
rect 192022 516698 192204 516934
rect 191604 481254 192204 516698
rect 191604 481018 191786 481254
rect 192022 481018 192204 481254
rect 191604 480934 192204 481018
rect 191604 480698 191786 480934
rect 192022 480698 192204 480934
rect 191604 445254 192204 480698
rect 191604 445018 191786 445254
rect 192022 445018 192204 445254
rect 191604 444934 192204 445018
rect 191604 444698 191786 444934
rect 192022 444698 192204 444934
rect 191604 409254 192204 444698
rect 191604 409018 191786 409254
rect 192022 409018 192204 409254
rect 191604 408934 192204 409018
rect 191604 408698 191786 408934
rect 192022 408698 192204 408934
rect 191604 373254 192204 408698
rect 191604 373018 191786 373254
rect 192022 373018 192204 373254
rect 191604 372934 192204 373018
rect 191604 372698 191786 372934
rect 192022 372698 192204 372934
rect 191604 337254 192204 372698
rect 191604 337018 191786 337254
rect 192022 337018 192204 337254
rect 191604 336934 192204 337018
rect 191604 336698 191786 336934
rect 192022 336698 192204 336934
rect 191604 301254 192204 336698
rect 191604 301018 191786 301254
rect 192022 301018 192204 301254
rect 191604 300934 192204 301018
rect 191604 300698 191786 300934
rect 192022 300698 192204 300934
rect 191604 265254 192204 300698
rect 191604 265018 191786 265254
rect 192022 265018 192204 265254
rect 191604 264934 192204 265018
rect 191604 264698 191786 264934
rect 192022 264698 192204 264934
rect 191604 229254 192204 264698
rect 191604 229018 191786 229254
rect 192022 229018 192204 229254
rect 191604 228934 192204 229018
rect 191604 228698 191786 228934
rect 192022 228698 192204 228934
rect 191604 193254 192204 228698
rect 191604 193018 191786 193254
rect 192022 193018 192204 193254
rect 191604 192934 192204 193018
rect 191604 192698 191786 192934
rect 192022 192698 192204 192934
rect 191604 157254 192204 192698
rect 191604 157018 191786 157254
rect 192022 157018 192204 157254
rect 191604 156934 192204 157018
rect 191604 156698 191786 156934
rect 192022 156698 192204 156934
rect 191604 121254 192204 156698
rect 191604 121018 191786 121254
rect 192022 121018 192204 121254
rect 191604 120934 192204 121018
rect 191604 120698 191786 120934
rect 192022 120698 192204 120934
rect 191604 85254 192204 120698
rect 191604 85018 191786 85254
rect 192022 85018 192204 85254
rect 191604 84934 192204 85018
rect 191604 84698 191786 84934
rect 192022 84698 192204 84934
rect 191604 49254 192204 84698
rect 191604 49018 191786 49254
rect 192022 49018 192204 49254
rect 191604 48934 192204 49018
rect 191604 48698 191786 48934
rect 192022 48698 192204 48934
rect 191604 13254 192204 48698
rect 191604 13018 191786 13254
rect 192022 13018 192204 13254
rect 191604 12934 192204 13018
rect 191604 12698 191786 12934
rect 192022 12698 192204 12934
rect 173604 -7022 173786 -6786
rect 174022 -7022 174204 -6786
rect 173604 -7106 174204 -7022
rect 173604 -7342 173786 -7106
rect 174022 -7342 174204 -7106
rect 173604 -7364 174204 -7342
rect 191604 -5866 192204 12698
rect 198804 560454 199404 595898
rect 198804 560218 198986 560454
rect 199222 560218 199404 560454
rect 198804 560134 199404 560218
rect 198804 559898 198986 560134
rect 199222 559898 199404 560134
rect 198804 524454 199404 559898
rect 198804 524218 198986 524454
rect 199222 524218 199404 524454
rect 198804 524134 199404 524218
rect 198804 523898 198986 524134
rect 199222 523898 199404 524134
rect 198804 488454 199404 523898
rect 198804 488218 198986 488454
rect 199222 488218 199404 488454
rect 198804 488134 199404 488218
rect 198804 487898 198986 488134
rect 199222 487898 199404 488134
rect 198804 452454 199404 487898
rect 198804 452218 198986 452454
rect 199222 452218 199404 452454
rect 198804 452134 199404 452218
rect 198804 451898 198986 452134
rect 199222 451898 199404 452134
rect 198804 416454 199404 451898
rect 198804 416218 198986 416454
rect 199222 416218 199404 416454
rect 198804 416134 199404 416218
rect 198804 415898 198986 416134
rect 199222 415898 199404 416134
rect 198804 380454 199404 415898
rect 198804 380218 198986 380454
rect 199222 380218 199404 380454
rect 198804 380134 199404 380218
rect 198804 379898 198986 380134
rect 199222 379898 199404 380134
rect 198804 344454 199404 379898
rect 198804 344218 198986 344454
rect 199222 344218 199404 344454
rect 198804 344134 199404 344218
rect 198804 343898 198986 344134
rect 199222 343898 199404 344134
rect 198804 308454 199404 343898
rect 198804 308218 198986 308454
rect 199222 308218 199404 308454
rect 198804 308134 199404 308218
rect 198804 307898 198986 308134
rect 199222 307898 199404 308134
rect 198804 272454 199404 307898
rect 198804 272218 198986 272454
rect 199222 272218 199404 272454
rect 198804 272134 199404 272218
rect 198804 271898 198986 272134
rect 199222 271898 199404 272134
rect 198804 236454 199404 271898
rect 198804 236218 198986 236454
rect 199222 236218 199404 236454
rect 198804 236134 199404 236218
rect 198804 235898 198986 236134
rect 199222 235898 199404 236134
rect 198804 200454 199404 235898
rect 198804 200218 198986 200454
rect 199222 200218 199404 200454
rect 198804 200134 199404 200218
rect 198804 199898 198986 200134
rect 199222 199898 199404 200134
rect 198804 164454 199404 199898
rect 198804 164218 198986 164454
rect 199222 164218 199404 164454
rect 198804 164134 199404 164218
rect 198804 163898 198986 164134
rect 199222 163898 199404 164134
rect 198804 128454 199404 163898
rect 198804 128218 198986 128454
rect 199222 128218 199404 128454
rect 198804 128134 199404 128218
rect 198804 127898 198986 128134
rect 199222 127898 199404 128134
rect 198804 92454 199404 127898
rect 198804 92218 198986 92454
rect 199222 92218 199404 92454
rect 198804 92134 199404 92218
rect 198804 91898 198986 92134
rect 199222 91898 199404 92134
rect 198804 56454 199404 91898
rect 198804 56218 198986 56454
rect 199222 56218 199404 56454
rect 198804 56134 199404 56218
rect 198804 55898 198986 56134
rect 199222 55898 199404 56134
rect 198804 20454 199404 55898
rect 198804 20218 198986 20454
rect 199222 20218 199404 20454
rect 198804 20134 199404 20218
rect 198804 19898 198986 20134
rect 199222 19898 199404 20134
rect 198804 -1266 199404 19898
rect 198804 -1502 198986 -1266
rect 199222 -1502 199404 -1266
rect 198804 -1586 199404 -1502
rect 198804 -1822 198986 -1586
rect 199222 -1822 199404 -1586
rect 198804 -1844 199404 -1822
rect 202404 672054 203004 707042
rect 202404 671818 202586 672054
rect 202822 671818 203004 672054
rect 202404 671734 203004 671818
rect 202404 671498 202586 671734
rect 202822 671498 203004 671734
rect 202404 636054 203004 671498
rect 202404 635818 202586 636054
rect 202822 635818 203004 636054
rect 202404 635734 203004 635818
rect 202404 635498 202586 635734
rect 202822 635498 203004 635734
rect 202404 600054 203004 635498
rect 202404 599818 202586 600054
rect 202822 599818 203004 600054
rect 202404 599734 203004 599818
rect 202404 599498 202586 599734
rect 202822 599498 203004 599734
rect 202404 564054 203004 599498
rect 202404 563818 202586 564054
rect 202822 563818 203004 564054
rect 202404 563734 203004 563818
rect 202404 563498 202586 563734
rect 202822 563498 203004 563734
rect 202404 528054 203004 563498
rect 206004 675654 206604 708882
rect 206004 675418 206186 675654
rect 206422 675418 206604 675654
rect 206004 675334 206604 675418
rect 206004 675098 206186 675334
rect 206422 675098 206604 675334
rect 206004 639654 206604 675098
rect 206004 639418 206186 639654
rect 206422 639418 206604 639654
rect 206004 639334 206604 639418
rect 206004 639098 206186 639334
rect 206422 639098 206604 639334
rect 206004 603654 206604 639098
rect 206004 603418 206186 603654
rect 206422 603418 206604 603654
rect 206004 603334 206604 603418
rect 206004 603098 206186 603334
rect 206422 603098 206604 603334
rect 206004 567654 206604 603098
rect 206004 567418 206186 567654
rect 206422 567418 206604 567654
rect 206004 567334 206604 567418
rect 206004 567098 206186 567334
rect 206422 567098 206604 567334
rect 202404 527818 202586 528054
rect 202822 527818 203004 528054
rect 202404 527734 203004 527818
rect 202404 527498 202586 527734
rect 202822 527498 203004 527734
rect 202404 492054 203004 527498
rect 202404 491818 202586 492054
rect 202822 491818 203004 492054
rect 202404 491734 203004 491818
rect 202404 491498 202586 491734
rect 202822 491498 203004 491734
rect 202404 456054 203004 491498
rect 202404 455818 202586 456054
rect 202822 455818 203004 456054
rect 202404 455734 203004 455818
rect 202404 455498 202586 455734
rect 202822 455498 203004 455734
rect 202404 420054 203004 455498
rect 202404 419818 202586 420054
rect 202822 419818 203004 420054
rect 202404 419734 203004 419818
rect 202404 419498 202586 419734
rect 202822 419498 203004 419734
rect 202404 384054 203004 419498
rect 202404 383818 202586 384054
rect 202822 383818 203004 384054
rect 202404 383734 203004 383818
rect 202404 383498 202586 383734
rect 202822 383498 203004 383734
rect 202404 348054 203004 383498
rect 202404 347818 202586 348054
rect 202822 347818 203004 348054
rect 202404 347734 203004 347818
rect 202404 347498 202586 347734
rect 202822 347498 203004 347734
rect 202404 312054 203004 347498
rect 202404 311818 202586 312054
rect 202822 311818 203004 312054
rect 202404 311734 203004 311818
rect 202404 311498 202586 311734
rect 202822 311498 203004 311734
rect 202404 276054 203004 311498
rect 202404 275818 202586 276054
rect 202822 275818 203004 276054
rect 202404 275734 203004 275818
rect 202404 275498 202586 275734
rect 202822 275498 203004 275734
rect 202404 240054 203004 275498
rect 202404 239818 202586 240054
rect 202822 239818 203004 240054
rect 202404 239734 203004 239818
rect 202404 239498 202586 239734
rect 202822 239498 203004 239734
rect 202404 204054 203004 239498
rect 202404 203818 202586 204054
rect 202822 203818 203004 204054
rect 202404 203734 203004 203818
rect 202404 203498 202586 203734
rect 202822 203498 203004 203734
rect 202404 168054 203004 203498
rect 202404 167818 202586 168054
rect 202822 167818 203004 168054
rect 202404 167734 203004 167818
rect 202404 167498 202586 167734
rect 202822 167498 203004 167734
rect 202404 132054 203004 167498
rect 202404 131818 202586 132054
rect 202822 131818 203004 132054
rect 202404 131734 203004 131818
rect 202404 131498 202586 131734
rect 202822 131498 203004 131734
rect 202404 96054 203004 131498
rect 202404 95818 202586 96054
rect 202822 95818 203004 96054
rect 202404 95734 203004 95818
rect 202404 95498 202586 95734
rect 202822 95498 203004 95734
rect 202404 60054 203004 95498
rect 202404 59818 202586 60054
rect 202822 59818 203004 60054
rect 202404 59734 203004 59818
rect 202404 59498 202586 59734
rect 202822 59498 203004 59734
rect 202404 24054 203004 59498
rect 202404 23818 202586 24054
rect 202822 23818 203004 24054
rect 202404 23734 203004 23818
rect 202404 23498 202586 23734
rect 202822 23498 203004 23734
rect 202404 -3106 203004 23498
rect 202404 -3342 202586 -3106
rect 202822 -3342 203004 -3106
rect 202404 -3426 203004 -3342
rect 202404 -3662 202586 -3426
rect 202822 -3662 203004 -3426
rect 202404 -3684 203004 -3662
rect 206004 531654 206604 567098
rect 209604 679254 210204 710722
rect 227604 710358 228204 711300
rect 227604 710122 227786 710358
rect 228022 710122 228204 710358
rect 227604 710038 228204 710122
rect 227604 709802 227786 710038
rect 228022 709802 228204 710038
rect 224004 708518 224604 709460
rect 224004 708282 224186 708518
rect 224422 708282 224604 708518
rect 224004 708198 224604 708282
rect 224004 707962 224186 708198
rect 224422 707962 224604 708198
rect 220404 706678 221004 707620
rect 220404 706442 220586 706678
rect 220822 706442 221004 706678
rect 220404 706358 221004 706442
rect 220404 706122 220586 706358
rect 220822 706122 221004 706358
rect 209604 679018 209786 679254
rect 210022 679018 210204 679254
rect 209604 678934 210204 679018
rect 209604 678698 209786 678934
rect 210022 678698 210204 678934
rect 209604 643254 210204 678698
rect 209604 643018 209786 643254
rect 210022 643018 210204 643254
rect 209604 642934 210204 643018
rect 209604 642698 209786 642934
rect 210022 642698 210204 642934
rect 209604 607254 210204 642698
rect 209604 607018 209786 607254
rect 210022 607018 210204 607254
rect 209604 606934 210204 607018
rect 209604 606698 209786 606934
rect 210022 606698 210204 606934
rect 209604 571254 210204 606698
rect 209604 571018 209786 571254
rect 210022 571018 210204 571254
rect 209604 570934 210204 571018
rect 209604 570698 209786 570934
rect 210022 570698 210204 570934
rect 207611 562732 207677 562733
rect 207611 562668 207612 562732
rect 207676 562668 207677 562732
rect 207611 562667 207677 562668
rect 207614 561458 207674 562667
rect 206004 531418 206186 531654
rect 206422 531418 206604 531654
rect 206004 531334 206604 531418
rect 206004 531098 206186 531334
rect 206422 531098 206604 531334
rect 206004 495654 206604 531098
rect 206004 495418 206186 495654
rect 206422 495418 206604 495654
rect 206004 495334 206604 495418
rect 206004 495098 206186 495334
rect 206422 495098 206604 495334
rect 206004 459654 206604 495098
rect 206004 459418 206186 459654
rect 206422 459418 206604 459654
rect 206004 459334 206604 459418
rect 206004 459098 206186 459334
rect 206422 459098 206604 459334
rect 206004 423654 206604 459098
rect 206004 423418 206186 423654
rect 206422 423418 206604 423654
rect 206004 423334 206604 423418
rect 206004 423098 206186 423334
rect 206422 423098 206604 423334
rect 206004 387654 206604 423098
rect 206004 387418 206186 387654
rect 206422 387418 206604 387654
rect 206004 387334 206604 387418
rect 206004 387098 206186 387334
rect 206422 387098 206604 387334
rect 206004 351654 206604 387098
rect 206004 351418 206186 351654
rect 206422 351418 206604 351654
rect 206004 351334 206604 351418
rect 206004 351098 206186 351334
rect 206422 351098 206604 351334
rect 206004 315654 206604 351098
rect 206004 315418 206186 315654
rect 206422 315418 206604 315654
rect 206004 315334 206604 315418
rect 206004 315098 206186 315334
rect 206422 315098 206604 315334
rect 206004 279654 206604 315098
rect 206004 279418 206186 279654
rect 206422 279418 206604 279654
rect 206004 279334 206604 279418
rect 206004 279098 206186 279334
rect 206422 279098 206604 279334
rect 206004 243654 206604 279098
rect 206004 243418 206186 243654
rect 206422 243418 206604 243654
rect 206004 243334 206604 243418
rect 206004 243098 206186 243334
rect 206422 243098 206604 243334
rect 206004 207654 206604 243098
rect 206004 207418 206186 207654
rect 206422 207418 206604 207654
rect 206004 207334 206604 207418
rect 206004 207098 206186 207334
rect 206422 207098 206604 207334
rect 206004 171654 206604 207098
rect 206004 171418 206186 171654
rect 206422 171418 206604 171654
rect 206004 171334 206604 171418
rect 206004 171098 206186 171334
rect 206422 171098 206604 171334
rect 206004 135654 206604 171098
rect 206004 135418 206186 135654
rect 206422 135418 206604 135654
rect 206004 135334 206604 135418
rect 206004 135098 206186 135334
rect 206422 135098 206604 135334
rect 206004 99654 206604 135098
rect 206004 99418 206186 99654
rect 206422 99418 206604 99654
rect 206004 99334 206604 99418
rect 206004 99098 206186 99334
rect 206422 99098 206604 99334
rect 206004 63654 206604 99098
rect 206004 63418 206186 63654
rect 206422 63418 206604 63654
rect 206004 63334 206604 63418
rect 206004 63098 206186 63334
rect 206422 63098 206604 63334
rect 206004 27654 206604 63098
rect 206004 27418 206186 27654
rect 206422 27418 206604 27654
rect 206004 27334 206604 27418
rect 206004 27098 206186 27334
rect 206422 27098 206604 27334
rect 206004 -4946 206604 27098
rect 206004 -5182 206186 -4946
rect 206422 -5182 206604 -4946
rect 206004 -5266 206604 -5182
rect 206004 -5502 206186 -5266
rect 206422 -5502 206604 -5266
rect 206004 -5524 206604 -5502
rect 209604 535254 210204 570698
rect 209604 535018 209786 535254
rect 210022 535018 210204 535254
rect 209604 534934 210204 535018
rect 209604 534698 209786 534934
rect 210022 534698 210204 534934
rect 209604 499254 210204 534698
rect 209604 499018 209786 499254
rect 210022 499018 210204 499254
rect 209604 498934 210204 499018
rect 209604 498698 209786 498934
rect 210022 498698 210204 498934
rect 209604 463254 210204 498698
rect 209604 463018 209786 463254
rect 210022 463018 210204 463254
rect 209604 462934 210204 463018
rect 209604 462698 209786 462934
rect 210022 462698 210204 462934
rect 209604 427254 210204 462698
rect 209604 427018 209786 427254
rect 210022 427018 210204 427254
rect 209604 426934 210204 427018
rect 209604 426698 209786 426934
rect 210022 426698 210204 426934
rect 209604 391254 210204 426698
rect 209604 391018 209786 391254
rect 210022 391018 210204 391254
rect 209604 390934 210204 391018
rect 209604 390698 209786 390934
rect 210022 390698 210204 390934
rect 209604 355254 210204 390698
rect 209604 355018 209786 355254
rect 210022 355018 210204 355254
rect 209604 354934 210204 355018
rect 209604 354698 209786 354934
rect 210022 354698 210204 354934
rect 209604 319254 210204 354698
rect 209604 319018 209786 319254
rect 210022 319018 210204 319254
rect 209604 318934 210204 319018
rect 209604 318698 209786 318934
rect 210022 318698 210204 318934
rect 209604 283254 210204 318698
rect 209604 283018 209786 283254
rect 210022 283018 210204 283254
rect 209604 282934 210204 283018
rect 209604 282698 209786 282934
rect 210022 282698 210204 282934
rect 209604 247254 210204 282698
rect 209604 247018 209786 247254
rect 210022 247018 210204 247254
rect 209604 246934 210204 247018
rect 209604 246698 209786 246934
rect 210022 246698 210204 246934
rect 209604 211254 210204 246698
rect 209604 211018 209786 211254
rect 210022 211018 210204 211254
rect 209604 210934 210204 211018
rect 209604 210698 209786 210934
rect 210022 210698 210204 210934
rect 209604 175254 210204 210698
rect 209604 175018 209786 175254
rect 210022 175018 210204 175254
rect 209604 174934 210204 175018
rect 209604 174698 209786 174934
rect 210022 174698 210204 174934
rect 209604 139254 210204 174698
rect 209604 139018 209786 139254
rect 210022 139018 210204 139254
rect 209604 138934 210204 139018
rect 209604 138698 209786 138934
rect 210022 138698 210204 138934
rect 209604 103254 210204 138698
rect 209604 103018 209786 103254
rect 210022 103018 210204 103254
rect 209604 102934 210204 103018
rect 209604 102698 209786 102934
rect 210022 102698 210204 102934
rect 209604 67254 210204 102698
rect 209604 67018 209786 67254
rect 210022 67018 210204 67254
rect 209604 66934 210204 67018
rect 209604 66698 209786 66934
rect 210022 66698 210204 66934
rect 209604 31254 210204 66698
rect 209604 31018 209786 31254
rect 210022 31018 210204 31254
rect 209604 30934 210204 31018
rect 209604 30698 209786 30934
rect 210022 30698 210204 30934
rect 191604 -6102 191786 -5866
rect 192022 -6102 192204 -5866
rect 191604 -6186 192204 -6102
rect 191604 -6422 191786 -6186
rect 192022 -6422 192204 -6186
rect 191604 -7364 192204 -6422
rect 209604 -6786 210204 30698
rect 216804 704838 217404 705780
rect 216804 704602 216986 704838
rect 217222 704602 217404 704838
rect 216804 704518 217404 704602
rect 216804 704282 216986 704518
rect 217222 704282 217404 704518
rect 216804 686454 217404 704282
rect 216804 686218 216986 686454
rect 217222 686218 217404 686454
rect 216804 686134 217404 686218
rect 216804 685898 216986 686134
rect 217222 685898 217404 686134
rect 216804 650454 217404 685898
rect 216804 650218 216986 650454
rect 217222 650218 217404 650454
rect 216804 650134 217404 650218
rect 216804 649898 216986 650134
rect 217222 649898 217404 650134
rect 216804 614454 217404 649898
rect 216804 614218 216986 614454
rect 217222 614218 217404 614454
rect 216804 614134 217404 614218
rect 216804 613898 216986 614134
rect 217222 613898 217404 614134
rect 216804 578454 217404 613898
rect 216804 578218 216986 578454
rect 217222 578218 217404 578454
rect 216804 578134 217404 578218
rect 216804 577898 216986 578134
rect 217222 577898 217404 578134
rect 216804 542454 217404 577898
rect 216804 542218 216986 542454
rect 217222 542218 217404 542454
rect 216804 542134 217404 542218
rect 216804 541898 216986 542134
rect 217222 541898 217404 542134
rect 216804 506454 217404 541898
rect 216804 506218 216986 506454
rect 217222 506218 217404 506454
rect 216804 506134 217404 506218
rect 216804 505898 216986 506134
rect 217222 505898 217404 506134
rect 216804 470454 217404 505898
rect 216804 470218 216986 470454
rect 217222 470218 217404 470454
rect 216804 470134 217404 470218
rect 216804 469898 216986 470134
rect 217222 469898 217404 470134
rect 216804 434454 217404 469898
rect 216804 434218 216986 434454
rect 217222 434218 217404 434454
rect 216804 434134 217404 434218
rect 216804 433898 216986 434134
rect 217222 433898 217404 434134
rect 216804 398454 217404 433898
rect 216804 398218 216986 398454
rect 217222 398218 217404 398454
rect 216804 398134 217404 398218
rect 216804 397898 216986 398134
rect 217222 397898 217404 398134
rect 216804 362454 217404 397898
rect 216804 362218 216986 362454
rect 217222 362218 217404 362454
rect 216804 362134 217404 362218
rect 216804 361898 216986 362134
rect 217222 361898 217404 362134
rect 216804 326454 217404 361898
rect 216804 326218 216986 326454
rect 217222 326218 217404 326454
rect 216804 326134 217404 326218
rect 216804 325898 216986 326134
rect 217222 325898 217404 326134
rect 216804 290454 217404 325898
rect 216804 290218 216986 290454
rect 217222 290218 217404 290454
rect 216804 290134 217404 290218
rect 216804 289898 216986 290134
rect 217222 289898 217404 290134
rect 216804 254454 217404 289898
rect 216804 254218 216986 254454
rect 217222 254218 217404 254454
rect 216804 254134 217404 254218
rect 216804 253898 216986 254134
rect 217222 253898 217404 254134
rect 216804 218454 217404 253898
rect 216804 218218 216986 218454
rect 217222 218218 217404 218454
rect 216804 218134 217404 218218
rect 216804 217898 216986 218134
rect 217222 217898 217404 218134
rect 216804 182454 217404 217898
rect 216804 182218 216986 182454
rect 217222 182218 217404 182454
rect 216804 182134 217404 182218
rect 216804 181898 216986 182134
rect 217222 181898 217404 182134
rect 216804 146454 217404 181898
rect 216804 146218 216986 146454
rect 217222 146218 217404 146454
rect 216804 146134 217404 146218
rect 216804 145898 216986 146134
rect 217222 145898 217404 146134
rect 216804 110454 217404 145898
rect 216804 110218 216986 110454
rect 217222 110218 217404 110454
rect 216804 110134 217404 110218
rect 216804 109898 216986 110134
rect 217222 109898 217404 110134
rect 216804 74454 217404 109898
rect 216804 74218 216986 74454
rect 217222 74218 217404 74454
rect 216804 74134 217404 74218
rect 216804 73898 216986 74134
rect 217222 73898 217404 74134
rect 216804 38454 217404 73898
rect 216804 38218 216986 38454
rect 217222 38218 217404 38454
rect 216804 38134 217404 38218
rect 216804 37898 216986 38134
rect 217222 37898 217404 38134
rect 216804 2454 217404 37898
rect 216804 2218 216986 2454
rect 217222 2218 217404 2454
rect 216804 2134 217404 2218
rect 216804 1898 216986 2134
rect 217222 1898 217404 2134
rect 216804 -346 217404 1898
rect 216804 -582 216986 -346
rect 217222 -582 217404 -346
rect 216804 -666 217404 -582
rect 216804 -902 216986 -666
rect 217222 -902 217404 -666
rect 216804 -1844 217404 -902
rect 220404 690054 221004 706122
rect 220404 689818 220586 690054
rect 220822 689818 221004 690054
rect 220404 689734 221004 689818
rect 220404 689498 220586 689734
rect 220822 689498 221004 689734
rect 220404 654054 221004 689498
rect 220404 653818 220586 654054
rect 220822 653818 221004 654054
rect 220404 653734 221004 653818
rect 220404 653498 220586 653734
rect 220822 653498 221004 653734
rect 220404 618054 221004 653498
rect 220404 617818 220586 618054
rect 220822 617818 221004 618054
rect 220404 617734 221004 617818
rect 220404 617498 220586 617734
rect 220822 617498 221004 617734
rect 220404 582054 221004 617498
rect 220404 581818 220586 582054
rect 220822 581818 221004 582054
rect 220404 581734 221004 581818
rect 220404 581498 220586 581734
rect 220822 581498 221004 581734
rect 220404 546054 221004 581498
rect 224004 693654 224604 707962
rect 224004 693418 224186 693654
rect 224422 693418 224604 693654
rect 224004 693334 224604 693418
rect 224004 693098 224186 693334
rect 224422 693098 224604 693334
rect 224004 657654 224604 693098
rect 224004 657418 224186 657654
rect 224422 657418 224604 657654
rect 224004 657334 224604 657418
rect 224004 657098 224186 657334
rect 224422 657098 224604 657334
rect 224004 621654 224604 657098
rect 224004 621418 224186 621654
rect 224422 621418 224604 621654
rect 224004 621334 224604 621418
rect 224004 621098 224186 621334
rect 224422 621098 224604 621334
rect 224004 585654 224604 621098
rect 224004 585418 224186 585654
rect 224422 585418 224604 585654
rect 224004 585334 224604 585418
rect 224004 585098 224186 585334
rect 224422 585098 224604 585334
rect 222147 559468 222213 559469
rect 222147 559404 222148 559468
rect 222212 559404 222213 559468
rect 222147 559403 222213 559404
rect 222150 559197 222210 559403
rect 222147 559196 222213 559197
rect 222147 559132 222148 559196
rect 222212 559132 222213 559196
rect 222147 559131 222213 559132
rect 220404 545818 220586 546054
rect 220822 545818 221004 546054
rect 220404 545734 221004 545818
rect 220404 545498 220586 545734
rect 220822 545498 221004 545734
rect 220404 510054 221004 545498
rect 220404 509818 220586 510054
rect 220822 509818 221004 510054
rect 220404 509734 221004 509818
rect 220404 509498 220586 509734
rect 220822 509498 221004 509734
rect 220404 474054 221004 509498
rect 220404 473818 220586 474054
rect 220822 473818 221004 474054
rect 220404 473734 221004 473818
rect 220404 473498 220586 473734
rect 220822 473498 221004 473734
rect 220404 438054 221004 473498
rect 220404 437818 220586 438054
rect 220822 437818 221004 438054
rect 220404 437734 221004 437818
rect 220404 437498 220586 437734
rect 220822 437498 221004 437734
rect 220404 402054 221004 437498
rect 220404 401818 220586 402054
rect 220822 401818 221004 402054
rect 220404 401734 221004 401818
rect 220404 401498 220586 401734
rect 220822 401498 221004 401734
rect 220404 366054 221004 401498
rect 220404 365818 220586 366054
rect 220822 365818 221004 366054
rect 220404 365734 221004 365818
rect 220404 365498 220586 365734
rect 220822 365498 221004 365734
rect 220404 330054 221004 365498
rect 220404 329818 220586 330054
rect 220822 329818 221004 330054
rect 220404 329734 221004 329818
rect 220404 329498 220586 329734
rect 220822 329498 221004 329734
rect 220404 294054 221004 329498
rect 220404 293818 220586 294054
rect 220822 293818 221004 294054
rect 220404 293734 221004 293818
rect 220404 293498 220586 293734
rect 220822 293498 221004 293734
rect 220404 258054 221004 293498
rect 220404 257818 220586 258054
rect 220822 257818 221004 258054
rect 220404 257734 221004 257818
rect 220404 257498 220586 257734
rect 220822 257498 221004 257734
rect 220404 222054 221004 257498
rect 220404 221818 220586 222054
rect 220822 221818 221004 222054
rect 220404 221734 221004 221818
rect 220404 221498 220586 221734
rect 220822 221498 221004 221734
rect 220404 186054 221004 221498
rect 220404 185818 220586 186054
rect 220822 185818 221004 186054
rect 220404 185734 221004 185818
rect 220404 185498 220586 185734
rect 220822 185498 221004 185734
rect 220404 150054 221004 185498
rect 220404 149818 220586 150054
rect 220822 149818 221004 150054
rect 220404 149734 221004 149818
rect 220404 149498 220586 149734
rect 220822 149498 221004 149734
rect 220404 114054 221004 149498
rect 220404 113818 220586 114054
rect 220822 113818 221004 114054
rect 220404 113734 221004 113818
rect 220404 113498 220586 113734
rect 220822 113498 221004 113734
rect 220404 78054 221004 113498
rect 220404 77818 220586 78054
rect 220822 77818 221004 78054
rect 220404 77734 221004 77818
rect 220404 77498 220586 77734
rect 220822 77498 221004 77734
rect 220404 42054 221004 77498
rect 220404 41818 220586 42054
rect 220822 41818 221004 42054
rect 220404 41734 221004 41818
rect 220404 41498 220586 41734
rect 220822 41498 221004 41734
rect 220404 6054 221004 41498
rect 220404 5818 220586 6054
rect 220822 5818 221004 6054
rect 220404 5734 221004 5818
rect 220404 5498 220586 5734
rect 220822 5498 221004 5734
rect 220404 -2186 221004 5498
rect 220404 -2422 220586 -2186
rect 220822 -2422 221004 -2186
rect 220404 -2506 221004 -2422
rect 220404 -2742 220586 -2506
rect 220822 -2742 221004 -2506
rect 220404 -3684 221004 -2742
rect 224004 549654 224604 585098
rect 227604 697254 228204 709802
rect 245604 711278 246204 711300
rect 245604 711042 245786 711278
rect 246022 711042 246204 711278
rect 245604 710958 246204 711042
rect 245604 710722 245786 710958
rect 246022 710722 246204 710958
rect 242004 709438 242604 709460
rect 242004 709202 242186 709438
rect 242422 709202 242604 709438
rect 242004 709118 242604 709202
rect 242004 708882 242186 709118
rect 242422 708882 242604 709118
rect 238404 707598 239004 707620
rect 238404 707362 238586 707598
rect 238822 707362 239004 707598
rect 238404 707278 239004 707362
rect 238404 707042 238586 707278
rect 238822 707042 239004 707278
rect 227604 697018 227786 697254
rect 228022 697018 228204 697254
rect 227604 696934 228204 697018
rect 227604 696698 227786 696934
rect 228022 696698 228204 696934
rect 227604 661254 228204 696698
rect 227604 661018 227786 661254
rect 228022 661018 228204 661254
rect 227604 660934 228204 661018
rect 227604 660698 227786 660934
rect 228022 660698 228204 660934
rect 227604 625254 228204 660698
rect 227604 625018 227786 625254
rect 228022 625018 228204 625254
rect 227604 624934 228204 625018
rect 227604 624698 227786 624934
rect 228022 624698 228204 624934
rect 227604 589254 228204 624698
rect 227604 589018 227786 589254
rect 228022 589018 228204 589254
rect 227604 588934 228204 589018
rect 227604 588698 227786 588934
rect 228022 588698 228204 588934
rect 225462 561373 225522 561902
rect 225459 561372 225525 561373
rect 225459 561308 225460 561372
rect 225524 561308 225525 561372
rect 225459 561307 225525 561308
rect 224004 549418 224186 549654
rect 224422 549418 224604 549654
rect 224004 549334 224604 549418
rect 224004 549098 224186 549334
rect 224422 549098 224604 549334
rect 224004 513654 224604 549098
rect 224004 513418 224186 513654
rect 224422 513418 224604 513654
rect 224004 513334 224604 513418
rect 224004 513098 224186 513334
rect 224422 513098 224604 513334
rect 224004 477654 224604 513098
rect 224004 477418 224186 477654
rect 224422 477418 224604 477654
rect 224004 477334 224604 477418
rect 224004 477098 224186 477334
rect 224422 477098 224604 477334
rect 224004 441654 224604 477098
rect 224004 441418 224186 441654
rect 224422 441418 224604 441654
rect 224004 441334 224604 441418
rect 224004 441098 224186 441334
rect 224422 441098 224604 441334
rect 224004 405654 224604 441098
rect 224004 405418 224186 405654
rect 224422 405418 224604 405654
rect 224004 405334 224604 405418
rect 224004 405098 224186 405334
rect 224422 405098 224604 405334
rect 224004 369654 224604 405098
rect 224004 369418 224186 369654
rect 224422 369418 224604 369654
rect 224004 369334 224604 369418
rect 224004 369098 224186 369334
rect 224422 369098 224604 369334
rect 224004 333654 224604 369098
rect 224004 333418 224186 333654
rect 224422 333418 224604 333654
rect 224004 333334 224604 333418
rect 224004 333098 224186 333334
rect 224422 333098 224604 333334
rect 224004 297654 224604 333098
rect 224004 297418 224186 297654
rect 224422 297418 224604 297654
rect 224004 297334 224604 297418
rect 224004 297098 224186 297334
rect 224422 297098 224604 297334
rect 224004 261654 224604 297098
rect 224004 261418 224186 261654
rect 224422 261418 224604 261654
rect 224004 261334 224604 261418
rect 224004 261098 224186 261334
rect 224422 261098 224604 261334
rect 224004 225654 224604 261098
rect 224004 225418 224186 225654
rect 224422 225418 224604 225654
rect 224004 225334 224604 225418
rect 224004 225098 224186 225334
rect 224422 225098 224604 225334
rect 224004 189654 224604 225098
rect 224004 189418 224186 189654
rect 224422 189418 224604 189654
rect 224004 189334 224604 189418
rect 224004 189098 224186 189334
rect 224422 189098 224604 189334
rect 224004 153654 224604 189098
rect 224004 153418 224186 153654
rect 224422 153418 224604 153654
rect 224004 153334 224604 153418
rect 224004 153098 224186 153334
rect 224422 153098 224604 153334
rect 224004 117654 224604 153098
rect 224004 117418 224186 117654
rect 224422 117418 224604 117654
rect 224004 117334 224604 117418
rect 224004 117098 224186 117334
rect 224422 117098 224604 117334
rect 224004 81654 224604 117098
rect 224004 81418 224186 81654
rect 224422 81418 224604 81654
rect 224004 81334 224604 81418
rect 224004 81098 224186 81334
rect 224422 81098 224604 81334
rect 224004 45654 224604 81098
rect 224004 45418 224186 45654
rect 224422 45418 224604 45654
rect 224004 45334 224604 45418
rect 224004 45098 224186 45334
rect 224422 45098 224604 45334
rect 224004 9654 224604 45098
rect 224004 9418 224186 9654
rect 224422 9418 224604 9654
rect 224004 9334 224604 9418
rect 224004 9098 224186 9334
rect 224422 9098 224604 9334
rect 224004 -4026 224604 9098
rect 224004 -4262 224186 -4026
rect 224422 -4262 224604 -4026
rect 224004 -4346 224604 -4262
rect 224004 -4582 224186 -4346
rect 224422 -4582 224604 -4346
rect 224004 -5524 224604 -4582
rect 227604 553254 228204 588698
rect 234804 705758 235404 705780
rect 234804 705522 234986 705758
rect 235222 705522 235404 705758
rect 234804 705438 235404 705522
rect 234804 705202 234986 705438
rect 235222 705202 235404 705438
rect 234804 668454 235404 705202
rect 234804 668218 234986 668454
rect 235222 668218 235404 668454
rect 234804 668134 235404 668218
rect 234804 667898 234986 668134
rect 235222 667898 235404 668134
rect 234804 632454 235404 667898
rect 234804 632218 234986 632454
rect 235222 632218 235404 632454
rect 234804 632134 235404 632218
rect 234804 631898 234986 632134
rect 235222 631898 235404 632134
rect 234804 596454 235404 631898
rect 234804 596218 234986 596454
rect 235222 596218 235404 596454
rect 234804 596134 235404 596218
rect 234804 595898 234986 596134
rect 235222 595898 235404 596134
rect 234804 560454 235404 595898
rect 238404 672054 239004 707042
rect 238404 671818 238586 672054
rect 238822 671818 239004 672054
rect 238404 671734 239004 671818
rect 238404 671498 238586 671734
rect 238822 671498 239004 671734
rect 238404 636054 239004 671498
rect 238404 635818 238586 636054
rect 238822 635818 239004 636054
rect 238404 635734 239004 635818
rect 238404 635498 238586 635734
rect 238822 635498 239004 635734
rect 238404 600054 239004 635498
rect 238404 599818 238586 600054
rect 238822 599818 239004 600054
rect 238404 599734 239004 599818
rect 238404 599498 238586 599734
rect 238822 599498 239004 599734
rect 238404 564054 239004 599498
rect 238404 563818 238586 564054
rect 238822 563818 239004 564054
rect 238404 563734 239004 563818
rect 238404 563498 238586 563734
rect 238822 563498 239004 563734
rect 237787 563004 237853 563005
rect 237787 562940 237788 563004
rect 237852 562940 237853 563004
rect 237787 562939 237853 562940
rect 236867 562868 236933 562869
rect 236867 562804 236868 562868
rect 236932 562804 236933 562868
rect 236867 562803 236933 562804
rect 236499 562732 236565 562733
rect 236499 562668 236500 562732
rect 236564 562668 236565 562732
rect 236499 562667 236565 562668
rect 234804 560218 234986 560454
rect 235222 560218 235404 560454
rect 234804 560134 235404 560218
rect 234804 559898 234986 560134
rect 235222 559898 235404 560134
rect 231715 559332 231781 559333
rect 231715 559268 231716 559332
rect 231780 559268 231781 559332
rect 231715 559267 231781 559268
rect 233003 559332 233069 559333
rect 233003 559268 233004 559332
rect 233068 559268 233069 559332
rect 233003 559267 233069 559268
rect 234291 559332 234357 559333
rect 234291 559268 234292 559332
rect 234356 559330 234357 559332
rect 234356 559270 234538 559330
rect 234356 559268 234357 559270
rect 234291 559267 234357 559268
rect 227604 553018 227786 553254
rect 228022 553018 228204 553254
rect 227604 552934 228204 553018
rect 227604 552698 227786 552934
rect 228022 552698 228204 552934
rect 227604 517254 228204 552698
rect 227604 517018 227786 517254
rect 228022 517018 228204 517254
rect 227604 516934 228204 517018
rect 227604 516698 227786 516934
rect 228022 516698 228204 516934
rect 227604 481254 228204 516698
rect 227604 481018 227786 481254
rect 228022 481018 228204 481254
rect 227604 480934 228204 481018
rect 227604 480698 227786 480934
rect 228022 480698 228204 480934
rect 227604 445254 228204 480698
rect 227604 445018 227786 445254
rect 228022 445018 228204 445254
rect 227604 444934 228204 445018
rect 227604 444698 227786 444934
rect 228022 444698 228204 444934
rect 227604 409254 228204 444698
rect 227604 409018 227786 409254
rect 228022 409018 228204 409254
rect 227604 408934 228204 409018
rect 227604 408698 227786 408934
rect 228022 408698 228204 408934
rect 227604 373254 228204 408698
rect 227604 373018 227786 373254
rect 228022 373018 228204 373254
rect 227604 372934 228204 373018
rect 227604 372698 227786 372934
rect 228022 372698 228204 372934
rect 227604 337254 228204 372698
rect 227604 337018 227786 337254
rect 228022 337018 228204 337254
rect 227604 336934 228204 337018
rect 227604 336698 227786 336934
rect 228022 336698 228204 336934
rect 227604 301254 228204 336698
rect 227604 301018 227786 301254
rect 228022 301018 228204 301254
rect 227604 300934 228204 301018
rect 227604 300698 227786 300934
rect 228022 300698 228204 300934
rect 227604 265254 228204 300698
rect 227604 265018 227786 265254
rect 228022 265018 228204 265254
rect 227604 264934 228204 265018
rect 227604 264698 227786 264934
rect 228022 264698 228204 264934
rect 227604 229254 228204 264698
rect 227604 229018 227786 229254
rect 228022 229018 228204 229254
rect 227604 228934 228204 229018
rect 227604 228698 227786 228934
rect 228022 228698 228204 228934
rect 227604 193254 228204 228698
rect 227604 193018 227786 193254
rect 228022 193018 228204 193254
rect 227604 192934 228204 193018
rect 227604 192698 227786 192934
rect 228022 192698 228204 192934
rect 227604 157254 228204 192698
rect 227604 157018 227786 157254
rect 228022 157018 228204 157254
rect 227604 156934 228204 157018
rect 227604 156698 227786 156934
rect 228022 156698 228204 156934
rect 227604 121254 228204 156698
rect 227604 121018 227786 121254
rect 228022 121018 228204 121254
rect 227604 120934 228204 121018
rect 227604 120698 227786 120934
rect 228022 120698 228204 120934
rect 227604 85254 228204 120698
rect 227604 85018 227786 85254
rect 228022 85018 228204 85254
rect 227604 84934 228204 85018
rect 227604 84698 227786 84934
rect 228022 84698 228204 84934
rect 227604 49254 228204 84698
rect 227604 49018 227786 49254
rect 228022 49018 228204 49254
rect 227604 48934 228204 49018
rect 227604 48698 227786 48934
rect 228022 48698 228204 48934
rect 227604 13254 228204 48698
rect 229323 22268 229389 22269
rect 229323 22204 229324 22268
rect 229388 22204 229389 22268
rect 229323 22203 229389 22204
rect 229326 18053 229386 22203
rect 229323 18052 229389 18053
rect 229323 17988 229324 18052
rect 229388 17988 229389 18052
rect 229323 17987 229389 17988
rect 231718 16693 231778 559267
rect 233006 40085 233066 559267
rect 233003 40084 233069 40085
rect 233003 40020 233004 40084
rect 233068 40020 233069 40084
rect 233003 40019 233069 40020
rect 234478 32605 234538 559270
rect 234804 524454 235404 559898
rect 234804 524218 234986 524454
rect 235222 524218 235404 524454
rect 234804 524134 235404 524218
rect 234804 523898 234986 524134
rect 235222 523898 235404 524134
rect 234804 488454 235404 523898
rect 234804 488218 234986 488454
rect 235222 488218 235404 488454
rect 234804 488134 235404 488218
rect 234804 487898 234986 488134
rect 235222 487898 235404 488134
rect 234804 452454 235404 487898
rect 234804 452218 234986 452454
rect 235222 452218 235404 452454
rect 234804 452134 235404 452218
rect 234804 451898 234986 452134
rect 235222 451898 235404 452134
rect 234804 416454 235404 451898
rect 234804 416218 234986 416454
rect 235222 416218 235404 416454
rect 234804 416134 235404 416218
rect 234804 415898 234986 416134
rect 235222 415898 235404 416134
rect 234804 380454 235404 415898
rect 234804 380218 234986 380454
rect 235222 380218 235404 380454
rect 234804 380134 235404 380218
rect 234804 379898 234986 380134
rect 235222 379898 235404 380134
rect 234804 344454 235404 379898
rect 234804 344218 234986 344454
rect 235222 344218 235404 344454
rect 234804 344134 235404 344218
rect 234804 343898 234986 344134
rect 235222 343898 235404 344134
rect 234804 308454 235404 343898
rect 234804 308218 234986 308454
rect 235222 308218 235404 308454
rect 234804 308134 235404 308218
rect 234804 307898 234986 308134
rect 235222 307898 235404 308134
rect 234804 272454 235404 307898
rect 234804 272218 234986 272454
rect 235222 272218 235404 272454
rect 234804 272134 235404 272218
rect 234804 271898 234986 272134
rect 235222 271898 235404 272134
rect 234804 236454 235404 271898
rect 236502 252517 236562 562667
rect 236683 559468 236749 559469
rect 236683 559404 236684 559468
rect 236748 559404 236749 559468
rect 236683 559403 236749 559404
rect 236686 309093 236746 559403
rect 236870 338061 236930 562803
rect 237235 559332 237301 559333
rect 237235 559268 237236 559332
rect 237300 559268 237301 559332
rect 237235 559267 237301 559268
rect 236867 338060 236933 338061
rect 236867 337996 236868 338060
rect 236932 337996 236933 338060
rect 236867 337995 236933 337996
rect 236683 309092 236749 309093
rect 236683 309028 236684 309092
rect 236748 309028 236749 309092
rect 236683 309027 236749 309028
rect 236499 252516 236565 252517
rect 236499 252452 236500 252516
rect 236564 252452 236565 252516
rect 236499 252451 236565 252452
rect 234804 236218 234986 236454
rect 235222 236218 235404 236454
rect 234804 236134 235404 236218
rect 234804 235898 234986 236134
rect 235222 235898 235404 236134
rect 234804 200454 235404 235898
rect 234804 200218 234986 200454
rect 235222 200218 235404 200454
rect 234804 200134 235404 200218
rect 234804 199898 234986 200134
rect 235222 199898 235404 200134
rect 234804 164454 235404 199898
rect 234804 164218 234986 164454
rect 235222 164218 235404 164454
rect 234804 164134 235404 164218
rect 234804 163898 234986 164134
rect 235222 163898 235404 164134
rect 234804 128454 235404 163898
rect 234804 128218 234986 128454
rect 235222 128218 235404 128454
rect 234804 128134 235404 128218
rect 234804 127898 234986 128134
rect 235222 127898 235404 128134
rect 234804 92454 235404 127898
rect 234804 92218 234986 92454
rect 235222 92218 235404 92454
rect 234804 92134 235404 92218
rect 234804 91898 234986 92134
rect 235222 91898 235404 92134
rect 234804 56454 235404 91898
rect 237238 63613 237298 559267
rect 237790 181117 237850 562939
rect 237971 562460 238037 562461
rect 237971 562396 237972 562460
rect 238036 562396 238037 562460
rect 237971 562395 238037 562396
rect 237787 181116 237853 181117
rect 237787 181052 237788 181116
rect 237852 181052 237853 181116
rect 237787 181051 237853 181052
rect 237974 133925 238034 562395
rect 238155 559332 238221 559333
rect 238155 559268 238156 559332
rect 238220 559268 238221 559332
rect 238155 559267 238221 559268
rect 237971 133924 238037 133925
rect 237971 133860 237972 133924
rect 238036 133860 238037 133924
rect 237971 133859 238037 133860
rect 238158 91221 238218 559267
rect 238404 528054 239004 563498
rect 238404 527818 238586 528054
rect 238822 527818 239004 528054
rect 238404 527734 239004 527818
rect 238404 527498 238586 527734
rect 238822 527498 239004 527734
rect 238404 492054 239004 527498
rect 238404 491818 238586 492054
rect 238822 491818 239004 492054
rect 238404 491734 239004 491818
rect 238404 491498 238586 491734
rect 238822 491498 239004 491734
rect 238404 456054 239004 491498
rect 238404 455818 238586 456054
rect 238822 455818 239004 456054
rect 238404 455734 239004 455818
rect 238404 455498 238586 455734
rect 238822 455498 239004 455734
rect 238404 420054 239004 455498
rect 238404 419818 238586 420054
rect 238822 419818 239004 420054
rect 238404 419734 239004 419818
rect 238404 419498 238586 419734
rect 238822 419498 239004 419734
rect 238404 384054 239004 419498
rect 238404 383818 238586 384054
rect 238822 383818 239004 384054
rect 238404 383734 239004 383818
rect 238404 383498 238586 383734
rect 238822 383498 239004 383734
rect 238404 348054 239004 383498
rect 238404 347818 238586 348054
rect 238822 347818 239004 348054
rect 238404 347734 239004 347818
rect 238404 347498 238586 347734
rect 238822 347498 239004 347734
rect 238404 312054 239004 347498
rect 238404 311818 238586 312054
rect 238822 311818 239004 312054
rect 238404 311734 239004 311818
rect 238404 311498 238586 311734
rect 238822 311498 239004 311734
rect 238404 276054 239004 311498
rect 238404 275818 238586 276054
rect 238822 275818 239004 276054
rect 238404 275734 239004 275818
rect 238404 275498 238586 275734
rect 238822 275498 239004 275734
rect 238404 240054 239004 275498
rect 238404 239818 238586 240054
rect 238822 239818 239004 240054
rect 238404 239734 239004 239818
rect 238404 239498 238586 239734
rect 238822 239498 239004 239734
rect 238404 204054 239004 239498
rect 238404 203818 238586 204054
rect 238822 203818 239004 204054
rect 238404 203734 239004 203818
rect 238404 203498 238586 203734
rect 238822 203498 239004 203734
rect 238404 168054 239004 203498
rect 242004 675654 242604 708882
rect 242004 675418 242186 675654
rect 242422 675418 242604 675654
rect 242004 675334 242604 675418
rect 242004 675098 242186 675334
rect 242422 675098 242604 675334
rect 242004 639654 242604 675098
rect 242004 639418 242186 639654
rect 242422 639418 242604 639654
rect 242004 639334 242604 639418
rect 242004 639098 242186 639334
rect 242422 639098 242604 639334
rect 242004 603654 242604 639098
rect 242004 603418 242186 603654
rect 242422 603418 242604 603654
rect 242004 603334 242604 603418
rect 242004 603098 242186 603334
rect 242422 603098 242604 603334
rect 242004 567654 242604 603098
rect 242004 567418 242186 567654
rect 242422 567418 242604 567654
rect 242004 567334 242604 567418
rect 242004 567098 242186 567334
rect 242422 567098 242604 567334
rect 242004 531654 242604 567098
rect 245604 679254 246204 710722
rect 263604 710358 264204 711300
rect 263604 710122 263786 710358
rect 264022 710122 264204 710358
rect 263604 710038 264204 710122
rect 263604 709802 263786 710038
rect 264022 709802 264204 710038
rect 260004 708518 260604 709460
rect 260004 708282 260186 708518
rect 260422 708282 260604 708518
rect 260004 708198 260604 708282
rect 260004 707962 260186 708198
rect 260422 707962 260604 708198
rect 256404 706678 257004 707620
rect 256404 706442 256586 706678
rect 256822 706442 257004 706678
rect 256404 706358 257004 706442
rect 256404 706122 256586 706358
rect 256822 706122 257004 706358
rect 245604 679018 245786 679254
rect 246022 679018 246204 679254
rect 245604 678934 246204 679018
rect 245604 678698 245786 678934
rect 246022 678698 246204 678934
rect 245604 643254 246204 678698
rect 245604 643018 245786 643254
rect 246022 643018 246204 643254
rect 245604 642934 246204 643018
rect 245604 642698 245786 642934
rect 246022 642698 246204 642934
rect 245604 607254 246204 642698
rect 245604 607018 245786 607254
rect 246022 607018 246204 607254
rect 245604 606934 246204 607018
rect 245604 606698 245786 606934
rect 246022 606698 246204 606934
rect 245604 571254 246204 606698
rect 245604 571018 245786 571254
rect 246022 571018 246204 571254
rect 245604 570934 246204 571018
rect 245604 570698 245786 570934
rect 246022 570698 246204 570934
rect 244043 559060 244109 559061
rect 244043 558996 244044 559060
rect 244108 558996 244109 559060
rect 244043 558995 244109 558996
rect 244046 558789 244106 558995
rect 244043 558788 244109 558789
rect 244043 558724 244044 558788
rect 244108 558724 244109 558788
rect 244043 558723 244109 558724
rect 242004 531418 242186 531654
rect 242422 531418 242604 531654
rect 242004 531334 242604 531418
rect 242004 531098 242186 531334
rect 242422 531098 242604 531334
rect 242004 495654 242604 531098
rect 242004 495418 242186 495654
rect 242422 495418 242604 495654
rect 242004 495334 242604 495418
rect 242004 495098 242186 495334
rect 242422 495098 242604 495334
rect 242004 459654 242604 495098
rect 242004 459418 242186 459654
rect 242422 459418 242604 459654
rect 242004 459334 242604 459418
rect 242004 459098 242186 459334
rect 242422 459098 242604 459334
rect 242004 423654 242604 459098
rect 242004 423418 242186 423654
rect 242422 423418 242604 423654
rect 242004 423334 242604 423418
rect 242004 423098 242186 423334
rect 242422 423098 242604 423334
rect 242004 387654 242604 423098
rect 242004 387418 242186 387654
rect 242422 387418 242604 387654
rect 242004 387334 242604 387418
rect 242004 387098 242186 387334
rect 242422 387098 242604 387334
rect 242004 351654 242604 387098
rect 242004 351418 242186 351654
rect 242422 351418 242604 351654
rect 242004 351334 242604 351418
rect 242004 351098 242186 351334
rect 242422 351098 242604 351334
rect 242004 315654 242604 351098
rect 242004 315418 242186 315654
rect 242422 315418 242604 315654
rect 242004 315334 242604 315418
rect 242004 315098 242186 315334
rect 242422 315098 242604 315334
rect 242004 279654 242604 315098
rect 242004 279418 242186 279654
rect 242422 279418 242604 279654
rect 242004 279334 242604 279418
rect 242004 279098 242186 279334
rect 242422 279098 242604 279334
rect 242004 243654 242604 279098
rect 242004 243418 242186 243654
rect 242422 243418 242604 243654
rect 242004 243334 242604 243418
rect 242004 243098 242186 243334
rect 242422 243098 242604 243334
rect 242004 207654 242604 243098
rect 242004 207418 242186 207654
rect 242422 207418 242604 207654
rect 242004 207334 242604 207418
rect 242004 207098 242186 207334
rect 242422 207098 242604 207334
rect 241467 181116 241533 181117
rect 241467 181052 241468 181116
rect 241532 181052 241533 181116
rect 241467 181051 241533 181052
rect 241470 180845 241530 181051
rect 241467 180844 241533 180845
rect 241467 180780 241468 180844
rect 241532 180780 241533 180844
rect 241467 180779 241533 180780
rect 238404 167818 238586 168054
rect 238822 167818 239004 168054
rect 238404 167734 239004 167818
rect 238404 167498 238586 167734
rect 238822 167498 239004 167734
rect 238404 132054 239004 167498
rect 238404 131818 238586 132054
rect 238822 131818 239004 132054
rect 238404 131734 239004 131818
rect 238404 131498 238586 131734
rect 238822 131498 239004 131734
rect 238404 96054 239004 131498
rect 238404 95818 238586 96054
rect 238822 95818 239004 96054
rect 238404 95734 239004 95818
rect 238404 95498 238586 95734
rect 238822 95498 239004 95734
rect 238155 91220 238221 91221
rect 238155 91156 238156 91220
rect 238220 91156 238221 91220
rect 238155 91155 238221 91156
rect 237235 63612 237301 63613
rect 237235 63548 237236 63612
rect 237300 63548 237301 63612
rect 237235 63547 237301 63548
rect 234804 56218 234986 56454
rect 235222 56218 235404 56454
rect 234804 56134 235404 56218
rect 234804 55898 234986 56134
rect 235222 55898 235404 56134
rect 234475 32604 234541 32605
rect 234475 32540 234476 32604
rect 234540 32540 234541 32604
rect 234475 32539 234541 32540
rect 234804 20454 235404 55898
rect 234804 20218 234986 20454
rect 235222 20218 235404 20454
rect 234804 20134 235404 20218
rect 234804 19898 234986 20134
rect 235222 19898 235404 20134
rect 231715 16692 231781 16693
rect 231715 16628 231716 16692
rect 231780 16628 231781 16692
rect 231715 16627 231781 16628
rect 227604 13018 227786 13254
rect 228022 13018 228204 13254
rect 227604 12934 228204 13018
rect 227604 12698 227786 12934
rect 228022 12698 228204 12934
rect 209604 -7022 209786 -6786
rect 210022 -7022 210204 -6786
rect 209604 -7106 210204 -7022
rect 209604 -7342 209786 -7106
rect 210022 -7342 210204 -7106
rect 209604 -7364 210204 -7342
rect 227604 -5866 228204 12698
rect 234804 -1266 235404 19898
rect 234804 -1502 234986 -1266
rect 235222 -1502 235404 -1266
rect 234804 -1586 235404 -1502
rect 234804 -1822 234986 -1586
rect 235222 -1822 235404 -1586
rect 234804 -1844 235404 -1822
rect 238404 60054 239004 95498
rect 238404 59818 238586 60054
rect 238822 59818 239004 60054
rect 238404 59734 239004 59818
rect 238404 59498 238586 59734
rect 238822 59498 239004 59734
rect 238404 24054 239004 59498
rect 238404 23818 238586 24054
rect 238822 23818 239004 24054
rect 238404 23734 239004 23818
rect 238404 23498 238586 23734
rect 238822 23498 239004 23734
rect 238404 -3106 239004 23498
rect 238404 -3342 238586 -3106
rect 238822 -3342 239004 -3106
rect 238404 -3426 239004 -3342
rect 238404 -3662 238586 -3426
rect 238822 -3662 239004 -3426
rect 238404 -3684 239004 -3662
rect 242004 171654 242604 207098
rect 242004 171418 242186 171654
rect 242422 171418 242604 171654
rect 242004 171334 242604 171418
rect 242004 171098 242186 171334
rect 242422 171098 242604 171334
rect 242004 135654 242604 171098
rect 242004 135418 242186 135654
rect 242422 135418 242604 135654
rect 242004 135334 242604 135418
rect 242004 135098 242186 135334
rect 242422 135098 242604 135334
rect 242004 99654 242604 135098
rect 242004 99418 242186 99654
rect 242422 99418 242604 99654
rect 242004 99334 242604 99418
rect 242004 99098 242186 99334
rect 242422 99098 242604 99334
rect 242004 63654 242604 99098
rect 242004 63418 242186 63654
rect 242422 63418 242604 63654
rect 242004 63334 242604 63418
rect 242004 63098 242186 63334
rect 242422 63098 242604 63334
rect 242004 27654 242604 63098
rect 242004 27418 242186 27654
rect 242422 27418 242604 27654
rect 242004 27334 242604 27418
rect 242004 27098 242186 27334
rect 242422 27098 242604 27334
rect 242004 -4946 242604 27098
rect 242004 -5182 242186 -4946
rect 242422 -5182 242604 -4946
rect 242004 -5266 242604 -5182
rect 242004 -5502 242186 -5266
rect 242422 -5502 242604 -5266
rect 242004 -5524 242604 -5502
rect 245604 535254 246204 570698
rect 252804 704838 253404 705780
rect 252804 704602 252986 704838
rect 253222 704602 253404 704838
rect 252804 704518 253404 704602
rect 252804 704282 252986 704518
rect 253222 704282 253404 704518
rect 252804 686454 253404 704282
rect 252804 686218 252986 686454
rect 253222 686218 253404 686454
rect 252804 686134 253404 686218
rect 252804 685898 252986 686134
rect 253222 685898 253404 686134
rect 252804 650454 253404 685898
rect 252804 650218 252986 650454
rect 253222 650218 253404 650454
rect 252804 650134 253404 650218
rect 252804 649898 252986 650134
rect 253222 649898 253404 650134
rect 252804 614454 253404 649898
rect 252804 614218 252986 614454
rect 253222 614218 253404 614454
rect 252804 614134 253404 614218
rect 252804 613898 252986 614134
rect 253222 613898 253404 614134
rect 252804 578454 253404 613898
rect 252804 578218 252986 578454
rect 253222 578218 253404 578454
rect 252804 578134 253404 578218
rect 252804 577898 252986 578134
rect 253222 577898 253404 578134
rect 252507 563004 252573 563005
rect 252507 562940 252508 563004
rect 252572 562940 252573 563004
rect 252507 562939 252573 562940
rect 252510 562138 252570 562939
rect 252507 559196 252573 559197
rect 252507 559132 252508 559196
rect 252572 559132 252573 559196
rect 252507 559131 252573 559132
rect 252510 558789 252570 559131
rect 252507 558788 252573 558789
rect 252507 558724 252508 558788
rect 252572 558724 252573 558788
rect 252507 558723 252573 558724
rect 245604 535018 245786 535254
rect 246022 535018 246204 535254
rect 245604 534934 246204 535018
rect 245604 534698 245786 534934
rect 246022 534698 246204 534934
rect 245604 499254 246204 534698
rect 245604 499018 245786 499254
rect 246022 499018 246204 499254
rect 245604 498934 246204 499018
rect 245604 498698 245786 498934
rect 246022 498698 246204 498934
rect 245604 463254 246204 498698
rect 245604 463018 245786 463254
rect 246022 463018 246204 463254
rect 245604 462934 246204 463018
rect 245604 462698 245786 462934
rect 246022 462698 246204 462934
rect 245604 427254 246204 462698
rect 245604 427018 245786 427254
rect 246022 427018 246204 427254
rect 245604 426934 246204 427018
rect 245604 426698 245786 426934
rect 246022 426698 246204 426934
rect 245604 391254 246204 426698
rect 245604 391018 245786 391254
rect 246022 391018 246204 391254
rect 245604 390934 246204 391018
rect 245604 390698 245786 390934
rect 246022 390698 246204 390934
rect 245604 355254 246204 390698
rect 245604 355018 245786 355254
rect 246022 355018 246204 355254
rect 245604 354934 246204 355018
rect 245604 354698 245786 354934
rect 246022 354698 246204 354934
rect 245604 319254 246204 354698
rect 245604 319018 245786 319254
rect 246022 319018 246204 319254
rect 245604 318934 246204 319018
rect 245604 318698 245786 318934
rect 246022 318698 246204 318934
rect 245604 283254 246204 318698
rect 245604 283018 245786 283254
rect 246022 283018 246204 283254
rect 245604 282934 246204 283018
rect 245604 282698 245786 282934
rect 246022 282698 246204 282934
rect 245604 247254 246204 282698
rect 245604 247018 245786 247254
rect 246022 247018 246204 247254
rect 245604 246934 246204 247018
rect 245604 246698 245786 246934
rect 246022 246698 246204 246934
rect 245604 211254 246204 246698
rect 245604 211018 245786 211254
rect 246022 211018 246204 211254
rect 245604 210934 246204 211018
rect 245604 210698 245786 210934
rect 246022 210698 246204 210934
rect 245604 175254 246204 210698
rect 245604 175018 245786 175254
rect 246022 175018 246204 175254
rect 245604 174934 246204 175018
rect 245604 174698 245786 174934
rect 246022 174698 246204 174934
rect 245604 139254 246204 174698
rect 245604 139018 245786 139254
rect 246022 139018 246204 139254
rect 245604 138934 246204 139018
rect 245604 138698 245786 138934
rect 246022 138698 246204 138934
rect 245604 103254 246204 138698
rect 245604 103018 245786 103254
rect 246022 103018 246204 103254
rect 245604 102934 246204 103018
rect 245604 102698 245786 102934
rect 246022 102698 246204 102934
rect 245604 67254 246204 102698
rect 245604 67018 245786 67254
rect 246022 67018 246204 67254
rect 245604 66934 246204 67018
rect 245604 66698 245786 66934
rect 246022 66698 246204 66934
rect 245604 31254 246204 66698
rect 252804 542454 253404 577898
rect 256404 690054 257004 706122
rect 256404 689818 256586 690054
rect 256822 689818 257004 690054
rect 256404 689734 257004 689818
rect 256404 689498 256586 689734
rect 256822 689498 257004 689734
rect 256404 654054 257004 689498
rect 256404 653818 256586 654054
rect 256822 653818 257004 654054
rect 256404 653734 257004 653818
rect 256404 653498 256586 653734
rect 256822 653498 257004 653734
rect 256404 618054 257004 653498
rect 256404 617818 256586 618054
rect 256822 617818 257004 618054
rect 256404 617734 257004 617818
rect 256404 617498 256586 617734
rect 256822 617498 257004 617734
rect 256404 582054 257004 617498
rect 256404 581818 256586 582054
rect 256822 581818 257004 582054
rect 256404 581734 257004 581818
rect 256404 581498 256586 581734
rect 256822 581498 257004 581734
rect 253611 563004 253677 563005
rect 253611 562940 253612 563004
rect 253676 562940 253677 563004
rect 253611 562939 253677 562940
rect 253614 562818 253674 562939
rect 252804 542218 252986 542454
rect 253222 542218 253404 542454
rect 252804 542134 253404 542218
rect 252804 541898 252986 542134
rect 253222 541898 253404 542134
rect 252804 506454 253404 541898
rect 252804 506218 252986 506454
rect 253222 506218 253404 506454
rect 252804 506134 253404 506218
rect 252804 505898 252986 506134
rect 253222 505898 253404 506134
rect 252804 470454 253404 505898
rect 252804 470218 252986 470454
rect 253222 470218 253404 470454
rect 252804 470134 253404 470218
rect 252804 469898 252986 470134
rect 253222 469898 253404 470134
rect 252804 434454 253404 469898
rect 252804 434218 252986 434454
rect 253222 434218 253404 434454
rect 252804 434134 253404 434218
rect 252804 433898 252986 434134
rect 253222 433898 253404 434134
rect 252804 398454 253404 433898
rect 252804 398218 252986 398454
rect 253222 398218 253404 398454
rect 252804 398134 253404 398218
rect 252804 397898 252986 398134
rect 253222 397898 253404 398134
rect 252804 362454 253404 397898
rect 252804 362218 252986 362454
rect 253222 362218 253404 362454
rect 252804 362134 253404 362218
rect 252804 361898 252986 362134
rect 253222 361898 253404 362134
rect 252804 326454 253404 361898
rect 252804 326218 252986 326454
rect 253222 326218 253404 326454
rect 252804 326134 253404 326218
rect 252804 325898 252986 326134
rect 253222 325898 253404 326134
rect 252804 290454 253404 325898
rect 252804 290218 252986 290454
rect 253222 290218 253404 290454
rect 252804 290134 253404 290218
rect 252804 289898 252986 290134
rect 253222 289898 253404 290134
rect 252804 254454 253404 289898
rect 252804 254218 252986 254454
rect 253222 254218 253404 254454
rect 252804 254134 253404 254218
rect 252804 253898 252986 254134
rect 253222 253898 253404 254134
rect 252804 218454 253404 253898
rect 252804 218218 252986 218454
rect 253222 218218 253404 218454
rect 252804 218134 253404 218218
rect 252804 217898 252986 218134
rect 253222 217898 253404 218134
rect 252804 182454 253404 217898
rect 252804 182218 252986 182454
rect 253222 182218 253404 182454
rect 252804 182134 253404 182218
rect 252804 181898 252986 182134
rect 253222 181898 253404 182134
rect 252804 146454 253404 181898
rect 252804 146218 252986 146454
rect 253222 146218 253404 146454
rect 252804 146134 253404 146218
rect 252804 145898 252986 146134
rect 253222 145898 253404 146134
rect 252804 110454 253404 145898
rect 252804 110218 252986 110454
rect 253222 110218 253404 110454
rect 252804 110134 253404 110218
rect 252804 109898 252986 110134
rect 253222 109898 253404 110134
rect 252804 74454 253404 109898
rect 252804 74218 252986 74454
rect 253222 74218 253404 74454
rect 252804 74134 253404 74218
rect 252804 73898 252986 74134
rect 253222 73898 253404 74134
rect 249747 40356 249813 40357
rect 249747 40292 249748 40356
rect 249812 40292 249813 40356
rect 249747 40291 249813 40292
rect 249750 40085 249810 40291
rect 249747 40084 249813 40085
rect 249747 40020 249748 40084
rect 249812 40020 249813 40084
rect 249747 40019 249813 40020
rect 245604 31018 245786 31254
rect 246022 31018 246204 31254
rect 245604 30934 246204 31018
rect 245604 30698 245786 30934
rect 246022 30698 246204 30934
rect 227604 -6102 227786 -5866
rect 228022 -6102 228204 -5866
rect 227604 -6186 228204 -6102
rect 227604 -6422 227786 -6186
rect 228022 -6422 228204 -6186
rect 227604 -7364 228204 -6422
rect 245604 -6786 246204 30698
rect 252804 38454 253404 73898
rect 252804 38218 252986 38454
rect 253222 38218 253404 38454
rect 252804 38134 253404 38218
rect 252804 37898 252986 38134
rect 253222 37898 253404 38134
rect 252804 2454 253404 37898
rect 252804 2218 252986 2454
rect 253222 2218 253404 2454
rect 252804 2134 253404 2218
rect 252804 1898 252986 2134
rect 253222 1898 253404 2134
rect 252804 -346 253404 1898
rect 252804 -582 252986 -346
rect 253222 -582 253404 -346
rect 252804 -666 253404 -582
rect 252804 -902 252986 -666
rect 253222 -902 253404 -666
rect 252804 -1844 253404 -902
rect 256404 546054 257004 581498
rect 256404 545818 256586 546054
rect 256822 545818 257004 546054
rect 256404 545734 257004 545818
rect 256404 545498 256586 545734
rect 256822 545498 257004 545734
rect 256404 510054 257004 545498
rect 256404 509818 256586 510054
rect 256822 509818 257004 510054
rect 256404 509734 257004 509818
rect 256404 509498 256586 509734
rect 256822 509498 257004 509734
rect 256404 474054 257004 509498
rect 256404 473818 256586 474054
rect 256822 473818 257004 474054
rect 256404 473734 257004 473818
rect 256404 473498 256586 473734
rect 256822 473498 257004 473734
rect 256404 438054 257004 473498
rect 256404 437818 256586 438054
rect 256822 437818 257004 438054
rect 256404 437734 257004 437818
rect 256404 437498 256586 437734
rect 256822 437498 257004 437734
rect 256404 402054 257004 437498
rect 256404 401818 256586 402054
rect 256822 401818 257004 402054
rect 256404 401734 257004 401818
rect 256404 401498 256586 401734
rect 256822 401498 257004 401734
rect 256404 366054 257004 401498
rect 256404 365818 256586 366054
rect 256822 365818 257004 366054
rect 256404 365734 257004 365818
rect 256404 365498 256586 365734
rect 256822 365498 257004 365734
rect 256404 330054 257004 365498
rect 256404 329818 256586 330054
rect 256822 329818 257004 330054
rect 256404 329734 257004 329818
rect 256404 329498 256586 329734
rect 256822 329498 257004 329734
rect 256404 294054 257004 329498
rect 256404 293818 256586 294054
rect 256822 293818 257004 294054
rect 256404 293734 257004 293818
rect 256404 293498 256586 293734
rect 256822 293498 257004 293734
rect 256404 258054 257004 293498
rect 256404 257818 256586 258054
rect 256822 257818 257004 258054
rect 256404 257734 257004 257818
rect 256404 257498 256586 257734
rect 256822 257498 257004 257734
rect 256404 222054 257004 257498
rect 256404 221818 256586 222054
rect 256822 221818 257004 222054
rect 256404 221734 257004 221818
rect 256404 221498 256586 221734
rect 256822 221498 257004 221734
rect 256404 186054 257004 221498
rect 256404 185818 256586 186054
rect 256822 185818 257004 186054
rect 256404 185734 257004 185818
rect 256404 185498 256586 185734
rect 256822 185498 257004 185734
rect 256404 150054 257004 185498
rect 256404 149818 256586 150054
rect 256822 149818 257004 150054
rect 256404 149734 257004 149818
rect 256404 149498 256586 149734
rect 256822 149498 257004 149734
rect 256404 114054 257004 149498
rect 256404 113818 256586 114054
rect 256822 113818 257004 114054
rect 256404 113734 257004 113818
rect 256404 113498 256586 113734
rect 256822 113498 257004 113734
rect 256404 78054 257004 113498
rect 256404 77818 256586 78054
rect 256822 77818 257004 78054
rect 256404 77734 257004 77818
rect 256404 77498 256586 77734
rect 256822 77498 257004 77734
rect 256404 42054 257004 77498
rect 256404 41818 256586 42054
rect 256822 41818 257004 42054
rect 256404 41734 257004 41818
rect 256404 41498 256586 41734
rect 256822 41498 257004 41734
rect 256404 6054 257004 41498
rect 256404 5818 256586 6054
rect 256822 5818 257004 6054
rect 256404 5734 257004 5818
rect 256404 5498 256586 5734
rect 256822 5498 257004 5734
rect 256404 -2186 257004 5498
rect 256404 -2422 256586 -2186
rect 256822 -2422 257004 -2186
rect 256404 -2506 257004 -2422
rect 256404 -2742 256586 -2506
rect 256822 -2742 257004 -2506
rect 256404 -3684 257004 -2742
rect 260004 693654 260604 707962
rect 260004 693418 260186 693654
rect 260422 693418 260604 693654
rect 260004 693334 260604 693418
rect 260004 693098 260186 693334
rect 260422 693098 260604 693334
rect 260004 657654 260604 693098
rect 260004 657418 260186 657654
rect 260422 657418 260604 657654
rect 260004 657334 260604 657418
rect 260004 657098 260186 657334
rect 260422 657098 260604 657334
rect 260004 621654 260604 657098
rect 260004 621418 260186 621654
rect 260422 621418 260604 621654
rect 260004 621334 260604 621418
rect 260004 621098 260186 621334
rect 260422 621098 260604 621334
rect 260004 585654 260604 621098
rect 260004 585418 260186 585654
rect 260422 585418 260604 585654
rect 260004 585334 260604 585418
rect 260004 585098 260186 585334
rect 260422 585098 260604 585334
rect 260004 549654 260604 585098
rect 260004 549418 260186 549654
rect 260422 549418 260604 549654
rect 260004 549334 260604 549418
rect 260004 549098 260186 549334
rect 260422 549098 260604 549334
rect 260004 513654 260604 549098
rect 260004 513418 260186 513654
rect 260422 513418 260604 513654
rect 260004 513334 260604 513418
rect 260004 513098 260186 513334
rect 260422 513098 260604 513334
rect 260004 477654 260604 513098
rect 260004 477418 260186 477654
rect 260422 477418 260604 477654
rect 260004 477334 260604 477418
rect 260004 477098 260186 477334
rect 260422 477098 260604 477334
rect 260004 441654 260604 477098
rect 260004 441418 260186 441654
rect 260422 441418 260604 441654
rect 260004 441334 260604 441418
rect 260004 441098 260186 441334
rect 260422 441098 260604 441334
rect 260004 405654 260604 441098
rect 260004 405418 260186 405654
rect 260422 405418 260604 405654
rect 260004 405334 260604 405418
rect 260004 405098 260186 405334
rect 260422 405098 260604 405334
rect 260004 369654 260604 405098
rect 260004 369418 260186 369654
rect 260422 369418 260604 369654
rect 260004 369334 260604 369418
rect 260004 369098 260186 369334
rect 260422 369098 260604 369334
rect 260004 333654 260604 369098
rect 260004 333418 260186 333654
rect 260422 333418 260604 333654
rect 260004 333334 260604 333418
rect 260004 333098 260186 333334
rect 260422 333098 260604 333334
rect 260004 297654 260604 333098
rect 260004 297418 260186 297654
rect 260422 297418 260604 297654
rect 260004 297334 260604 297418
rect 260004 297098 260186 297334
rect 260422 297098 260604 297334
rect 260004 261654 260604 297098
rect 260004 261418 260186 261654
rect 260422 261418 260604 261654
rect 260004 261334 260604 261418
rect 260004 261098 260186 261334
rect 260422 261098 260604 261334
rect 260004 225654 260604 261098
rect 260004 225418 260186 225654
rect 260422 225418 260604 225654
rect 260004 225334 260604 225418
rect 260004 225098 260186 225334
rect 260422 225098 260604 225334
rect 260004 189654 260604 225098
rect 260004 189418 260186 189654
rect 260422 189418 260604 189654
rect 260004 189334 260604 189418
rect 260004 189098 260186 189334
rect 260422 189098 260604 189334
rect 260004 153654 260604 189098
rect 260004 153418 260186 153654
rect 260422 153418 260604 153654
rect 260004 153334 260604 153418
rect 260004 153098 260186 153334
rect 260422 153098 260604 153334
rect 260004 117654 260604 153098
rect 260004 117418 260186 117654
rect 260422 117418 260604 117654
rect 260004 117334 260604 117418
rect 260004 117098 260186 117334
rect 260422 117098 260604 117334
rect 260004 81654 260604 117098
rect 260004 81418 260186 81654
rect 260422 81418 260604 81654
rect 260004 81334 260604 81418
rect 260004 81098 260186 81334
rect 260422 81098 260604 81334
rect 260004 45654 260604 81098
rect 260004 45418 260186 45654
rect 260422 45418 260604 45654
rect 260004 45334 260604 45418
rect 260004 45098 260186 45334
rect 260422 45098 260604 45334
rect 260004 9654 260604 45098
rect 260004 9418 260186 9654
rect 260422 9418 260604 9654
rect 260004 9334 260604 9418
rect 260004 9098 260186 9334
rect 260422 9098 260604 9334
rect 260004 -4026 260604 9098
rect 260004 -4262 260186 -4026
rect 260422 -4262 260604 -4026
rect 260004 -4346 260604 -4262
rect 260004 -4582 260186 -4346
rect 260422 -4582 260604 -4346
rect 260004 -5524 260604 -4582
rect 263604 697254 264204 709802
rect 281604 711278 282204 711300
rect 281604 711042 281786 711278
rect 282022 711042 282204 711278
rect 281604 710958 282204 711042
rect 281604 710722 281786 710958
rect 282022 710722 282204 710958
rect 278004 709438 278604 709460
rect 278004 709202 278186 709438
rect 278422 709202 278604 709438
rect 278004 709118 278604 709202
rect 278004 708882 278186 709118
rect 278422 708882 278604 709118
rect 274404 707598 275004 707620
rect 274404 707362 274586 707598
rect 274822 707362 275004 707598
rect 274404 707278 275004 707362
rect 274404 707042 274586 707278
rect 274822 707042 275004 707278
rect 263604 697018 263786 697254
rect 264022 697018 264204 697254
rect 263604 696934 264204 697018
rect 263604 696698 263786 696934
rect 264022 696698 264204 696934
rect 263604 661254 264204 696698
rect 263604 661018 263786 661254
rect 264022 661018 264204 661254
rect 263604 660934 264204 661018
rect 263604 660698 263786 660934
rect 264022 660698 264204 660934
rect 263604 625254 264204 660698
rect 263604 625018 263786 625254
rect 264022 625018 264204 625254
rect 263604 624934 264204 625018
rect 263604 624698 263786 624934
rect 264022 624698 264204 624934
rect 263604 589254 264204 624698
rect 263604 589018 263786 589254
rect 264022 589018 264204 589254
rect 263604 588934 264204 589018
rect 263604 588698 263786 588934
rect 264022 588698 264204 588934
rect 263604 553254 264204 588698
rect 270804 705758 271404 705780
rect 270804 705522 270986 705758
rect 271222 705522 271404 705758
rect 270804 705438 271404 705522
rect 270804 705202 270986 705438
rect 271222 705202 271404 705438
rect 270804 668454 271404 705202
rect 270804 668218 270986 668454
rect 271222 668218 271404 668454
rect 270804 668134 271404 668218
rect 270804 667898 270986 668134
rect 271222 667898 271404 668134
rect 270804 632454 271404 667898
rect 270804 632218 270986 632454
rect 271222 632218 271404 632454
rect 270804 632134 271404 632218
rect 270804 631898 270986 632134
rect 271222 631898 271404 632134
rect 270804 596454 271404 631898
rect 270804 596218 270986 596454
rect 271222 596218 271404 596454
rect 270804 596134 271404 596218
rect 270804 595898 270986 596134
rect 271222 595898 271404 596134
rect 266307 563004 266373 563005
rect 266307 562940 266308 563004
rect 266372 562940 266373 563004
rect 266307 562939 266373 562940
rect 266310 562138 266370 562939
rect 263604 553018 263786 553254
rect 264022 553018 264204 553254
rect 263604 552934 264204 553018
rect 263604 552698 263786 552934
rect 264022 552698 264204 552934
rect 263604 517254 264204 552698
rect 263604 517018 263786 517254
rect 264022 517018 264204 517254
rect 263604 516934 264204 517018
rect 263604 516698 263786 516934
rect 264022 516698 264204 516934
rect 263604 481254 264204 516698
rect 263604 481018 263786 481254
rect 264022 481018 264204 481254
rect 263604 480934 264204 481018
rect 263604 480698 263786 480934
rect 264022 480698 264204 480934
rect 263604 445254 264204 480698
rect 263604 445018 263786 445254
rect 264022 445018 264204 445254
rect 263604 444934 264204 445018
rect 263604 444698 263786 444934
rect 264022 444698 264204 444934
rect 263604 409254 264204 444698
rect 263604 409018 263786 409254
rect 264022 409018 264204 409254
rect 263604 408934 264204 409018
rect 263604 408698 263786 408934
rect 264022 408698 264204 408934
rect 263604 373254 264204 408698
rect 263604 373018 263786 373254
rect 264022 373018 264204 373254
rect 263604 372934 264204 373018
rect 263604 372698 263786 372934
rect 264022 372698 264204 372934
rect 263604 337254 264204 372698
rect 263604 337018 263786 337254
rect 264022 337018 264204 337254
rect 263604 336934 264204 337018
rect 263604 336698 263786 336934
rect 264022 336698 264204 336934
rect 263604 301254 264204 336698
rect 263604 301018 263786 301254
rect 264022 301018 264204 301254
rect 263604 300934 264204 301018
rect 263604 300698 263786 300934
rect 264022 300698 264204 300934
rect 263604 265254 264204 300698
rect 263604 265018 263786 265254
rect 264022 265018 264204 265254
rect 263604 264934 264204 265018
rect 263604 264698 263786 264934
rect 264022 264698 264204 264934
rect 263604 229254 264204 264698
rect 263604 229018 263786 229254
rect 264022 229018 264204 229254
rect 263604 228934 264204 229018
rect 263604 228698 263786 228934
rect 264022 228698 264204 228934
rect 263604 193254 264204 228698
rect 263604 193018 263786 193254
rect 264022 193018 264204 193254
rect 263604 192934 264204 193018
rect 263604 192698 263786 192934
rect 264022 192698 264204 192934
rect 263604 157254 264204 192698
rect 263604 157018 263786 157254
rect 264022 157018 264204 157254
rect 263604 156934 264204 157018
rect 263604 156698 263786 156934
rect 264022 156698 264204 156934
rect 263604 121254 264204 156698
rect 263604 121018 263786 121254
rect 264022 121018 264204 121254
rect 263604 120934 264204 121018
rect 263604 120698 263786 120934
rect 264022 120698 264204 120934
rect 263604 85254 264204 120698
rect 270804 560454 271404 595898
rect 270804 560218 270986 560454
rect 271222 560218 271404 560454
rect 270804 560134 271404 560218
rect 270804 559898 270986 560134
rect 271222 559898 271404 560134
rect 270804 524454 271404 559898
rect 270804 524218 270986 524454
rect 271222 524218 271404 524454
rect 270804 524134 271404 524218
rect 270804 523898 270986 524134
rect 271222 523898 271404 524134
rect 270804 488454 271404 523898
rect 270804 488218 270986 488454
rect 271222 488218 271404 488454
rect 270804 488134 271404 488218
rect 270804 487898 270986 488134
rect 271222 487898 271404 488134
rect 270804 452454 271404 487898
rect 270804 452218 270986 452454
rect 271222 452218 271404 452454
rect 270804 452134 271404 452218
rect 270804 451898 270986 452134
rect 271222 451898 271404 452134
rect 270804 416454 271404 451898
rect 270804 416218 270986 416454
rect 271222 416218 271404 416454
rect 270804 416134 271404 416218
rect 270804 415898 270986 416134
rect 271222 415898 271404 416134
rect 270804 380454 271404 415898
rect 270804 380218 270986 380454
rect 271222 380218 271404 380454
rect 270804 380134 271404 380218
rect 270804 379898 270986 380134
rect 271222 379898 271404 380134
rect 270804 344454 271404 379898
rect 270804 344218 270986 344454
rect 271222 344218 271404 344454
rect 270804 344134 271404 344218
rect 270804 343898 270986 344134
rect 271222 343898 271404 344134
rect 270804 308454 271404 343898
rect 270804 308218 270986 308454
rect 271222 308218 271404 308454
rect 270804 308134 271404 308218
rect 270804 307898 270986 308134
rect 271222 307898 271404 308134
rect 270804 272454 271404 307898
rect 270804 272218 270986 272454
rect 271222 272218 271404 272454
rect 270804 272134 271404 272218
rect 270804 271898 270986 272134
rect 271222 271898 271404 272134
rect 270804 236454 271404 271898
rect 270804 236218 270986 236454
rect 271222 236218 271404 236454
rect 270804 236134 271404 236218
rect 270804 235898 270986 236134
rect 271222 235898 271404 236134
rect 270804 200454 271404 235898
rect 270804 200218 270986 200454
rect 271222 200218 271404 200454
rect 270804 200134 271404 200218
rect 270804 199898 270986 200134
rect 271222 199898 271404 200134
rect 270804 164454 271404 199898
rect 270804 164218 270986 164454
rect 271222 164218 271404 164454
rect 270804 164134 271404 164218
rect 270804 163898 270986 164134
rect 271222 163898 271404 164134
rect 270804 128454 271404 163898
rect 270804 128218 270986 128454
rect 271222 128218 271404 128454
rect 270804 128134 271404 128218
rect 270804 127898 270986 128134
rect 271222 127898 271404 128134
rect 270804 92454 271404 127898
rect 270804 92218 270986 92454
rect 271222 92218 271404 92454
rect 270804 92134 271404 92218
rect 270804 91898 270986 92134
rect 271222 91898 271404 92134
rect 269067 87276 269133 87277
rect 269067 87212 269068 87276
rect 269132 87212 269133 87276
rect 269067 87211 269133 87212
rect 269070 87005 269130 87211
rect 269067 87004 269133 87005
rect 269067 86940 269068 87004
rect 269132 86940 269133 87004
rect 269067 86939 269133 86940
rect 263604 85018 263786 85254
rect 264022 85018 264204 85254
rect 263604 84934 264204 85018
rect 263604 84698 263786 84934
rect 264022 84698 264204 84934
rect 263604 49254 264204 84698
rect 263604 49018 263786 49254
rect 264022 49018 264204 49254
rect 263604 48934 264204 49018
rect 263604 48698 263786 48934
rect 264022 48698 264204 48934
rect 263604 13254 264204 48698
rect 263604 13018 263786 13254
rect 264022 13018 264204 13254
rect 263604 12934 264204 13018
rect 263604 12698 263786 12934
rect 264022 12698 264204 12934
rect 245604 -7022 245786 -6786
rect 246022 -7022 246204 -6786
rect 245604 -7106 246204 -7022
rect 245604 -7342 245786 -7106
rect 246022 -7342 246204 -7106
rect 245604 -7364 246204 -7342
rect 263604 -5866 264204 12698
rect 270804 56454 271404 91898
rect 270804 56218 270986 56454
rect 271222 56218 271404 56454
rect 270804 56134 271404 56218
rect 270804 55898 270986 56134
rect 271222 55898 271404 56134
rect 270804 20454 271404 55898
rect 270804 20218 270986 20454
rect 271222 20218 271404 20454
rect 270804 20134 271404 20218
rect 270804 19898 270986 20134
rect 271222 19898 271404 20134
rect 270804 -1266 271404 19898
rect 270804 -1502 270986 -1266
rect 271222 -1502 271404 -1266
rect 270804 -1586 271404 -1502
rect 270804 -1822 270986 -1586
rect 271222 -1822 271404 -1586
rect 270804 -1844 271404 -1822
rect 274404 672054 275004 707042
rect 274404 671818 274586 672054
rect 274822 671818 275004 672054
rect 274404 671734 275004 671818
rect 274404 671498 274586 671734
rect 274822 671498 275004 671734
rect 274404 636054 275004 671498
rect 274404 635818 274586 636054
rect 274822 635818 275004 636054
rect 274404 635734 275004 635818
rect 274404 635498 274586 635734
rect 274822 635498 275004 635734
rect 274404 600054 275004 635498
rect 274404 599818 274586 600054
rect 274822 599818 275004 600054
rect 274404 599734 275004 599818
rect 274404 599498 274586 599734
rect 274822 599498 275004 599734
rect 274404 564054 275004 599498
rect 274404 563818 274586 564054
rect 274822 563818 275004 564054
rect 274404 563734 275004 563818
rect 274404 563498 274586 563734
rect 274822 563498 275004 563734
rect 274404 528054 275004 563498
rect 278004 675654 278604 708882
rect 278004 675418 278186 675654
rect 278422 675418 278604 675654
rect 278004 675334 278604 675418
rect 278004 675098 278186 675334
rect 278422 675098 278604 675334
rect 278004 639654 278604 675098
rect 278004 639418 278186 639654
rect 278422 639418 278604 639654
rect 278004 639334 278604 639418
rect 278004 639098 278186 639334
rect 278422 639098 278604 639334
rect 278004 603654 278604 639098
rect 278004 603418 278186 603654
rect 278422 603418 278604 603654
rect 278004 603334 278604 603418
rect 278004 603098 278186 603334
rect 278422 603098 278604 603334
rect 278004 567654 278604 603098
rect 278004 567418 278186 567654
rect 278422 567418 278604 567654
rect 278004 567334 278604 567418
rect 278004 567098 278186 567334
rect 278422 567098 278604 567334
rect 275875 563004 275941 563005
rect 275875 562940 275876 563004
rect 275940 562940 275941 563004
rect 275875 562939 275941 562940
rect 275878 562818 275938 562939
rect 274404 527818 274586 528054
rect 274822 527818 275004 528054
rect 274404 527734 275004 527818
rect 274404 527498 274586 527734
rect 274822 527498 275004 527734
rect 274404 492054 275004 527498
rect 274404 491818 274586 492054
rect 274822 491818 275004 492054
rect 274404 491734 275004 491818
rect 274404 491498 274586 491734
rect 274822 491498 275004 491734
rect 274404 456054 275004 491498
rect 274404 455818 274586 456054
rect 274822 455818 275004 456054
rect 274404 455734 275004 455818
rect 274404 455498 274586 455734
rect 274822 455498 275004 455734
rect 274404 420054 275004 455498
rect 274404 419818 274586 420054
rect 274822 419818 275004 420054
rect 274404 419734 275004 419818
rect 274404 419498 274586 419734
rect 274822 419498 275004 419734
rect 274404 384054 275004 419498
rect 274404 383818 274586 384054
rect 274822 383818 275004 384054
rect 274404 383734 275004 383818
rect 274404 383498 274586 383734
rect 274822 383498 275004 383734
rect 274404 348054 275004 383498
rect 274404 347818 274586 348054
rect 274822 347818 275004 348054
rect 274404 347734 275004 347818
rect 274404 347498 274586 347734
rect 274822 347498 275004 347734
rect 274404 312054 275004 347498
rect 274404 311818 274586 312054
rect 274822 311818 275004 312054
rect 274404 311734 275004 311818
rect 274404 311498 274586 311734
rect 274822 311498 275004 311734
rect 274404 276054 275004 311498
rect 274404 275818 274586 276054
rect 274822 275818 275004 276054
rect 274404 275734 275004 275818
rect 274404 275498 274586 275734
rect 274822 275498 275004 275734
rect 274404 240054 275004 275498
rect 274404 239818 274586 240054
rect 274822 239818 275004 240054
rect 274404 239734 275004 239818
rect 274404 239498 274586 239734
rect 274822 239498 275004 239734
rect 274404 204054 275004 239498
rect 274404 203818 274586 204054
rect 274822 203818 275004 204054
rect 274404 203734 275004 203818
rect 274404 203498 274586 203734
rect 274822 203498 275004 203734
rect 274404 168054 275004 203498
rect 274404 167818 274586 168054
rect 274822 167818 275004 168054
rect 274404 167734 275004 167818
rect 274404 167498 274586 167734
rect 274822 167498 275004 167734
rect 274404 132054 275004 167498
rect 274404 131818 274586 132054
rect 274822 131818 275004 132054
rect 274404 131734 275004 131818
rect 274404 131498 274586 131734
rect 274822 131498 275004 131734
rect 274404 96054 275004 131498
rect 274404 95818 274586 96054
rect 274822 95818 275004 96054
rect 274404 95734 275004 95818
rect 274404 95498 274586 95734
rect 274822 95498 275004 95734
rect 274404 60054 275004 95498
rect 274404 59818 274586 60054
rect 274822 59818 275004 60054
rect 274404 59734 275004 59818
rect 274404 59498 274586 59734
rect 274822 59498 275004 59734
rect 274404 24054 275004 59498
rect 274404 23818 274586 24054
rect 274822 23818 275004 24054
rect 274404 23734 275004 23818
rect 274404 23498 274586 23734
rect 274822 23498 275004 23734
rect 274404 -3106 275004 23498
rect 274404 -3342 274586 -3106
rect 274822 -3342 275004 -3106
rect 274404 -3426 275004 -3342
rect 274404 -3662 274586 -3426
rect 274822 -3662 275004 -3426
rect 274404 -3684 275004 -3662
rect 278004 531654 278604 567098
rect 281604 679254 282204 710722
rect 299604 710358 300204 711300
rect 299604 710122 299786 710358
rect 300022 710122 300204 710358
rect 299604 710038 300204 710122
rect 299604 709802 299786 710038
rect 300022 709802 300204 710038
rect 296004 708518 296604 709460
rect 296004 708282 296186 708518
rect 296422 708282 296604 708518
rect 296004 708198 296604 708282
rect 296004 707962 296186 708198
rect 296422 707962 296604 708198
rect 292404 706678 293004 707620
rect 292404 706442 292586 706678
rect 292822 706442 293004 706678
rect 292404 706358 293004 706442
rect 292404 706122 292586 706358
rect 292822 706122 293004 706358
rect 281604 679018 281786 679254
rect 282022 679018 282204 679254
rect 281604 678934 282204 679018
rect 281604 678698 281786 678934
rect 282022 678698 282204 678934
rect 281604 643254 282204 678698
rect 281604 643018 281786 643254
rect 282022 643018 282204 643254
rect 281604 642934 282204 643018
rect 281604 642698 281786 642934
rect 282022 642698 282204 642934
rect 281604 607254 282204 642698
rect 281604 607018 281786 607254
rect 282022 607018 282204 607254
rect 281604 606934 282204 607018
rect 281604 606698 281786 606934
rect 282022 606698 282204 606934
rect 281604 571254 282204 606698
rect 281604 571018 281786 571254
rect 282022 571018 282204 571254
rect 281604 570934 282204 571018
rect 281604 570698 281786 570934
rect 282022 570698 282204 570934
rect 280107 560828 280173 560829
rect 280107 560764 280108 560828
rect 280172 560764 280173 560828
rect 280107 560763 280173 560764
rect 280110 560557 280170 560763
rect 280107 560556 280173 560557
rect 280107 560492 280108 560556
rect 280172 560492 280173 560556
rect 280107 560491 280173 560492
rect 278004 531418 278186 531654
rect 278422 531418 278604 531654
rect 278004 531334 278604 531418
rect 278004 531098 278186 531334
rect 278422 531098 278604 531334
rect 278004 495654 278604 531098
rect 278004 495418 278186 495654
rect 278422 495418 278604 495654
rect 278004 495334 278604 495418
rect 278004 495098 278186 495334
rect 278422 495098 278604 495334
rect 278004 459654 278604 495098
rect 278004 459418 278186 459654
rect 278422 459418 278604 459654
rect 278004 459334 278604 459418
rect 278004 459098 278186 459334
rect 278422 459098 278604 459334
rect 278004 423654 278604 459098
rect 278004 423418 278186 423654
rect 278422 423418 278604 423654
rect 278004 423334 278604 423418
rect 278004 423098 278186 423334
rect 278422 423098 278604 423334
rect 278004 387654 278604 423098
rect 278004 387418 278186 387654
rect 278422 387418 278604 387654
rect 278004 387334 278604 387418
rect 278004 387098 278186 387334
rect 278422 387098 278604 387334
rect 278004 351654 278604 387098
rect 278004 351418 278186 351654
rect 278422 351418 278604 351654
rect 278004 351334 278604 351418
rect 278004 351098 278186 351334
rect 278422 351098 278604 351334
rect 278004 315654 278604 351098
rect 278004 315418 278186 315654
rect 278422 315418 278604 315654
rect 278004 315334 278604 315418
rect 278004 315098 278186 315334
rect 278422 315098 278604 315334
rect 278004 279654 278604 315098
rect 278004 279418 278186 279654
rect 278422 279418 278604 279654
rect 278004 279334 278604 279418
rect 278004 279098 278186 279334
rect 278422 279098 278604 279334
rect 278004 243654 278604 279098
rect 278004 243418 278186 243654
rect 278422 243418 278604 243654
rect 278004 243334 278604 243418
rect 278004 243098 278186 243334
rect 278422 243098 278604 243334
rect 278004 207654 278604 243098
rect 278004 207418 278186 207654
rect 278422 207418 278604 207654
rect 278004 207334 278604 207418
rect 278004 207098 278186 207334
rect 278422 207098 278604 207334
rect 278004 171654 278604 207098
rect 278004 171418 278186 171654
rect 278422 171418 278604 171654
rect 278004 171334 278604 171418
rect 278004 171098 278186 171334
rect 278422 171098 278604 171334
rect 278004 135654 278604 171098
rect 278004 135418 278186 135654
rect 278422 135418 278604 135654
rect 278004 135334 278604 135418
rect 278004 135098 278186 135334
rect 278422 135098 278604 135334
rect 278004 99654 278604 135098
rect 278004 99418 278186 99654
rect 278422 99418 278604 99654
rect 278004 99334 278604 99418
rect 278004 99098 278186 99334
rect 278422 99098 278604 99334
rect 278004 63654 278604 99098
rect 278004 63418 278186 63654
rect 278422 63418 278604 63654
rect 278004 63334 278604 63418
rect 278004 63098 278186 63334
rect 278422 63098 278604 63334
rect 278004 27654 278604 63098
rect 278004 27418 278186 27654
rect 278422 27418 278604 27654
rect 278004 27334 278604 27418
rect 278004 27098 278186 27334
rect 278422 27098 278604 27334
rect 278004 -4946 278604 27098
rect 278004 -5182 278186 -4946
rect 278422 -5182 278604 -4946
rect 278004 -5266 278604 -5182
rect 278004 -5502 278186 -5266
rect 278422 -5502 278604 -5266
rect 278004 -5524 278604 -5502
rect 281604 535254 282204 570698
rect 288804 704838 289404 705780
rect 288804 704602 288986 704838
rect 289222 704602 289404 704838
rect 288804 704518 289404 704602
rect 288804 704282 288986 704518
rect 289222 704282 289404 704518
rect 288804 686454 289404 704282
rect 288804 686218 288986 686454
rect 289222 686218 289404 686454
rect 288804 686134 289404 686218
rect 288804 685898 288986 686134
rect 289222 685898 289404 686134
rect 288804 650454 289404 685898
rect 288804 650218 288986 650454
rect 289222 650218 289404 650454
rect 288804 650134 289404 650218
rect 288804 649898 288986 650134
rect 289222 649898 289404 650134
rect 288804 614454 289404 649898
rect 288804 614218 288986 614454
rect 289222 614218 289404 614454
rect 288804 614134 289404 614218
rect 288804 613898 288986 614134
rect 289222 613898 289404 614134
rect 288804 578454 289404 613898
rect 288804 578218 288986 578454
rect 289222 578218 289404 578454
rect 288804 578134 289404 578218
rect 288804 577898 288986 578134
rect 289222 577898 289404 578134
rect 288390 561645 288450 561902
rect 288387 561644 288453 561645
rect 288387 561580 288388 561644
rect 288452 561580 288453 561644
rect 288387 561579 288453 561580
rect 281604 535018 281786 535254
rect 282022 535018 282204 535254
rect 281604 534934 282204 535018
rect 281604 534698 281786 534934
rect 282022 534698 282204 534934
rect 281604 499254 282204 534698
rect 281604 499018 281786 499254
rect 282022 499018 282204 499254
rect 281604 498934 282204 499018
rect 281604 498698 281786 498934
rect 282022 498698 282204 498934
rect 281604 463254 282204 498698
rect 281604 463018 281786 463254
rect 282022 463018 282204 463254
rect 281604 462934 282204 463018
rect 281604 462698 281786 462934
rect 282022 462698 282204 462934
rect 281604 427254 282204 462698
rect 281604 427018 281786 427254
rect 282022 427018 282204 427254
rect 281604 426934 282204 427018
rect 281604 426698 281786 426934
rect 282022 426698 282204 426934
rect 281604 391254 282204 426698
rect 281604 391018 281786 391254
rect 282022 391018 282204 391254
rect 281604 390934 282204 391018
rect 281604 390698 281786 390934
rect 282022 390698 282204 390934
rect 281604 355254 282204 390698
rect 281604 355018 281786 355254
rect 282022 355018 282204 355254
rect 281604 354934 282204 355018
rect 281604 354698 281786 354934
rect 282022 354698 282204 354934
rect 281604 319254 282204 354698
rect 281604 319018 281786 319254
rect 282022 319018 282204 319254
rect 281604 318934 282204 319018
rect 281604 318698 281786 318934
rect 282022 318698 282204 318934
rect 281604 283254 282204 318698
rect 281604 283018 281786 283254
rect 282022 283018 282204 283254
rect 281604 282934 282204 283018
rect 281604 282698 281786 282934
rect 282022 282698 282204 282934
rect 281604 247254 282204 282698
rect 281604 247018 281786 247254
rect 282022 247018 282204 247254
rect 281604 246934 282204 247018
rect 281604 246698 281786 246934
rect 282022 246698 282204 246934
rect 281604 211254 282204 246698
rect 281604 211018 281786 211254
rect 282022 211018 282204 211254
rect 281604 210934 282204 211018
rect 281604 210698 281786 210934
rect 282022 210698 282204 210934
rect 281604 175254 282204 210698
rect 281604 175018 281786 175254
rect 282022 175018 282204 175254
rect 281604 174934 282204 175018
rect 281604 174698 281786 174934
rect 282022 174698 282204 174934
rect 281604 139254 282204 174698
rect 281604 139018 281786 139254
rect 282022 139018 282204 139254
rect 281604 138934 282204 139018
rect 281604 138698 281786 138934
rect 282022 138698 282204 138934
rect 281604 103254 282204 138698
rect 281604 103018 281786 103254
rect 282022 103018 282204 103254
rect 281604 102934 282204 103018
rect 281604 102698 281786 102934
rect 282022 102698 282204 102934
rect 281604 67254 282204 102698
rect 281604 67018 281786 67254
rect 282022 67018 282204 67254
rect 281604 66934 282204 67018
rect 281604 66698 281786 66934
rect 282022 66698 282204 66934
rect 281604 31254 282204 66698
rect 281604 31018 281786 31254
rect 282022 31018 282204 31254
rect 281604 30934 282204 31018
rect 281604 30698 281786 30934
rect 282022 30698 282204 30934
rect 263604 -6102 263786 -5866
rect 264022 -6102 264204 -5866
rect 263604 -6186 264204 -6102
rect 263604 -6422 263786 -6186
rect 264022 -6422 264204 -6186
rect 263604 -7364 264204 -6422
rect 281604 -6786 282204 30698
rect 288804 542454 289404 577898
rect 288804 542218 288986 542454
rect 289222 542218 289404 542454
rect 288804 542134 289404 542218
rect 288804 541898 288986 542134
rect 289222 541898 289404 542134
rect 288804 506454 289404 541898
rect 288804 506218 288986 506454
rect 289222 506218 289404 506454
rect 288804 506134 289404 506218
rect 288804 505898 288986 506134
rect 289222 505898 289404 506134
rect 288804 470454 289404 505898
rect 288804 470218 288986 470454
rect 289222 470218 289404 470454
rect 288804 470134 289404 470218
rect 288804 469898 288986 470134
rect 289222 469898 289404 470134
rect 288804 434454 289404 469898
rect 288804 434218 288986 434454
rect 289222 434218 289404 434454
rect 288804 434134 289404 434218
rect 288804 433898 288986 434134
rect 289222 433898 289404 434134
rect 288804 398454 289404 433898
rect 288804 398218 288986 398454
rect 289222 398218 289404 398454
rect 288804 398134 289404 398218
rect 288804 397898 288986 398134
rect 289222 397898 289404 398134
rect 288804 362454 289404 397898
rect 288804 362218 288986 362454
rect 289222 362218 289404 362454
rect 288804 362134 289404 362218
rect 288804 361898 288986 362134
rect 289222 361898 289404 362134
rect 288804 326454 289404 361898
rect 288804 326218 288986 326454
rect 289222 326218 289404 326454
rect 288804 326134 289404 326218
rect 288804 325898 288986 326134
rect 289222 325898 289404 326134
rect 288804 290454 289404 325898
rect 288804 290218 288986 290454
rect 289222 290218 289404 290454
rect 288804 290134 289404 290218
rect 288804 289898 288986 290134
rect 289222 289898 289404 290134
rect 288804 254454 289404 289898
rect 288804 254218 288986 254454
rect 289222 254218 289404 254454
rect 288804 254134 289404 254218
rect 288804 253898 288986 254134
rect 289222 253898 289404 254134
rect 288804 218454 289404 253898
rect 288804 218218 288986 218454
rect 289222 218218 289404 218454
rect 288804 218134 289404 218218
rect 288804 217898 288986 218134
rect 289222 217898 289404 218134
rect 288804 182454 289404 217898
rect 288804 182218 288986 182454
rect 289222 182218 289404 182454
rect 288804 182134 289404 182218
rect 288804 181898 288986 182134
rect 289222 181898 289404 182134
rect 288804 146454 289404 181898
rect 288804 146218 288986 146454
rect 289222 146218 289404 146454
rect 288804 146134 289404 146218
rect 288804 145898 288986 146134
rect 289222 145898 289404 146134
rect 288804 110454 289404 145898
rect 288804 110218 288986 110454
rect 289222 110218 289404 110454
rect 288804 110134 289404 110218
rect 288804 109898 288986 110134
rect 289222 109898 289404 110134
rect 288804 74454 289404 109898
rect 288804 74218 288986 74454
rect 289222 74218 289404 74454
rect 288804 74134 289404 74218
rect 288804 73898 288986 74134
rect 289222 73898 289404 74134
rect 288804 38454 289404 73898
rect 288804 38218 288986 38454
rect 289222 38218 289404 38454
rect 288804 38134 289404 38218
rect 288804 37898 288986 38134
rect 289222 37898 289404 38134
rect 288804 2454 289404 37898
rect 288804 2218 288986 2454
rect 289222 2218 289404 2454
rect 288804 2134 289404 2218
rect 288804 1898 288986 2134
rect 289222 1898 289404 2134
rect 288804 -346 289404 1898
rect 288804 -582 288986 -346
rect 289222 -582 289404 -346
rect 288804 -666 289404 -582
rect 288804 -902 288986 -666
rect 289222 -902 289404 -666
rect 288804 -1844 289404 -902
rect 292404 690054 293004 706122
rect 292404 689818 292586 690054
rect 292822 689818 293004 690054
rect 292404 689734 293004 689818
rect 292404 689498 292586 689734
rect 292822 689498 293004 689734
rect 292404 654054 293004 689498
rect 292404 653818 292586 654054
rect 292822 653818 293004 654054
rect 292404 653734 293004 653818
rect 292404 653498 292586 653734
rect 292822 653498 293004 653734
rect 292404 618054 293004 653498
rect 292404 617818 292586 618054
rect 292822 617818 293004 618054
rect 292404 617734 293004 617818
rect 292404 617498 292586 617734
rect 292822 617498 293004 617734
rect 292404 582054 293004 617498
rect 292404 581818 292586 582054
rect 292822 581818 293004 582054
rect 292404 581734 293004 581818
rect 292404 581498 292586 581734
rect 292822 581498 293004 581734
rect 292404 546054 293004 581498
rect 296004 693654 296604 707962
rect 296004 693418 296186 693654
rect 296422 693418 296604 693654
rect 296004 693334 296604 693418
rect 296004 693098 296186 693334
rect 296422 693098 296604 693334
rect 296004 657654 296604 693098
rect 296004 657418 296186 657654
rect 296422 657418 296604 657654
rect 296004 657334 296604 657418
rect 296004 657098 296186 657334
rect 296422 657098 296604 657334
rect 296004 621654 296604 657098
rect 296004 621418 296186 621654
rect 296422 621418 296604 621654
rect 296004 621334 296604 621418
rect 296004 621098 296186 621334
rect 296422 621098 296604 621334
rect 296004 585654 296604 621098
rect 296004 585418 296186 585654
rect 296422 585418 296604 585654
rect 296004 585334 296604 585418
rect 296004 585098 296186 585334
rect 296422 585098 296604 585334
rect 293174 561645 293234 562582
rect 293171 561644 293237 561645
rect 293171 561580 293172 561644
rect 293236 561580 293237 561644
rect 293171 561579 293237 561580
rect 292404 545818 292586 546054
rect 292822 545818 293004 546054
rect 292404 545734 293004 545818
rect 292404 545498 292586 545734
rect 292822 545498 293004 545734
rect 292404 510054 293004 545498
rect 292404 509818 292586 510054
rect 292822 509818 293004 510054
rect 292404 509734 293004 509818
rect 292404 509498 292586 509734
rect 292822 509498 293004 509734
rect 292404 474054 293004 509498
rect 292404 473818 292586 474054
rect 292822 473818 293004 474054
rect 292404 473734 293004 473818
rect 292404 473498 292586 473734
rect 292822 473498 293004 473734
rect 292404 438054 293004 473498
rect 292404 437818 292586 438054
rect 292822 437818 293004 438054
rect 292404 437734 293004 437818
rect 292404 437498 292586 437734
rect 292822 437498 293004 437734
rect 292404 402054 293004 437498
rect 292404 401818 292586 402054
rect 292822 401818 293004 402054
rect 292404 401734 293004 401818
rect 292404 401498 292586 401734
rect 292822 401498 293004 401734
rect 292404 366054 293004 401498
rect 292404 365818 292586 366054
rect 292822 365818 293004 366054
rect 292404 365734 293004 365818
rect 292404 365498 292586 365734
rect 292822 365498 293004 365734
rect 292404 330054 293004 365498
rect 292404 329818 292586 330054
rect 292822 329818 293004 330054
rect 292404 329734 293004 329818
rect 292404 329498 292586 329734
rect 292822 329498 293004 329734
rect 292404 294054 293004 329498
rect 292404 293818 292586 294054
rect 292822 293818 293004 294054
rect 292404 293734 293004 293818
rect 292404 293498 292586 293734
rect 292822 293498 293004 293734
rect 292404 258054 293004 293498
rect 292404 257818 292586 258054
rect 292822 257818 293004 258054
rect 292404 257734 293004 257818
rect 292404 257498 292586 257734
rect 292822 257498 293004 257734
rect 292404 222054 293004 257498
rect 292404 221818 292586 222054
rect 292822 221818 293004 222054
rect 292404 221734 293004 221818
rect 292404 221498 292586 221734
rect 292822 221498 293004 221734
rect 292404 186054 293004 221498
rect 292404 185818 292586 186054
rect 292822 185818 293004 186054
rect 292404 185734 293004 185818
rect 292404 185498 292586 185734
rect 292822 185498 293004 185734
rect 292404 150054 293004 185498
rect 292404 149818 292586 150054
rect 292822 149818 293004 150054
rect 292404 149734 293004 149818
rect 292404 149498 292586 149734
rect 292822 149498 293004 149734
rect 292404 114054 293004 149498
rect 292404 113818 292586 114054
rect 292822 113818 293004 114054
rect 292404 113734 293004 113818
rect 292404 113498 292586 113734
rect 292822 113498 293004 113734
rect 292404 78054 293004 113498
rect 292404 77818 292586 78054
rect 292822 77818 293004 78054
rect 292404 77734 293004 77818
rect 292404 77498 292586 77734
rect 292822 77498 293004 77734
rect 292404 42054 293004 77498
rect 292404 41818 292586 42054
rect 292822 41818 293004 42054
rect 292404 41734 293004 41818
rect 292404 41498 292586 41734
rect 292822 41498 293004 41734
rect 292404 6054 293004 41498
rect 292404 5818 292586 6054
rect 292822 5818 293004 6054
rect 292404 5734 293004 5818
rect 292404 5498 292586 5734
rect 292822 5498 293004 5734
rect 292404 -2186 293004 5498
rect 292404 -2422 292586 -2186
rect 292822 -2422 293004 -2186
rect 292404 -2506 293004 -2422
rect 292404 -2742 292586 -2506
rect 292822 -2742 293004 -2506
rect 292404 -3684 293004 -2742
rect 296004 549654 296604 585098
rect 299604 697254 300204 709802
rect 317604 711278 318204 711300
rect 317604 711042 317786 711278
rect 318022 711042 318204 711278
rect 317604 710958 318204 711042
rect 317604 710722 317786 710958
rect 318022 710722 318204 710958
rect 314004 709438 314604 709460
rect 314004 709202 314186 709438
rect 314422 709202 314604 709438
rect 314004 709118 314604 709202
rect 314004 708882 314186 709118
rect 314422 708882 314604 709118
rect 310404 707598 311004 707620
rect 310404 707362 310586 707598
rect 310822 707362 311004 707598
rect 310404 707278 311004 707362
rect 310404 707042 310586 707278
rect 310822 707042 311004 707278
rect 299604 697018 299786 697254
rect 300022 697018 300204 697254
rect 299604 696934 300204 697018
rect 299604 696698 299786 696934
rect 300022 696698 300204 696934
rect 299604 661254 300204 696698
rect 299604 661018 299786 661254
rect 300022 661018 300204 661254
rect 299604 660934 300204 661018
rect 299604 660698 299786 660934
rect 300022 660698 300204 660934
rect 299604 625254 300204 660698
rect 299604 625018 299786 625254
rect 300022 625018 300204 625254
rect 299604 624934 300204 625018
rect 299604 624698 299786 624934
rect 300022 624698 300204 624934
rect 299604 589254 300204 624698
rect 299604 589018 299786 589254
rect 300022 589018 300204 589254
rect 299604 588934 300204 589018
rect 299604 588698 299786 588934
rect 300022 588698 300204 588934
rect 299427 559876 299493 559877
rect 299427 559812 299428 559876
rect 299492 559812 299493 559876
rect 299427 559811 299493 559812
rect 299430 559605 299490 559811
rect 299427 559604 299493 559605
rect 299427 559540 299428 559604
rect 299492 559540 299493 559604
rect 299427 559539 299493 559540
rect 299427 559332 299493 559333
rect 299427 559268 299428 559332
rect 299492 559268 299493 559332
rect 299427 559267 299493 559268
rect 299430 559061 299490 559267
rect 299427 559060 299493 559061
rect 299427 558996 299428 559060
rect 299492 558996 299493 559060
rect 299427 558995 299493 558996
rect 296004 549418 296186 549654
rect 296422 549418 296604 549654
rect 296004 549334 296604 549418
rect 296004 549098 296186 549334
rect 296422 549098 296604 549334
rect 296004 513654 296604 549098
rect 296004 513418 296186 513654
rect 296422 513418 296604 513654
rect 296004 513334 296604 513418
rect 296004 513098 296186 513334
rect 296422 513098 296604 513334
rect 296004 477654 296604 513098
rect 296004 477418 296186 477654
rect 296422 477418 296604 477654
rect 296004 477334 296604 477418
rect 296004 477098 296186 477334
rect 296422 477098 296604 477334
rect 296004 441654 296604 477098
rect 296004 441418 296186 441654
rect 296422 441418 296604 441654
rect 296004 441334 296604 441418
rect 296004 441098 296186 441334
rect 296422 441098 296604 441334
rect 296004 405654 296604 441098
rect 296004 405418 296186 405654
rect 296422 405418 296604 405654
rect 296004 405334 296604 405418
rect 296004 405098 296186 405334
rect 296422 405098 296604 405334
rect 296004 369654 296604 405098
rect 296004 369418 296186 369654
rect 296422 369418 296604 369654
rect 296004 369334 296604 369418
rect 296004 369098 296186 369334
rect 296422 369098 296604 369334
rect 296004 333654 296604 369098
rect 296004 333418 296186 333654
rect 296422 333418 296604 333654
rect 296004 333334 296604 333418
rect 296004 333098 296186 333334
rect 296422 333098 296604 333334
rect 296004 297654 296604 333098
rect 296004 297418 296186 297654
rect 296422 297418 296604 297654
rect 296004 297334 296604 297418
rect 296004 297098 296186 297334
rect 296422 297098 296604 297334
rect 296004 261654 296604 297098
rect 296004 261418 296186 261654
rect 296422 261418 296604 261654
rect 296004 261334 296604 261418
rect 296004 261098 296186 261334
rect 296422 261098 296604 261334
rect 296004 225654 296604 261098
rect 296004 225418 296186 225654
rect 296422 225418 296604 225654
rect 296004 225334 296604 225418
rect 296004 225098 296186 225334
rect 296422 225098 296604 225334
rect 296004 189654 296604 225098
rect 296004 189418 296186 189654
rect 296422 189418 296604 189654
rect 296004 189334 296604 189418
rect 296004 189098 296186 189334
rect 296422 189098 296604 189334
rect 296004 153654 296604 189098
rect 299604 553254 300204 588698
rect 299604 553018 299786 553254
rect 300022 553018 300204 553254
rect 299604 552934 300204 553018
rect 299604 552698 299786 552934
rect 300022 552698 300204 552934
rect 299604 517254 300204 552698
rect 299604 517018 299786 517254
rect 300022 517018 300204 517254
rect 299604 516934 300204 517018
rect 299604 516698 299786 516934
rect 300022 516698 300204 516934
rect 299604 481254 300204 516698
rect 299604 481018 299786 481254
rect 300022 481018 300204 481254
rect 299604 480934 300204 481018
rect 299604 480698 299786 480934
rect 300022 480698 300204 480934
rect 299604 445254 300204 480698
rect 299604 445018 299786 445254
rect 300022 445018 300204 445254
rect 299604 444934 300204 445018
rect 299604 444698 299786 444934
rect 300022 444698 300204 444934
rect 299604 409254 300204 444698
rect 299604 409018 299786 409254
rect 300022 409018 300204 409254
rect 299604 408934 300204 409018
rect 299604 408698 299786 408934
rect 300022 408698 300204 408934
rect 299604 373254 300204 408698
rect 299604 373018 299786 373254
rect 300022 373018 300204 373254
rect 299604 372934 300204 373018
rect 299604 372698 299786 372934
rect 300022 372698 300204 372934
rect 299604 337254 300204 372698
rect 299604 337018 299786 337254
rect 300022 337018 300204 337254
rect 299604 336934 300204 337018
rect 299604 336698 299786 336934
rect 300022 336698 300204 336934
rect 299604 301254 300204 336698
rect 299604 301018 299786 301254
rect 300022 301018 300204 301254
rect 299604 300934 300204 301018
rect 299604 300698 299786 300934
rect 300022 300698 300204 300934
rect 299604 265254 300204 300698
rect 299604 265018 299786 265254
rect 300022 265018 300204 265254
rect 299604 264934 300204 265018
rect 299604 264698 299786 264934
rect 300022 264698 300204 264934
rect 299604 229254 300204 264698
rect 299604 229018 299786 229254
rect 300022 229018 300204 229254
rect 299604 228934 300204 229018
rect 299604 228698 299786 228934
rect 300022 228698 300204 228934
rect 299604 193254 300204 228698
rect 299604 193018 299786 193254
rect 300022 193018 300204 193254
rect 299604 192934 300204 193018
rect 299604 192698 299786 192934
rect 300022 192698 300204 192934
rect 299243 181252 299309 181253
rect 299243 181188 299244 181252
rect 299308 181250 299309 181252
rect 299308 181190 299490 181250
rect 299308 181188 299309 181190
rect 299243 181187 299309 181188
rect 299430 181117 299490 181190
rect 299427 181116 299493 181117
rect 299427 181052 299428 181116
rect 299492 181052 299493 181116
rect 299427 181051 299493 181052
rect 296004 153418 296186 153654
rect 296422 153418 296604 153654
rect 296004 153334 296604 153418
rect 296004 153098 296186 153334
rect 296422 153098 296604 153334
rect 296004 117654 296604 153098
rect 296004 117418 296186 117654
rect 296422 117418 296604 117654
rect 296004 117334 296604 117418
rect 296004 117098 296186 117334
rect 296422 117098 296604 117334
rect 296004 81654 296604 117098
rect 299604 157254 300204 192698
rect 299604 157018 299786 157254
rect 300022 157018 300204 157254
rect 299604 156934 300204 157018
rect 299604 156698 299786 156934
rect 300022 156698 300204 156934
rect 299604 121254 300204 156698
rect 299604 121018 299786 121254
rect 300022 121018 300204 121254
rect 299604 120934 300204 121018
rect 299604 120698 299786 120934
rect 300022 120698 300204 120934
rect 299427 87548 299493 87549
rect 299427 87484 299428 87548
rect 299492 87484 299493 87548
rect 299427 87483 299493 87484
rect 299430 87277 299490 87483
rect 299427 87276 299493 87277
rect 299427 87212 299428 87276
rect 299492 87212 299493 87276
rect 299427 87211 299493 87212
rect 296004 81418 296186 81654
rect 296422 81418 296604 81654
rect 296004 81334 296604 81418
rect 296004 81098 296186 81334
rect 296422 81098 296604 81334
rect 296004 45654 296604 81098
rect 296004 45418 296186 45654
rect 296422 45418 296604 45654
rect 296004 45334 296604 45418
rect 296004 45098 296186 45334
rect 296422 45098 296604 45334
rect 296004 9654 296604 45098
rect 296004 9418 296186 9654
rect 296422 9418 296604 9654
rect 296004 9334 296604 9418
rect 296004 9098 296186 9334
rect 296422 9098 296604 9334
rect 296004 -4026 296604 9098
rect 296004 -4262 296186 -4026
rect 296422 -4262 296604 -4026
rect 296004 -4346 296604 -4262
rect 296004 -4582 296186 -4346
rect 296422 -4582 296604 -4346
rect 296004 -5524 296604 -4582
rect 299604 85254 300204 120698
rect 299604 85018 299786 85254
rect 300022 85018 300204 85254
rect 299604 84934 300204 85018
rect 299604 84698 299786 84934
rect 300022 84698 300204 84934
rect 299604 49254 300204 84698
rect 299604 49018 299786 49254
rect 300022 49018 300204 49254
rect 299604 48934 300204 49018
rect 299604 48698 299786 48934
rect 300022 48698 300204 48934
rect 299604 13254 300204 48698
rect 299604 13018 299786 13254
rect 300022 13018 300204 13254
rect 299604 12934 300204 13018
rect 299604 12698 299786 12934
rect 300022 12698 300204 12934
rect 281604 -7022 281786 -6786
rect 282022 -7022 282204 -6786
rect 281604 -7106 282204 -7022
rect 281604 -7342 281786 -7106
rect 282022 -7342 282204 -7106
rect 281604 -7364 282204 -7342
rect 299604 -5866 300204 12698
rect 306804 705758 307404 705780
rect 306804 705522 306986 705758
rect 307222 705522 307404 705758
rect 306804 705438 307404 705522
rect 306804 705202 306986 705438
rect 307222 705202 307404 705438
rect 306804 668454 307404 705202
rect 306804 668218 306986 668454
rect 307222 668218 307404 668454
rect 306804 668134 307404 668218
rect 306804 667898 306986 668134
rect 307222 667898 307404 668134
rect 306804 632454 307404 667898
rect 306804 632218 306986 632454
rect 307222 632218 307404 632454
rect 306804 632134 307404 632218
rect 306804 631898 306986 632134
rect 307222 631898 307404 632134
rect 306804 596454 307404 631898
rect 306804 596218 306986 596454
rect 307222 596218 307404 596454
rect 306804 596134 307404 596218
rect 306804 595898 306986 596134
rect 307222 595898 307404 596134
rect 306804 560454 307404 595898
rect 310404 672054 311004 707042
rect 310404 671818 310586 672054
rect 310822 671818 311004 672054
rect 310404 671734 311004 671818
rect 310404 671498 310586 671734
rect 310822 671498 311004 671734
rect 310404 636054 311004 671498
rect 310404 635818 310586 636054
rect 310822 635818 311004 636054
rect 310404 635734 311004 635818
rect 310404 635498 310586 635734
rect 310822 635498 311004 635734
rect 310404 600054 311004 635498
rect 310404 599818 310586 600054
rect 310822 599818 311004 600054
rect 310404 599734 311004 599818
rect 310404 599498 310586 599734
rect 310822 599498 311004 599734
rect 310404 564054 311004 599498
rect 310404 563818 310586 564054
rect 310822 563818 311004 564054
rect 310404 563734 311004 563818
rect 310404 563498 310586 563734
rect 310822 563498 311004 563734
rect 308995 560556 309061 560557
rect 308995 560492 308996 560556
rect 309060 560492 309061 560556
rect 308995 560491 309061 560492
rect 306804 560218 306986 560454
rect 307222 560218 307404 560454
rect 308998 560421 309058 560491
rect 308995 560420 309061 560421
rect 308995 560356 308996 560420
rect 309060 560356 309061 560420
rect 308995 560355 309061 560356
rect 306804 560134 307404 560218
rect 306804 559898 306986 560134
rect 307222 559898 307404 560134
rect 306804 524454 307404 559898
rect 307707 559468 307773 559469
rect 307707 559404 307708 559468
rect 307772 559404 307773 559468
rect 307707 559403 307773 559404
rect 307710 559330 307770 559403
rect 307891 559332 307957 559333
rect 307891 559330 307892 559332
rect 307710 559270 307892 559330
rect 307891 559268 307892 559270
rect 307956 559268 307957 559332
rect 307891 559267 307957 559268
rect 306804 524218 306986 524454
rect 307222 524218 307404 524454
rect 306804 524134 307404 524218
rect 306804 523898 306986 524134
rect 307222 523898 307404 524134
rect 306804 488454 307404 523898
rect 306804 488218 306986 488454
rect 307222 488218 307404 488454
rect 306804 488134 307404 488218
rect 306804 487898 306986 488134
rect 307222 487898 307404 488134
rect 306804 452454 307404 487898
rect 306804 452218 306986 452454
rect 307222 452218 307404 452454
rect 306804 452134 307404 452218
rect 306804 451898 306986 452134
rect 307222 451898 307404 452134
rect 306804 416454 307404 451898
rect 306804 416218 306986 416454
rect 307222 416218 307404 416454
rect 306804 416134 307404 416218
rect 306804 415898 306986 416134
rect 307222 415898 307404 416134
rect 306804 380454 307404 415898
rect 306804 380218 306986 380454
rect 307222 380218 307404 380454
rect 306804 380134 307404 380218
rect 306804 379898 306986 380134
rect 307222 379898 307404 380134
rect 306804 344454 307404 379898
rect 306804 344218 306986 344454
rect 307222 344218 307404 344454
rect 306804 344134 307404 344218
rect 306804 343898 306986 344134
rect 307222 343898 307404 344134
rect 306804 308454 307404 343898
rect 306804 308218 306986 308454
rect 307222 308218 307404 308454
rect 306804 308134 307404 308218
rect 306804 307898 306986 308134
rect 307222 307898 307404 308134
rect 306804 272454 307404 307898
rect 306804 272218 306986 272454
rect 307222 272218 307404 272454
rect 306804 272134 307404 272218
rect 306804 271898 306986 272134
rect 307222 271898 307404 272134
rect 306804 236454 307404 271898
rect 306804 236218 306986 236454
rect 307222 236218 307404 236454
rect 306804 236134 307404 236218
rect 306804 235898 306986 236134
rect 307222 235898 307404 236134
rect 306804 200454 307404 235898
rect 306804 200218 306986 200454
rect 307222 200218 307404 200454
rect 306804 200134 307404 200218
rect 306804 199898 306986 200134
rect 307222 199898 307404 200134
rect 306804 164454 307404 199898
rect 306804 164218 306986 164454
rect 307222 164218 307404 164454
rect 306804 164134 307404 164218
rect 306804 163898 306986 164134
rect 307222 163898 307404 164134
rect 306804 128454 307404 163898
rect 306804 128218 306986 128454
rect 307222 128218 307404 128454
rect 306804 128134 307404 128218
rect 306804 127898 306986 128134
rect 307222 127898 307404 128134
rect 306804 92454 307404 127898
rect 306804 92218 306986 92454
rect 307222 92218 307404 92454
rect 306804 92134 307404 92218
rect 306804 91898 306986 92134
rect 307222 91898 307404 92134
rect 306804 56454 307404 91898
rect 306804 56218 306986 56454
rect 307222 56218 307404 56454
rect 306804 56134 307404 56218
rect 306804 55898 306986 56134
rect 307222 55898 307404 56134
rect 306804 20454 307404 55898
rect 306804 20218 306986 20454
rect 307222 20218 307404 20454
rect 306804 20134 307404 20218
rect 306804 19898 306986 20134
rect 307222 19898 307404 20134
rect 306804 -1266 307404 19898
rect 306804 -1502 306986 -1266
rect 307222 -1502 307404 -1266
rect 306804 -1586 307404 -1502
rect 306804 -1822 306986 -1586
rect 307222 -1822 307404 -1586
rect 306804 -1844 307404 -1822
rect 310404 528054 311004 563498
rect 314004 675654 314604 708882
rect 314004 675418 314186 675654
rect 314422 675418 314604 675654
rect 314004 675334 314604 675418
rect 314004 675098 314186 675334
rect 314422 675098 314604 675334
rect 314004 639654 314604 675098
rect 314004 639418 314186 639654
rect 314422 639418 314604 639654
rect 314004 639334 314604 639418
rect 314004 639098 314186 639334
rect 314422 639098 314604 639334
rect 314004 603654 314604 639098
rect 314004 603418 314186 603654
rect 314422 603418 314604 603654
rect 314004 603334 314604 603418
rect 314004 603098 314186 603334
rect 314422 603098 314604 603334
rect 314004 567654 314604 603098
rect 314004 567418 314186 567654
rect 314422 567418 314604 567654
rect 314004 567334 314604 567418
rect 314004 567098 314186 567334
rect 314422 567098 314604 567334
rect 311758 559270 312002 559330
rect 311758 559061 311818 559270
rect 311942 559197 312002 559270
rect 311939 559196 312005 559197
rect 311939 559132 311940 559196
rect 312004 559132 312005 559196
rect 311939 559131 312005 559132
rect 311755 559060 311821 559061
rect 311755 558996 311756 559060
rect 311820 558996 311821 559060
rect 311755 558995 311821 558996
rect 310404 527818 310586 528054
rect 310822 527818 311004 528054
rect 310404 527734 311004 527818
rect 310404 527498 310586 527734
rect 310822 527498 311004 527734
rect 310404 492054 311004 527498
rect 310404 491818 310586 492054
rect 310822 491818 311004 492054
rect 310404 491734 311004 491818
rect 310404 491498 310586 491734
rect 310822 491498 311004 491734
rect 310404 456054 311004 491498
rect 310404 455818 310586 456054
rect 310822 455818 311004 456054
rect 310404 455734 311004 455818
rect 310404 455498 310586 455734
rect 310822 455498 311004 455734
rect 310404 420054 311004 455498
rect 310404 419818 310586 420054
rect 310822 419818 311004 420054
rect 310404 419734 311004 419818
rect 310404 419498 310586 419734
rect 310822 419498 311004 419734
rect 310404 384054 311004 419498
rect 310404 383818 310586 384054
rect 310822 383818 311004 384054
rect 310404 383734 311004 383818
rect 310404 383498 310586 383734
rect 310822 383498 311004 383734
rect 310404 348054 311004 383498
rect 310404 347818 310586 348054
rect 310822 347818 311004 348054
rect 310404 347734 311004 347818
rect 310404 347498 310586 347734
rect 310822 347498 311004 347734
rect 310404 312054 311004 347498
rect 310404 311818 310586 312054
rect 310822 311818 311004 312054
rect 310404 311734 311004 311818
rect 310404 311498 310586 311734
rect 310822 311498 311004 311734
rect 310404 276054 311004 311498
rect 310404 275818 310586 276054
rect 310822 275818 311004 276054
rect 310404 275734 311004 275818
rect 310404 275498 310586 275734
rect 310822 275498 311004 275734
rect 310404 240054 311004 275498
rect 310404 239818 310586 240054
rect 310822 239818 311004 240054
rect 310404 239734 311004 239818
rect 310404 239498 310586 239734
rect 310822 239498 311004 239734
rect 310404 204054 311004 239498
rect 310404 203818 310586 204054
rect 310822 203818 311004 204054
rect 310404 203734 311004 203818
rect 310404 203498 310586 203734
rect 310822 203498 311004 203734
rect 310404 168054 311004 203498
rect 310404 167818 310586 168054
rect 310822 167818 311004 168054
rect 310404 167734 311004 167818
rect 310404 167498 310586 167734
rect 310822 167498 311004 167734
rect 310404 132054 311004 167498
rect 310404 131818 310586 132054
rect 310822 131818 311004 132054
rect 310404 131734 311004 131818
rect 310404 131498 310586 131734
rect 310822 131498 311004 131734
rect 310404 96054 311004 131498
rect 310404 95818 310586 96054
rect 310822 95818 311004 96054
rect 310404 95734 311004 95818
rect 310404 95498 310586 95734
rect 310822 95498 311004 95734
rect 310404 60054 311004 95498
rect 310404 59818 310586 60054
rect 310822 59818 311004 60054
rect 310404 59734 311004 59818
rect 310404 59498 310586 59734
rect 310822 59498 311004 59734
rect 310404 24054 311004 59498
rect 310404 23818 310586 24054
rect 310822 23818 311004 24054
rect 310404 23734 311004 23818
rect 310404 23498 310586 23734
rect 310822 23498 311004 23734
rect 310404 -3106 311004 23498
rect 310404 -3342 310586 -3106
rect 310822 -3342 311004 -3106
rect 310404 -3426 311004 -3342
rect 310404 -3662 310586 -3426
rect 310822 -3662 311004 -3426
rect 310404 -3684 311004 -3662
rect 314004 531654 314604 567098
rect 314004 531418 314186 531654
rect 314422 531418 314604 531654
rect 314004 531334 314604 531418
rect 314004 531098 314186 531334
rect 314422 531098 314604 531334
rect 314004 495654 314604 531098
rect 314004 495418 314186 495654
rect 314422 495418 314604 495654
rect 314004 495334 314604 495418
rect 314004 495098 314186 495334
rect 314422 495098 314604 495334
rect 314004 459654 314604 495098
rect 314004 459418 314186 459654
rect 314422 459418 314604 459654
rect 314004 459334 314604 459418
rect 314004 459098 314186 459334
rect 314422 459098 314604 459334
rect 314004 423654 314604 459098
rect 314004 423418 314186 423654
rect 314422 423418 314604 423654
rect 314004 423334 314604 423418
rect 314004 423098 314186 423334
rect 314422 423098 314604 423334
rect 314004 387654 314604 423098
rect 314004 387418 314186 387654
rect 314422 387418 314604 387654
rect 314004 387334 314604 387418
rect 314004 387098 314186 387334
rect 314422 387098 314604 387334
rect 314004 351654 314604 387098
rect 314004 351418 314186 351654
rect 314422 351418 314604 351654
rect 314004 351334 314604 351418
rect 314004 351098 314186 351334
rect 314422 351098 314604 351334
rect 314004 315654 314604 351098
rect 314004 315418 314186 315654
rect 314422 315418 314604 315654
rect 314004 315334 314604 315418
rect 314004 315098 314186 315334
rect 314422 315098 314604 315334
rect 314004 279654 314604 315098
rect 314004 279418 314186 279654
rect 314422 279418 314604 279654
rect 314004 279334 314604 279418
rect 314004 279098 314186 279334
rect 314422 279098 314604 279334
rect 314004 243654 314604 279098
rect 314004 243418 314186 243654
rect 314422 243418 314604 243654
rect 314004 243334 314604 243418
rect 314004 243098 314186 243334
rect 314422 243098 314604 243334
rect 314004 207654 314604 243098
rect 314004 207418 314186 207654
rect 314422 207418 314604 207654
rect 314004 207334 314604 207418
rect 314004 207098 314186 207334
rect 314422 207098 314604 207334
rect 314004 171654 314604 207098
rect 314004 171418 314186 171654
rect 314422 171418 314604 171654
rect 314004 171334 314604 171418
rect 314004 171098 314186 171334
rect 314422 171098 314604 171334
rect 314004 135654 314604 171098
rect 314004 135418 314186 135654
rect 314422 135418 314604 135654
rect 314004 135334 314604 135418
rect 314004 135098 314186 135334
rect 314422 135098 314604 135334
rect 314004 99654 314604 135098
rect 314004 99418 314186 99654
rect 314422 99418 314604 99654
rect 314004 99334 314604 99418
rect 314004 99098 314186 99334
rect 314422 99098 314604 99334
rect 314004 63654 314604 99098
rect 317604 679254 318204 710722
rect 335604 710358 336204 711300
rect 335604 710122 335786 710358
rect 336022 710122 336204 710358
rect 335604 710038 336204 710122
rect 335604 709802 335786 710038
rect 336022 709802 336204 710038
rect 332004 708518 332604 709460
rect 332004 708282 332186 708518
rect 332422 708282 332604 708518
rect 332004 708198 332604 708282
rect 332004 707962 332186 708198
rect 332422 707962 332604 708198
rect 328404 706678 329004 707620
rect 328404 706442 328586 706678
rect 328822 706442 329004 706678
rect 328404 706358 329004 706442
rect 328404 706122 328586 706358
rect 328822 706122 329004 706358
rect 317604 679018 317786 679254
rect 318022 679018 318204 679254
rect 317604 678934 318204 679018
rect 317604 678698 317786 678934
rect 318022 678698 318204 678934
rect 317604 643254 318204 678698
rect 317604 643018 317786 643254
rect 318022 643018 318204 643254
rect 317604 642934 318204 643018
rect 317604 642698 317786 642934
rect 318022 642698 318204 642934
rect 317604 607254 318204 642698
rect 317604 607018 317786 607254
rect 318022 607018 318204 607254
rect 317604 606934 318204 607018
rect 317604 606698 317786 606934
rect 318022 606698 318204 606934
rect 317604 571254 318204 606698
rect 317604 571018 317786 571254
rect 318022 571018 318204 571254
rect 317604 570934 318204 571018
rect 317604 570698 317786 570934
rect 318022 570698 318204 570934
rect 317604 535254 318204 570698
rect 324804 704838 325404 705780
rect 324804 704602 324986 704838
rect 325222 704602 325404 704838
rect 324804 704518 325404 704602
rect 324804 704282 324986 704518
rect 325222 704282 325404 704518
rect 324804 686454 325404 704282
rect 324804 686218 324986 686454
rect 325222 686218 325404 686454
rect 324804 686134 325404 686218
rect 324804 685898 324986 686134
rect 325222 685898 325404 686134
rect 324804 650454 325404 685898
rect 324804 650218 324986 650454
rect 325222 650218 325404 650454
rect 324804 650134 325404 650218
rect 324804 649898 324986 650134
rect 325222 649898 325404 650134
rect 324804 614454 325404 649898
rect 324804 614218 324986 614454
rect 325222 614218 325404 614454
rect 324804 614134 325404 614218
rect 324804 613898 324986 614134
rect 325222 613898 325404 614134
rect 324804 578454 325404 613898
rect 324804 578218 324986 578454
rect 325222 578218 325404 578454
rect 324804 578134 325404 578218
rect 324804 577898 324986 578134
rect 325222 577898 325404 578134
rect 318714 561310 319214 561370
rect 318747 559060 318813 559061
rect 318747 558996 318748 559060
rect 318812 558996 318813 559060
rect 318747 558995 318813 558996
rect 318750 558789 318810 558995
rect 318747 558788 318813 558789
rect 318747 558724 318748 558788
rect 318812 558724 318813 558788
rect 318747 558723 318813 558724
rect 317604 535018 317786 535254
rect 318022 535018 318204 535254
rect 317604 534934 318204 535018
rect 317604 534698 317786 534934
rect 318022 534698 318204 534934
rect 317604 499254 318204 534698
rect 317604 499018 317786 499254
rect 318022 499018 318204 499254
rect 317604 498934 318204 499018
rect 317604 498698 317786 498934
rect 318022 498698 318204 498934
rect 317604 463254 318204 498698
rect 317604 463018 317786 463254
rect 318022 463018 318204 463254
rect 317604 462934 318204 463018
rect 317604 462698 317786 462934
rect 318022 462698 318204 462934
rect 317604 427254 318204 462698
rect 317604 427018 317786 427254
rect 318022 427018 318204 427254
rect 317604 426934 318204 427018
rect 317604 426698 317786 426934
rect 318022 426698 318204 426934
rect 317604 391254 318204 426698
rect 317604 391018 317786 391254
rect 318022 391018 318204 391254
rect 317604 390934 318204 391018
rect 317604 390698 317786 390934
rect 318022 390698 318204 390934
rect 317604 355254 318204 390698
rect 317604 355018 317786 355254
rect 318022 355018 318204 355254
rect 317604 354934 318204 355018
rect 317604 354698 317786 354934
rect 318022 354698 318204 354934
rect 317604 319254 318204 354698
rect 317604 319018 317786 319254
rect 318022 319018 318204 319254
rect 317604 318934 318204 319018
rect 317604 318698 317786 318934
rect 318022 318698 318204 318934
rect 317604 283254 318204 318698
rect 317604 283018 317786 283254
rect 318022 283018 318204 283254
rect 317604 282934 318204 283018
rect 317604 282698 317786 282934
rect 318022 282698 318204 282934
rect 317604 247254 318204 282698
rect 317604 247018 317786 247254
rect 318022 247018 318204 247254
rect 317604 246934 318204 247018
rect 317604 246698 317786 246934
rect 318022 246698 318204 246934
rect 317604 211254 318204 246698
rect 317604 211018 317786 211254
rect 318022 211018 318204 211254
rect 317604 210934 318204 211018
rect 317604 210698 317786 210934
rect 318022 210698 318204 210934
rect 317604 175254 318204 210698
rect 317604 175018 317786 175254
rect 318022 175018 318204 175254
rect 317604 174934 318204 175018
rect 317604 174698 317786 174934
rect 318022 174698 318204 174934
rect 317604 139254 318204 174698
rect 317604 139018 317786 139254
rect 318022 139018 318204 139254
rect 317604 138934 318204 139018
rect 317604 138698 317786 138934
rect 318022 138698 318204 138934
rect 317604 103254 318204 138698
rect 317604 103018 317786 103254
rect 318022 103018 318204 103254
rect 317604 102934 318204 103018
rect 317604 102698 317786 102934
rect 318022 102698 318204 102934
rect 317459 87276 317525 87277
rect 317459 87212 317460 87276
rect 317524 87212 317525 87276
rect 317459 87211 317525 87212
rect 317462 87005 317522 87211
rect 317459 87004 317525 87005
rect 317459 86940 317460 87004
rect 317524 86940 317525 87004
rect 317459 86939 317525 86940
rect 314004 63418 314186 63654
rect 314422 63418 314604 63654
rect 314004 63334 314604 63418
rect 314004 63098 314186 63334
rect 314422 63098 314604 63334
rect 314004 27654 314604 63098
rect 317604 67254 318204 102698
rect 317604 67018 317786 67254
rect 318022 67018 318204 67254
rect 317604 66934 318204 67018
rect 317604 66698 317786 66934
rect 318022 66698 318204 66934
rect 317604 31254 318204 66698
rect 317604 31018 317786 31254
rect 318022 31018 318204 31254
rect 317604 30934 318204 31018
rect 317604 30698 317786 30934
rect 318022 30698 318204 30934
rect 315987 29612 316053 29613
rect 315987 29548 315988 29612
rect 316052 29548 316053 29612
rect 315987 29547 316053 29548
rect 315990 29205 316050 29547
rect 315987 29204 316053 29205
rect 315987 29140 315988 29204
rect 316052 29140 316053 29204
rect 315987 29139 316053 29140
rect 314004 27418 314186 27654
rect 314422 27418 314604 27654
rect 314004 27334 314604 27418
rect 314004 27098 314186 27334
rect 314422 27098 314604 27334
rect 314004 -4946 314604 27098
rect 314004 -5182 314186 -4946
rect 314422 -5182 314604 -4946
rect 314004 -5266 314604 -5182
rect 314004 -5502 314186 -5266
rect 314422 -5502 314604 -5266
rect 314004 -5524 314604 -5502
rect 299604 -6102 299786 -5866
rect 300022 -6102 300204 -5866
rect 299604 -6186 300204 -6102
rect 299604 -6422 299786 -6186
rect 300022 -6422 300204 -6186
rect 299604 -7364 300204 -6422
rect 317604 -6786 318204 30698
rect 324804 542454 325404 577898
rect 328404 690054 329004 706122
rect 328404 689818 328586 690054
rect 328822 689818 329004 690054
rect 328404 689734 329004 689818
rect 328404 689498 328586 689734
rect 328822 689498 329004 689734
rect 328404 654054 329004 689498
rect 328404 653818 328586 654054
rect 328822 653818 329004 654054
rect 328404 653734 329004 653818
rect 328404 653498 328586 653734
rect 328822 653498 329004 653734
rect 328404 618054 329004 653498
rect 328404 617818 328586 618054
rect 328822 617818 329004 618054
rect 328404 617734 329004 617818
rect 328404 617498 328586 617734
rect 328822 617498 329004 617734
rect 328404 582054 329004 617498
rect 328404 581818 328586 582054
rect 328822 581818 329004 582054
rect 328404 581734 329004 581818
rect 328404 581498 328586 581734
rect 328822 581498 329004 581734
rect 324804 542218 324986 542454
rect 325222 542218 325404 542454
rect 324804 542134 325404 542218
rect 324804 541898 324986 542134
rect 325222 541898 325404 542134
rect 324804 506454 325404 541898
rect 324804 506218 324986 506454
rect 325222 506218 325404 506454
rect 324804 506134 325404 506218
rect 324804 505898 324986 506134
rect 325222 505898 325404 506134
rect 324804 470454 325404 505898
rect 324804 470218 324986 470454
rect 325222 470218 325404 470454
rect 324804 470134 325404 470218
rect 324804 469898 324986 470134
rect 325222 469898 325404 470134
rect 324804 434454 325404 469898
rect 324804 434218 324986 434454
rect 325222 434218 325404 434454
rect 324804 434134 325404 434218
rect 324804 433898 324986 434134
rect 325222 433898 325404 434134
rect 324804 398454 325404 433898
rect 324804 398218 324986 398454
rect 325222 398218 325404 398454
rect 324804 398134 325404 398218
rect 324804 397898 324986 398134
rect 325222 397898 325404 398134
rect 324804 362454 325404 397898
rect 324804 362218 324986 362454
rect 325222 362218 325404 362454
rect 324804 362134 325404 362218
rect 324804 361898 324986 362134
rect 325222 361898 325404 362134
rect 324804 326454 325404 361898
rect 324804 326218 324986 326454
rect 325222 326218 325404 326454
rect 324804 326134 325404 326218
rect 324804 325898 324986 326134
rect 325222 325898 325404 326134
rect 324804 290454 325404 325898
rect 324804 290218 324986 290454
rect 325222 290218 325404 290454
rect 324804 290134 325404 290218
rect 324804 289898 324986 290134
rect 325222 289898 325404 290134
rect 324804 254454 325404 289898
rect 324804 254218 324986 254454
rect 325222 254218 325404 254454
rect 324804 254134 325404 254218
rect 324804 253898 324986 254134
rect 325222 253898 325404 254134
rect 324804 218454 325404 253898
rect 324804 218218 324986 218454
rect 325222 218218 325404 218454
rect 324804 218134 325404 218218
rect 324804 217898 324986 218134
rect 325222 217898 325404 218134
rect 324804 182454 325404 217898
rect 324804 182218 324986 182454
rect 325222 182218 325404 182454
rect 324804 182134 325404 182218
rect 324804 181898 324986 182134
rect 325222 181898 325404 182134
rect 324804 146454 325404 181898
rect 324804 146218 324986 146454
rect 325222 146218 325404 146454
rect 324804 146134 325404 146218
rect 324804 145898 324986 146134
rect 325222 145898 325404 146134
rect 324804 110454 325404 145898
rect 328404 546054 329004 581498
rect 328404 545818 328586 546054
rect 328822 545818 329004 546054
rect 328404 545734 329004 545818
rect 328404 545498 328586 545734
rect 328822 545498 329004 545734
rect 328404 510054 329004 545498
rect 328404 509818 328586 510054
rect 328822 509818 329004 510054
rect 328404 509734 329004 509818
rect 328404 509498 328586 509734
rect 328822 509498 329004 509734
rect 328404 474054 329004 509498
rect 328404 473818 328586 474054
rect 328822 473818 329004 474054
rect 328404 473734 329004 473818
rect 328404 473498 328586 473734
rect 328822 473498 329004 473734
rect 328404 438054 329004 473498
rect 328404 437818 328586 438054
rect 328822 437818 329004 438054
rect 328404 437734 329004 437818
rect 328404 437498 328586 437734
rect 328822 437498 329004 437734
rect 328404 402054 329004 437498
rect 328404 401818 328586 402054
rect 328822 401818 329004 402054
rect 328404 401734 329004 401818
rect 328404 401498 328586 401734
rect 328822 401498 329004 401734
rect 328404 366054 329004 401498
rect 328404 365818 328586 366054
rect 328822 365818 329004 366054
rect 328404 365734 329004 365818
rect 328404 365498 328586 365734
rect 328822 365498 329004 365734
rect 328404 330054 329004 365498
rect 328404 329818 328586 330054
rect 328822 329818 329004 330054
rect 328404 329734 329004 329818
rect 328404 329498 328586 329734
rect 328822 329498 329004 329734
rect 328404 294054 329004 329498
rect 328404 293818 328586 294054
rect 328822 293818 329004 294054
rect 328404 293734 329004 293818
rect 328404 293498 328586 293734
rect 328822 293498 329004 293734
rect 328404 258054 329004 293498
rect 328404 257818 328586 258054
rect 328822 257818 329004 258054
rect 328404 257734 329004 257818
rect 328404 257498 328586 257734
rect 328822 257498 329004 257734
rect 328404 222054 329004 257498
rect 328404 221818 328586 222054
rect 328822 221818 329004 222054
rect 328404 221734 329004 221818
rect 328404 221498 328586 221734
rect 328822 221498 329004 221734
rect 328404 186054 329004 221498
rect 328404 185818 328586 186054
rect 328822 185818 329004 186054
rect 328404 185734 329004 185818
rect 328404 185498 328586 185734
rect 328822 185498 329004 185734
rect 328404 150054 329004 185498
rect 328404 149818 328586 150054
rect 328822 149818 329004 150054
rect 328404 149734 329004 149818
rect 328404 149498 328586 149734
rect 328822 149498 329004 149734
rect 327395 138276 327461 138277
rect 327395 138212 327396 138276
rect 327460 138212 327461 138276
rect 327395 138211 327461 138212
rect 327398 135285 327458 138211
rect 327395 135284 327461 135285
rect 327395 135220 327396 135284
rect 327460 135220 327461 135284
rect 327395 135219 327461 135220
rect 324804 110218 324986 110454
rect 325222 110218 325404 110454
rect 324804 110134 325404 110218
rect 324804 109898 324986 110134
rect 325222 109898 325404 110134
rect 324804 74454 325404 109898
rect 324804 74218 324986 74454
rect 325222 74218 325404 74454
rect 324804 74134 325404 74218
rect 324804 73898 324986 74134
rect 325222 73898 325404 74134
rect 324804 38454 325404 73898
rect 324804 38218 324986 38454
rect 325222 38218 325404 38454
rect 324804 38134 325404 38218
rect 324804 37898 324986 38134
rect 325222 37898 325404 38134
rect 324804 2454 325404 37898
rect 328404 114054 329004 149498
rect 328404 113818 328586 114054
rect 328822 113818 329004 114054
rect 328404 113734 329004 113818
rect 328404 113498 328586 113734
rect 328822 113498 329004 113734
rect 328404 78054 329004 113498
rect 328404 77818 328586 78054
rect 328822 77818 329004 78054
rect 328404 77734 329004 77818
rect 328404 77498 328586 77734
rect 328822 77498 329004 77734
rect 328404 42054 329004 77498
rect 328404 41818 328586 42054
rect 328822 41818 329004 42054
rect 328404 41734 329004 41818
rect 328404 41498 328586 41734
rect 328822 41498 329004 41734
rect 327027 29204 327093 29205
rect 327027 29140 327028 29204
rect 327092 29140 327093 29204
rect 327027 29139 327093 29140
rect 327211 29204 327277 29205
rect 327211 29140 327212 29204
rect 327276 29140 327277 29204
rect 327211 29139 327277 29140
rect 327030 28930 327090 29139
rect 327214 28930 327274 29139
rect 327030 28870 327274 28930
rect 324804 2218 324986 2454
rect 325222 2218 325404 2454
rect 324804 2134 325404 2218
rect 324804 1898 324986 2134
rect 325222 1898 325404 2134
rect 324804 -346 325404 1898
rect 324804 -582 324986 -346
rect 325222 -582 325404 -346
rect 324804 -666 325404 -582
rect 324804 -902 324986 -666
rect 325222 -902 325404 -666
rect 324804 -1844 325404 -902
rect 328404 6054 329004 41498
rect 328404 5818 328586 6054
rect 328822 5818 329004 6054
rect 328404 5734 329004 5818
rect 328404 5498 328586 5734
rect 328822 5498 329004 5734
rect 328404 -2186 329004 5498
rect 328404 -2422 328586 -2186
rect 328822 -2422 329004 -2186
rect 328404 -2506 329004 -2422
rect 328404 -2742 328586 -2506
rect 328822 -2742 329004 -2506
rect 328404 -3684 329004 -2742
rect 332004 693654 332604 707962
rect 332004 693418 332186 693654
rect 332422 693418 332604 693654
rect 332004 693334 332604 693418
rect 332004 693098 332186 693334
rect 332422 693098 332604 693334
rect 332004 657654 332604 693098
rect 332004 657418 332186 657654
rect 332422 657418 332604 657654
rect 332004 657334 332604 657418
rect 332004 657098 332186 657334
rect 332422 657098 332604 657334
rect 332004 621654 332604 657098
rect 332004 621418 332186 621654
rect 332422 621418 332604 621654
rect 332004 621334 332604 621418
rect 332004 621098 332186 621334
rect 332422 621098 332604 621334
rect 332004 585654 332604 621098
rect 332004 585418 332186 585654
rect 332422 585418 332604 585654
rect 332004 585334 332604 585418
rect 332004 585098 332186 585334
rect 332422 585098 332604 585334
rect 332004 549654 332604 585098
rect 335604 697254 336204 709802
rect 353604 711278 354204 711300
rect 353604 711042 353786 711278
rect 354022 711042 354204 711278
rect 353604 710958 354204 711042
rect 353604 710722 353786 710958
rect 354022 710722 354204 710958
rect 350004 709438 350604 709460
rect 350004 709202 350186 709438
rect 350422 709202 350604 709438
rect 350004 709118 350604 709202
rect 350004 708882 350186 709118
rect 350422 708882 350604 709118
rect 346404 707598 347004 707620
rect 346404 707362 346586 707598
rect 346822 707362 347004 707598
rect 346404 707278 347004 707362
rect 346404 707042 346586 707278
rect 346822 707042 347004 707278
rect 335604 697018 335786 697254
rect 336022 697018 336204 697254
rect 335604 696934 336204 697018
rect 335604 696698 335786 696934
rect 336022 696698 336204 696934
rect 335604 661254 336204 696698
rect 335604 661018 335786 661254
rect 336022 661018 336204 661254
rect 335604 660934 336204 661018
rect 335604 660698 335786 660934
rect 336022 660698 336204 660934
rect 335604 625254 336204 660698
rect 335604 625018 335786 625254
rect 336022 625018 336204 625254
rect 335604 624934 336204 625018
rect 335604 624698 335786 624934
rect 336022 624698 336204 624934
rect 335604 589254 336204 624698
rect 335604 589018 335786 589254
rect 336022 589018 336204 589254
rect 335604 588934 336204 589018
rect 335604 588698 335786 588934
rect 336022 588698 336204 588934
rect 335126 561373 335186 562582
rect 335123 561372 335189 561373
rect 335123 561308 335124 561372
rect 335188 561308 335189 561372
rect 335123 561307 335189 561308
rect 335123 560964 335189 560965
rect 335123 560900 335124 560964
rect 335188 560900 335189 560964
rect 335123 560899 335189 560900
rect 335126 560690 335186 560899
rect 335307 560692 335373 560693
rect 335307 560690 335308 560692
rect 335126 560630 335308 560690
rect 335307 560628 335308 560630
rect 335372 560628 335373 560692
rect 335307 560627 335373 560628
rect 332004 549418 332186 549654
rect 332422 549418 332604 549654
rect 332004 549334 332604 549418
rect 332004 549098 332186 549334
rect 332422 549098 332604 549334
rect 332004 513654 332604 549098
rect 332004 513418 332186 513654
rect 332422 513418 332604 513654
rect 332004 513334 332604 513418
rect 332004 513098 332186 513334
rect 332422 513098 332604 513334
rect 332004 477654 332604 513098
rect 332004 477418 332186 477654
rect 332422 477418 332604 477654
rect 332004 477334 332604 477418
rect 332004 477098 332186 477334
rect 332422 477098 332604 477334
rect 332004 441654 332604 477098
rect 332004 441418 332186 441654
rect 332422 441418 332604 441654
rect 332004 441334 332604 441418
rect 332004 441098 332186 441334
rect 332422 441098 332604 441334
rect 332004 405654 332604 441098
rect 332004 405418 332186 405654
rect 332422 405418 332604 405654
rect 332004 405334 332604 405418
rect 332004 405098 332186 405334
rect 332422 405098 332604 405334
rect 332004 369654 332604 405098
rect 332004 369418 332186 369654
rect 332422 369418 332604 369654
rect 332004 369334 332604 369418
rect 332004 369098 332186 369334
rect 332422 369098 332604 369334
rect 332004 333654 332604 369098
rect 332004 333418 332186 333654
rect 332422 333418 332604 333654
rect 332004 333334 332604 333418
rect 332004 333098 332186 333334
rect 332422 333098 332604 333334
rect 332004 297654 332604 333098
rect 332004 297418 332186 297654
rect 332422 297418 332604 297654
rect 332004 297334 332604 297418
rect 332004 297098 332186 297334
rect 332422 297098 332604 297334
rect 332004 261654 332604 297098
rect 332004 261418 332186 261654
rect 332422 261418 332604 261654
rect 332004 261334 332604 261418
rect 332004 261098 332186 261334
rect 332422 261098 332604 261334
rect 332004 225654 332604 261098
rect 332004 225418 332186 225654
rect 332422 225418 332604 225654
rect 332004 225334 332604 225418
rect 332004 225098 332186 225334
rect 332422 225098 332604 225334
rect 332004 189654 332604 225098
rect 332004 189418 332186 189654
rect 332422 189418 332604 189654
rect 332004 189334 332604 189418
rect 332004 189098 332186 189334
rect 332422 189098 332604 189334
rect 332004 153654 332604 189098
rect 332004 153418 332186 153654
rect 332422 153418 332604 153654
rect 332004 153334 332604 153418
rect 332004 153098 332186 153334
rect 332422 153098 332604 153334
rect 332004 117654 332604 153098
rect 332004 117418 332186 117654
rect 332422 117418 332604 117654
rect 332004 117334 332604 117418
rect 332004 117098 332186 117334
rect 332422 117098 332604 117334
rect 332004 81654 332604 117098
rect 332004 81418 332186 81654
rect 332422 81418 332604 81654
rect 332004 81334 332604 81418
rect 332004 81098 332186 81334
rect 332422 81098 332604 81334
rect 332004 45654 332604 81098
rect 332004 45418 332186 45654
rect 332422 45418 332604 45654
rect 332004 45334 332604 45418
rect 332004 45098 332186 45334
rect 332422 45098 332604 45334
rect 332004 9654 332604 45098
rect 332004 9418 332186 9654
rect 332422 9418 332604 9654
rect 332004 9334 332604 9418
rect 332004 9098 332186 9334
rect 332422 9098 332604 9334
rect 332004 -4026 332604 9098
rect 332004 -4262 332186 -4026
rect 332422 -4262 332604 -4026
rect 332004 -4346 332604 -4262
rect 332004 -4582 332186 -4346
rect 332422 -4582 332604 -4346
rect 332004 -5524 332604 -4582
rect 335604 553254 336204 588698
rect 342804 705758 343404 705780
rect 342804 705522 342986 705758
rect 343222 705522 343404 705758
rect 342804 705438 343404 705522
rect 342804 705202 342986 705438
rect 343222 705202 343404 705438
rect 342804 668454 343404 705202
rect 342804 668218 342986 668454
rect 343222 668218 343404 668454
rect 342804 668134 343404 668218
rect 342804 667898 342986 668134
rect 343222 667898 343404 668134
rect 342804 632454 343404 667898
rect 342804 632218 342986 632454
rect 343222 632218 343404 632454
rect 342804 632134 343404 632218
rect 342804 631898 342986 632134
rect 343222 631898 343404 632134
rect 342804 596454 343404 631898
rect 342804 596218 342986 596454
rect 343222 596218 343404 596454
rect 342804 596134 343404 596218
rect 342804 595898 342986 596134
rect 343222 595898 343404 596134
rect 336930 562670 337394 562730
rect 337334 562138 337394 562670
rect 342804 560454 343404 595898
rect 342804 560218 342986 560454
rect 343222 560218 343404 560454
rect 342804 560134 343404 560218
rect 342804 559898 342986 560134
rect 343222 559898 343404 560134
rect 338067 559060 338133 559061
rect 338067 558996 338068 559060
rect 338132 558996 338133 559060
rect 338067 558995 338133 558996
rect 338070 558789 338130 558995
rect 338067 558788 338133 558789
rect 338067 558724 338068 558788
rect 338132 558724 338133 558788
rect 338067 558723 338133 558724
rect 335604 553018 335786 553254
rect 336022 553018 336204 553254
rect 335604 552934 336204 553018
rect 335604 552698 335786 552934
rect 336022 552698 336204 552934
rect 335604 517254 336204 552698
rect 335604 517018 335786 517254
rect 336022 517018 336204 517254
rect 335604 516934 336204 517018
rect 335604 516698 335786 516934
rect 336022 516698 336204 516934
rect 335604 481254 336204 516698
rect 335604 481018 335786 481254
rect 336022 481018 336204 481254
rect 335604 480934 336204 481018
rect 335604 480698 335786 480934
rect 336022 480698 336204 480934
rect 335604 445254 336204 480698
rect 335604 445018 335786 445254
rect 336022 445018 336204 445254
rect 335604 444934 336204 445018
rect 335604 444698 335786 444934
rect 336022 444698 336204 444934
rect 335604 409254 336204 444698
rect 335604 409018 335786 409254
rect 336022 409018 336204 409254
rect 335604 408934 336204 409018
rect 335604 408698 335786 408934
rect 336022 408698 336204 408934
rect 335604 373254 336204 408698
rect 335604 373018 335786 373254
rect 336022 373018 336204 373254
rect 335604 372934 336204 373018
rect 335604 372698 335786 372934
rect 336022 372698 336204 372934
rect 335604 337254 336204 372698
rect 335604 337018 335786 337254
rect 336022 337018 336204 337254
rect 335604 336934 336204 337018
rect 335604 336698 335786 336934
rect 336022 336698 336204 336934
rect 335604 301254 336204 336698
rect 335604 301018 335786 301254
rect 336022 301018 336204 301254
rect 335604 300934 336204 301018
rect 335604 300698 335786 300934
rect 336022 300698 336204 300934
rect 335604 265254 336204 300698
rect 335604 265018 335786 265254
rect 336022 265018 336204 265254
rect 335604 264934 336204 265018
rect 335604 264698 335786 264934
rect 336022 264698 336204 264934
rect 335604 229254 336204 264698
rect 335604 229018 335786 229254
rect 336022 229018 336204 229254
rect 335604 228934 336204 229018
rect 335604 228698 335786 228934
rect 336022 228698 336204 228934
rect 335604 193254 336204 228698
rect 335604 193018 335786 193254
rect 336022 193018 336204 193254
rect 335604 192934 336204 193018
rect 335604 192698 335786 192934
rect 336022 192698 336204 192934
rect 335604 157254 336204 192698
rect 335604 157018 335786 157254
rect 336022 157018 336204 157254
rect 335604 156934 336204 157018
rect 335604 156698 335786 156934
rect 336022 156698 336204 156934
rect 335604 121254 336204 156698
rect 335604 121018 335786 121254
rect 336022 121018 336204 121254
rect 335604 120934 336204 121018
rect 335604 120698 335786 120934
rect 336022 120698 336204 120934
rect 335604 85254 336204 120698
rect 335604 85018 335786 85254
rect 336022 85018 336204 85254
rect 335604 84934 336204 85018
rect 335604 84698 335786 84934
rect 336022 84698 336204 84934
rect 335604 49254 336204 84698
rect 335604 49018 335786 49254
rect 336022 49018 336204 49254
rect 335604 48934 336204 49018
rect 335604 48698 335786 48934
rect 336022 48698 336204 48934
rect 335604 13254 336204 48698
rect 335604 13018 335786 13254
rect 336022 13018 336204 13254
rect 335604 12934 336204 13018
rect 335604 12698 335786 12934
rect 336022 12698 336204 12934
rect 317604 -7022 317786 -6786
rect 318022 -7022 318204 -6786
rect 317604 -7106 318204 -7022
rect 317604 -7342 317786 -7106
rect 318022 -7342 318204 -7106
rect 317604 -7364 318204 -7342
rect 335604 -5866 336204 12698
rect 342804 524454 343404 559898
rect 342804 524218 342986 524454
rect 343222 524218 343404 524454
rect 342804 524134 343404 524218
rect 342804 523898 342986 524134
rect 343222 523898 343404 524134
rect 342804 488454 343404 523898
rect 342804 488218 342986 488454
rect 343222 488218 343404 488454
rect 342804 488134 343404 488218
rect 342804 487898 342986 488134
rect 343222 487898 343404 488134
rect 342804 452454 343404 487898
rect 342804 452218 342986 452454
rect 343222 452218 343404 452454
rect 342804 452134 343404 452218
rect 342804 451898 342986 452134
rect 343222 451898 343404 452134
rect 342804 416454 343404 451898
rect 342804 416218 342986 416454
rect 343222 416218 343404 416454
rect 342804 416134 343404 416218
rect 342804 415898 342986 416134
rect 343222 415898 343404 416134
rect 342804 380454 343404 415898
rect 342804 380218 342986 380454
rect 343222 380218 343404 380454
rect 342804 380134 343404 380218
rect 342804 379898 342986 380134
rect 343222 379898 343404 380134
rect 342804 344454 343404 379898
rect 342804 344218 342986 344454
rect 343222 344218 343404 344454
rect 342804 344134 343404 344218
rect 342804 343898 342986 344134
rect 343222 343898 343404 344134
rect 342804 308454 343404 343898
rect 342804 308218 342986 308454
rect 343222 308218 343404 308454
rect 342804 308134 343404 308218
rect 342804 307898 342986 308134
rect 343222 307898 343404 308134
rect 342804 272454 343404 307898
rect 342804 272218 342986 272454
rect 343222 272218 343404 272454
rect 342804 272134 343404 272218
rect 342804 271898 342986 272134
rect 343222 271898 343404 272134
rect 342804 236454 343404 271898
rect 342804 236218 342986 236454
rect 343222 236218 343404 236454
rect 342804 236134 343404 236218
rect 342804 235898 342986 236134
rect 343222 235898 343404 236134
rect 342804 200454 343404 235898
rect 342804 200218 342986 200454
rect 343222 200218 343404 200454
rect 342804 200134 343404 200218
rect 342804 199898 342986 200134
rect 343222 199898 343404 200134
rect 342804 164454 343404 199898
rect 342804 164218 342986 164454
rect 343222 164218 343404 164454
rect 342804 164134 343404 164218
rect 342804 163898 342986 164134
rect 343222 163898 343404 164134
rect 342804 128454 343404 163898
rect 342804 128218 342986 128454
rect 343222 128218 343404 128454
rect 342804 128134 343404 128218
rect 342804 127898 342986 128134
rect 343222 127898 343404 128134
rect 342804 92454 343404 127898
rect 342804 92218 342986 92454
rect 343222 92218 343404 92454
rect 342804 92134 343404 92218
rect 342804 91898 342986 92134
rect 343222 91898 343404 92134
rect 342804 56454 343404 91898
rect 346404 672054 347004 707042
rect 346404 671818 346586 672054
rect 346822 671818 347004 672054
rect 346404 671734 347004 671818
rect 346404 671498 346586 671734
rect 346822 671498 347004 671734
rect 346404 636054 347004 671498
rect 346404 635818 346586 636054
rect 346822 635818 347004 636054
rect 346404 635734 347004 635818
rect 346404 635498 346586 635734
rect 346822 635498 347004 635734
rect 346404 600054 347004 635498
rect 346404 599818 346586 600054
rect 346822 599818 347004 600054
rect 346404 599734 347004 599818
rect 346404 599498 346586 599734
rect 346822 599498 347004 599734
rect 346404 564054 347004 599498
rect 346404 563818 346586 564054
rect 346822 563818 347004 564054
rect 346404 563734 347004 563818
rect 346404 563498 346586 563734
rect 346822 563498 347004 563734
rect 346404 528054 347004 563498
rect 346404 527818 346586 528054
rect 346822 527818 347004 528054
rect 346404 527734 347004 527818
rect 346404 527498 346586 527734
rect 346822 527498 347004 527734
rect 346404 492054 347004 527498
rect 346404 491818 346586 492054
rect 346822 491818 347004 492054
rect 346404 491734 347004 491818
rect 346404 491498 346586 491734
rect 346822 491498 347004 491734
rect 346404 456054 347004 491498
rect 346404 455818 346586 456054
rect 346822 455818 347004 456054
rect 346404 455734 347004 455818
rect 346404 455498 346586 455734
rect 346822 455498 347004 455734
rect 346404 420054 347004 455498
rect 346404 419818 346586 420054
rect 346822 419818 347004 420054
rect 346404 419734 347004 419818
rect 346404 419498 346586 419734
rect 346822 419498 347004 419734
rect 346404 384054 347004 419498
rect 346404 383818 346586 384054
rect 346822 383818 347004 384054
rect 346404 383734 347004 383818
rect 346404 383498 346586 383734
rect 346822 383498 347004 383734
rect 346404 348054 347004 383498
rect 346404 347818 346586 348054
rect 346822 347818 347004 348054
rect 346404 347734 347004 347818
rect 346404 347498 346586 347734
rect 346822 347498 347004 347734
rect 346404 312054 347004 347498
rect 346404 311818 346586 312054
rect 346822 311818 347004 312054
rect 346404 311734 347004 311818
rect 346404 311498 346586 311734
rect 346822 311498 347004 311734
rect 346404 276054 347004 311498
rect 346404 275818 346586 276054
rect 346822 275818 347004 276054
rect 346404 275734 347004 275818
rect 346404 275498 346586 275734
rect 346822 275498 347004 275734
rect 346404 240054 347004 275498
rect 346404 239818 346586 240054
rect 346822 239818 347004 240054
rect 346404 239734 347004 239818
rect 346404 239498 346586 239734
rect 346822 239498 347004 239734
rect 346404 204054 347004 239498
rect 346404 203818 346586 204054
rect 346822 203818 347004 204054
rect 346404 203734 347004 203818
rect 346404 203498 346586 203734
rect 346822 203498 347004 203734
rect 346404 168054 347004 203498
rect 346404 167818 346586 168054
rect 346822 167818 347004 168054
rect 346404 167734 347004 167818
rect 346404 167498 346586 167734
rect 346822 167498 347004 167734
rect 346404 132054 347004 167498
rect 346404 131818 346586 132054
rect 346822 131818 347004 132054
rect 346404 131734 347004 131818
rect 346404 131498 346586 131734
rect 346822 131498 347004 131734
rect 346404 96054 347004 131498
rect 346404 95818 346586 96054
rect 346822 95818 347004 96054
rect 346404 95734 347004 95818
rect 346404 95498 346586 95734
rect 346822 95498 347004 95734
rect 343587 64020 343653 64021
rect 343587 63956 343588 64020
rect 343652 63956 343653 64020
rect 343587 63955 343653 63956
rect 343590 63749 343650 63955
rect 343587 63748 343653 63749
rect 343587 63684 343588 63748
rect 343652 63684 343653 63748
rect 343587 63683 343653 63684
rect 342804 56218 342986 56454
rect 343222 56218 343404 56454
rect 342804 56134 343404 56218
rect 342804 55898 342986 56134
rect 343222 55898 343404 56134
rect 342804 20454 343404 55898
rect 342804 20218 342986 20454
rect 343222 20218 343404 20454
rect 342804 20134 343404 20218
rect 342804 19898 342986 20134
rect 343222 19898 343404 20134
rect 342804 -1266 343404 19898
rect 342804 -1502 342986 -1266
rect 343222 -1502 343404 -1266
rect 342804 -1586 343404 -1502
rect 342804 -1822 342986 -1586
rect 343222 -1822 343404 -1586
rect 342804 -1844 343404 -1822
rect 346404 60054 347004 95498
rect 346404 59818 346586 60054
rect 346822 59818 347004 60054
rect 346404 59734 347004 59818
rect 346404 59498 346586 59734
rect 346822 59498 347004 59734
rect 346404 24054 347004 59498
rect 346404 23818 346586 24054
rect 346822 23818 347004 24054
rect 346404 23734 347004 23818
rect 346404 23498 346586 23734
rect 346822 23498 347004 23734
rect 346404 -3106 347004 23498
rect 346404 -3342 346586 -3106
rect 346822 -3342 347004 -3106
rect 346404 -3426 347004 -3342
rect 346404 -3662 346586 -3426
rect 346822 -3662 347004 -3426
rect 346404 -3684 347004 -3662
rect 350004 675654 350604 708882
rect 350004 675418 350186 675654
rect 350422 675418 350604 675654
rect 350004 675334 350604 675418
rect 350004 675098 350186 675334
rect 350422 675098 350604 675334
rect 350004 639654 350604 675098
rect 350004 639418 350186 639654
rect 350422 639418 350604 639654
rect 350004 639334 350604 639418
rect 350004 639098 350186 639334
rect 350422 639098 350604 639334
rect 350004 603654 350604 639098
rect 350004 603418 350186 603654
rect 350422 603418 350604 603654
rect 350004 603334 350604 603418
rect 350004 603098 350186 603334
rect 350422 603098 350604 603334
rect 350004 567654 350604 603098
rect 350004 567418 350186 567654
rect 350422 567418 350604 567654
rect 350004 567334 350604 567418
rect 350004 567098 350186 567334
rect 350422 567098 350604 567334
rect 350004 531654 350604 567098
rect 353604 679254 354204 710722
rect 371604 710358 372204 711300
rect 371604 710122 371786 710358
rect 372022 710122 372204 710358
rect 371604 710038 372204 710122
rect 371604 709802 371786 710038
rect 372022 709802 372204 710038
rect 368004 708518 368604 709460
rect 368004 708282 368186 708518
rect 368422 708282 368604 708518
rect 368004 708198 368604 708282
rect 368004 707962 368186 708198
rect 368422 707962 368604 708198
rect 364404 706678 365004 707620
rect 364404 706442 364586 706678
rect 364822 706442 365004 706678
rect 364404 706358 365004 706442
rect 364404 706122 364586 706358
rect 364822 706122 365004 706358
rect 353604 679018 353786 679254
rect 354022 679018 354204 679254
rect 353604 678934 354204 679018
rect 353604 678698 353786 678934
rect 354022 678698 354204 678934
rect 353604 643254 354204 678698
rect 353604 643018 353786 643254
rect 354022 643018 354204 643254
rect 353604 642934 354204 643018
rect 353604 642698 353786 642934
rect 354022 642698 354204 642934
rect 353604 607254 354204 642698
rect 353604 607018 353786 607254
rect 354022 607018 354204 607254
rect 353604 606934 354204 607018
rect 353604 606698 353786 606934
rect 354022 606698 354204 606934
rect 353604 571254 354204 606698
rect 353604 571018 353786 571254
rect 354022 571018 354204 571254
rect 353604 570934 354204 571018
rect 353604 570698 353786 570934
rect 354022 570698 354204 570934
rect 351870 559270 352114 559330
rect 351870 559061 351930 559270
rect 352054 559197 352114 559270
rect 352051 559196 352117 559197
rect 352051 559132 352052 559196
rect 352116 559132 352117 559196
rect 352051 559131 352117 559132
rect 351867 559060 351933 559061
rect 351867 558996 351868 559060
rect 351932 558996 351933 559060
rect 351867 558995 351933 558996
rect 350004 531418 350186 531654
rect 350422 531418 350604 531654
rect 350004 531334 350604 531418
rect 350004 531098 350186 531334
rect 350422 531098 350604 531334
rect 350004 495654 350604 531098
rect 350004 495418 350186 495654
rect 350422 495418 350604 495654
rect 350004 495334 350604 495418
rect 350004 495098 350186 495334
rect 350422 495098 350604 495334
rect 350004 459654 350604 495098
rect 350004 459418 350186 459654
rect 350422 459418 350604 459654
rect 350004 459334 350604 459418
rect 350004 459098 350186 459334
rect 350422 459098 350604 459334
rect 350004 423654 350604 459098
rect 350004 423418 350186 423654
rect 350422 423418 350604 423654
rect 350004 423334 350604 423418
rect 350004 423098 350186 423334
rect 350422 423098 350604 423334
rect 350004 387654 350604 423098
rect 350004 387418 350186 387654
rect 350422 387418 350604 387654
rect 350004 387334 350604 387418
rect 350004 387098 350186 387334
rect 350422 387098 350604 387334
rect 350004 351654 350604 387098
rect 350004 351418 350186 351654
rect 350422 351418 350604 351654
rect 350004 351334 350604 351418
rect 350004 351098 350186 351334
rect 350422 351098 350604 351334
rect 350004 315654 350604 351098
rect 350004 315418 350186 315654
rect 350422 315418 350604 315654
rect 350004 315334 350604 315418
rect 350004 315098 350186 315334
rect 350422 315098 350604 315334
rect 350004 279654 350604 315098
rect 350004 279418 350186 279654
rect 350422 279418 350604 279654
rect 350004 279334 350604 279418
rect 350004 279098 350186 279334
rect 350422 279098 350604 279334
rect 350004 243654 350604 279098
rect 350004 243418 350186 243654
rect 350422 243418 350604 243654
rect 350004 243334 350604 243418
rect 350004 243098 350186 243334
rect 350422 243098 350604 243334
rect 350004 207654 350604 243098
rect 350004 207418 350186 207654
rect 350422 207418 350604 207654
rect 350004 207334 350604 207418
rect 350004 207098 350186 207334
rect 350422 207098 350604 207334
rect 350004 171654 350604 207098
rect 350004 171418 350186 171654
rect 350422 171418 350604 171654
rect 350004 171334 350604 171418
rect 350004 171098 350186 171334
rect 350422 171098 350604 171334
rect 350004 135654 350604 171098
rect 350004 135418 350186 135654
rect 350422 135418 350604 135654
rect 350004 135334 350604 135418
rect 350004 135098 350186 135334
rect 350422 135098 350604 135334
rect 350004 99654 350604 135098
rect 350004 99418 350186 99654
rect 350422 99418 350604 99654
rect 350004 99334 350604 99418
rect 350004 99098 350186 99334
rect 350422 99098 350604 99334
rect 350004 63654 350604 99098
rect 350004 63418 350186 63654
rect 350422 63418 350604 63654
rect 350004 63334 350604 63418
rect 350004 63098 350186 63334
rect 350422 63098 350604 63334
rect 350004 27654 350604 63098
rect 350004 27418 350186 27654
rect 350422 27418 350604 27654
rect 350004 27334 350604 27418
rect 350004 27098 350186 27334
rect 350422 27098 350604 27334
rect 350004 -4946 350604 27098
rect 350004 -5182 350186 -4946
rect 350422 -5182 350604 -4946
rect 350004 -5266 350604 -5182
rect 350004 -5502 350186 -5266
rect 350422 -5502 350604 -5266
rect 350004 -5524 350604 -5502
rect 353604 535254 354204 570698
rect 360804 704838 361404 705780
rect 360804 704602 360986 704838
rect 361222 704602 361404 704838
rect 360804 704518 361404 704602
rect 360804 704282 360986 704518
rect 361222 704282 361404 704518
rect 360804 686454 361404 704282
rect 360804 686218 360986 686454
rect 361222 686218 361404 686454
rect 360804 686134 361404 686218
rect 360804 685898 360986 686134
rect 361222 685898 361404 686134
rect 360804 650454 361404 685898
rect 360804 650218 360986 650454
rect 361222 650218 361404 650454
rect 360804 650134 361404 650218
rect 360804 649898 360986 650134
rect 361222 649898 361404 650134
rect 360804 614454 361404 649898
rect 360804 614218 360986 614454
rect 361222 614218 361404 614454
rect 360804 614134 361404 614218
rect 360804 613898 360986 614134
rect 361222 613898 361404 614134
rect 360804 578454 361404 613898
rect 360804 578218 360986 578454
rect 361222 578218 361404 578454
rect 360804 578134 361404 578218
rect 360804 577898 360986 578134
rect 361222 577898 361404 578134
rect 357387 563140 357453 563141
rect 357387 563076 357388 563140
rect 357452 563076 357453 563140
rect 357387 563075 357453 563076
rect 357390 562818 357450 563075
rect 357387 560828 357453 560829
rect 357387 560764 357388 560828
rect 357452 560764 357453 560828
rect 357387 560763 357453 560764
rect 357390 560557 357450 560763
rect 357387 560556 357453 560557
rect 357387 560492 357388 560556
rect 357452 560492 357453 560556
rect 357387 560491 357453 560492
rect 353604 535018 353786 535254
rect 354022 535018 354204 535254
rect 353604 534934 354204 535018
rect 353604 534698 353786 534934
rect 354022 534698 354204 534934
rect 353604 499254 354204 534698
rect 353604 499018 353786 499254
rect 354022 499018 354204 499254
rect 353604 498934 354204 499018
rect 353604 498698 353786 498934
rect 354022 498698 354204 498934
rect 353604 463254 354204 498698
rect 353604 463018 353786 463254
rect 354022 463018 354204 463254
rect 353604 462934 354204 463018
rect 353604 462698 353786 462934
rect 354022 462698 354204 462934
rect 353604 427254 354204 462698
rect 353604 427018 353786 427254
rect 354022 427018 354204 427254
rect 353604 426934 354204 427018
rect 353604 426698 353786 426934
rect 354022 426698 354204 426934
rect 353604 391254 354204 426698
rect 353604 391018 353786 391254
rect 354022 391018 354204 391254
rect 353604 390934 354204 391018
rect 353604 390698 353786 390934
rect 354022 390698 354204 390934
rect 353604 355254 354204 390698
rect 353604 355018 353786 355254
rect 354022 355018 354204 355254
rect 353604 354934 354204 355018
rect 353604 354698 353786 354934
rect 354022 354698 354204 354934
rect 353604 319254 354204 354698
rect 353604 319018 353786 319254
rect 354022 319018 354204 319254
rect 353604 318934 354204 319018
rect 353604 318698 353786 318934
rect 354022 318698 354204 318934
rect 353604 283254 354204 318698
rect 353604 283018 353786 283254
rect 354022 283018 354204 283254
rect 353604 282934 354204 283018
rect 353604 282698 353786 282934
rect 354022 282698 354204 282934
rect 353604 247254 354204 282698
rect 353604 247018 353786 247254
rect 354022 247018 354204 247254
rect 353604 246934 354204 247018
rect 353604 246698 353786 246934
rect 354022 246698 354204 246934
rect 353604 211254 354204 246698
rect 353604 211018 353786 211254
rect 354022 211018 354204 211254
rect 353604 210934 354204 211018
rect 353604 210698 353786 210934
rect 354022 210698 354204 210934
rect 353604 175254 354204 210698
rect 360804 542454 361404 577898
rect 360804 542218 360986 542454
rect 361222 542218 361404 542454
rect 360804 542134 361404 542218
rect 360804 541898 360986 542134
rect 361222 541898 361404 542134
rect 360804 506454 361404 541898
rect 360804 506218 360986 506454
rect 361222 506218 361404 506454
rect 360804 506134 361404 506218
rect 360804 505898 360986 506134
rect 361222 505898 361404 506134
rect 360804 470454 361404 505898
rect 360804 470218 360986 470454
rect 361222 470218 361404 470454
rect 360804 470134 361404 470218
rect 360804 469898 360986 470134
rect 361222 469898 361404 470134
rect 360804 434454 361404 469898
rect 360804 434218 360986 434454
rect 361222 434218 361404 434454
rect 360804 434134 361404 434218
rect 360804 433898 360986 434134
rect 361222 433898 361404 434134
rect 360804 398454 361404 433898
rect 360804 398218 360986 398454
rect 361222 398218 361404 398454
rect 360804 398134 361404 398218
rect 360804 397898 360986 398134
rect 361222 397898 361404 398134
rect 360804 362454 361404 397898
rect 360804 362218 360986 362454
rect 361222 362218 361404 362454
rect 360804 362134 361404 362218
rect 360804 361898 360986 362134
rect 361222 361898 361404 362134
rect 360804 326454 361404 361898
rect 360804 326218 360986 326454
rect 361222 326218 361404 326454
rect 360804 326134 361404 326218
rect 360804 325898 360986 326134
rect 361222 325898 361404 326134
rect 360804 290454 361404 325898
rect 360804 290218 360986 290454
rect 361222 290218 361404 290454
rect 360804 290134 361404 290218
rect 360804 289898 360986 290134
rect 361222 289898 361404 290134
rect 360804 254454 361404 289898
rect 360804 254218 360986 254454
rect 361222 254218 361404 254454
rect 360804 254134 361404 254218
rect 360804 253898 360986 254134
rect 361222 253898 361404 254134
rect 360804 218454 361404 253898
rect 360804 218218 360986 218454
rect 361222 218218 361404 218454
rect 360804 218134 361404 218218
rect 360804 217898 360986 218134
rect 361222 217898 361404 218134
rect 360804 182454 361404 217898
rect 360804 182218 360986 182454
rect 361222 182218 361404 182454
rect 360804 182134 361404 182218
rect 360804 181898 360986 182134
rect 361222 181898 361404 182134
rect 357387 181524 357453 181525
rect 357387 181460 357388 181524
rect 357452 181460 357453 181524
rect 357387 181459 357453 181460
rect 357390 181253 357450 181459
rect 357387 181252 357453 181253
rect 357387 181188 357388 181252
rect 357452 181188 357453 181252
rect 357387 181187 357453 181188
rect 353604 175018 353786 175254
rect 354022 175018 354204 175254
rect 353604 174934 354204 175018
rect 353604 174698 353786 174934
rect 354022 174698 354204 174934
rect 353604 139254 354204 174698
rect 353604 139018 353786 139254
rect 354022 139018 354204 139254
rect 353604 138934 354204 139018
rect 353604 138698 353786 138934
rect 354022 138698 354204 138934
rect 353604 103254 354204 138698
rect 353604 103018 353786 103254
rect 354022 103018 354204 103254
rect 353604 102934 354204 103018
rect 353604 102698 353786 102934
rect 354022 102698 354204 102934
rect 353604 67254 354204 102698
rect 353604 67018 353786 67254
rect 354022 67018 354204 67254
rect 353604 66934 354204 67018
rect 353604 66698 353786 66934
rect 354022 66698 354204 66934
rect 353604 31254 354204 66698
rect 353604 31018 353786 31254
rect 354022 31018 354204 31254
rect 353604 30934 354204 31018
rect 353604 30698 353786 30934
rect 354022 30698 354204 30934
rect 335604 -6102 335786 -5866
rect 336022 -6102 336204 -5866
rect 335604 -6186 336204 -6102
rect 335604 -6422 335786 -6186
rect 336022 -6422 336204 -6186
rect 335604 -7364 336204 -6422
rect 353604 -6786 354204 30698
rect 360804 146454 361404 181898
rect 360804 146218 360986 146454
rect 361222 146218 361404 146454
rect 360804 146134 361404 146218
rect 360804 145898 360986 146134
rect 361222 145898 361404 146134
rect 360804 110454 361404 145898
rect 360804 110218 360986 110454
rect 361222 110218 361404 110454
rect 360804 110134 361404 110218
rect 360804 109898 360986 110134
rect 361222 109898 361404 110134
rect 360804 74454 361404 109898
rect 360804 74218 360986 74454
rect 361222 74218 361404 74454
rect 360804 74134 361404 74218
rect 360804 73898 360986 74134
rect 361222 73898 361404 74134
rect 360804 38454 361404 73898
rect 360804 38218 360986 38454
rect 361222 38218 361404 38454
rect 360804 38134 361404 38218
rect 360804 37898 360986 38134
rect 361222 37898 361404 38134
rect 360804 2454 361404 37898
rect 360804 2218 360986 2454
rect 361222 2218 361404 2454
rect 360804 2134 361404 2218
rect 360804 1898 360986 2134
rect 361222 1898 361404 2134
rect 360804 -346 361404 1898
rect 360804 -582 360986 -346
rect 361222 -582 361404 -346
rect 360804 -666 361404 -582
rect 360804 -902 360986 -666
rect 361222 -902 361404 -666
rect 360804 -1844 361404 -902
rect 364404 690054 365004 706122
rect 364404 689818 364586 690054
rect 364822 689818 365004 690054
rect 364404 689734 365004 689818
rect 364404 689498 364586 689734
rect 364822 689498 365004 689734
rect 364404 654054 365004 689498
rect 364404 653818 364586 654054
rect 364822 653818 365004 654054
rect 364404 653734 365004 653818
rect 364404 653498 364586 653734
rect 364822 653498 365004 653734
rect 364404 618054 365004 653498
rect 364404 617818 364586 618054
rect 364822 617818 365004 618054
rect 364404 617734 365004 617818
rect 364404 617498 364586 617734
rect 364822 617498 365004 617734
rect 364404 582054 365004 617498
rect 364404 581818 364586 582054
rect 364822 581818 365004 582054
rect 364404 581734 365004 581818
rect 364404 581498 364586 581734
rect 364822 581498 365004 581734
rect 364404 546054 365004 581498
rect 368004 693654 368604 707962
rect 368004 693418 368186 693654
rect 368422 693418 368604 693654
rect 368004 693334 368604 693418
rect 368004 693098 368186 693334
rect 368422 693098 368604 693334
rect 368004 657654 368604 693098
rect 368004 657418 368186 657654
rect 368422 657418 368604 657654
rect 368004 657334 368604 657418
rect 368004 657098 368186 657334
rect 368422 657098 368604 657334
rect 368004 621654 368604 657098
rect 368004 621418 368186 621654
rect 368422 621418 368604 621654
rect 368004 621334 368604 621418
rect 368004 621098 368186 621334
rect 368422 621098 368604 621334
rect 368004 585654 368604 621098
rect 368004 585418 368186 585654
rect 368422 585418 368604 585654
rect 368004 585334 368604 585418
rect 368004 585098 368186 585334
rect 368422 585098 368604 585334
rect 366955 563140 367021 563141
rect 366955 563076 366956 563140
rect 367020 563076 367021 563140
rect 366955 563075 367021 563076
rect 366958 562138 367018 563075
rect 364404 545818 364586 546054
rect 364822 545818 365004 546054
rect 364404 545734 365004 545818
rect 364404 545498 364586 545734
rect 364822 545498 365004 545734
rect 364404 510054 365004 545498
rect 364404 509818 364586 510054
rect 364822 509818 365004 510054
rect 364404 509734 365004 509818
rect 364404 509498 364586 509734
rect 364822 509498 365004 509734
rect 364404 474054 365004 509498
rect 364404 473818 364586 474054
rect 364822 473818 365004 474054
rect 364404 473734 365004 473818
rect 364404 473498 364586 473734
rect 364822 473498 365004 473734
rect 364404 438054 365004 473498
rect 364404 437818 364586 438054
rect 364822 437818 365004 438054
rect 364404 437734 365004 437818
rect 364404 437498 364586 437734
rect 364822 437498 365004 437734
rect 364404 402054 365004 437498
rect 364404 401818 364586 402054
rect 364822 401818 365004 402054
rect 364404 401734 365004 401818
rect 364404 401498 364586 401734
rect 364822 401498 365004 401734
rect 364404 366054 365004 401498
rect 364404 365818 364586 366054
rect 364822 365818 365004 366054
rect 364404 365734 365004 365818
rect 364404 365498 364586 365734
rect 364822 365498 365004 365734
rect 364404 330054 365004 365498
rect 364404 329818 364586 330054
rect 364822 329818 365004 330054
rect 364404 329734 365004 329818
rect 364404 329498 364586 329734
rect 364822 329498 365004 329734
rect 364404 294054 365004 329498
rect 364404 293818 364586 294054
rect 364822 293818 365004 294054
rect 364404 293734 365004 293818
rect 364404 293498 364586 293734
rect 364822 293498 365004 293734
rect 364404 258054 365004 293498
rect 364404 257818 364586 258054
rect 364822 257818 365004 258054
rect 364404 257734 365004 257818
rect 364404 257498 364586 257734
rect 364822 257498 365004 257734
rect 364404 222054 365004 257498
rect 364404 221818 364586 222054
rect 364822 221818 365004 222054
rect 364404 221734 365004 221818
rect 364404 221498 364586 221734
rect 364822 221498 365004 221734
rect 364404 186054 365004 221498
rect 364404 185818 364586 186054
rect 364822 185818 365004 186054
rect 364404 185734 365004 185818
rect 364404 185498 364586 185734
rect 364822 185498 365004 185734
rect 364404 150054 365004 185498
rect 364404 149818 364586 150054
rect 364822 149818 365004 150054
rect 364404 149734 365004 149818
rect 364404 149498 364586 149734
rect 364822 149498 365004 149734
rect 364404 114054 365004 149498
rect 364404 113818 364586 114054
rect 364822 113818 365004 114054
rect 364404 113734 365004 113818
rect 364404 113498 364586 113734
rect 364822 113498 365004 113734
rect 364404 78054 365004 113498
rect 368004 549654 368604 585098
rect 371604 697254 372204 709802
rect 389604 711278 390204 711300
rect 389604 711042 389786 711278
rect 390022 711042 390204 711278
rect 389604 710958 390204 711042
rect 389604 710722 389786 710958
rect 390022 710722 390204 710958
rect 386004 709438 386604 709460
rect 386004 709202 386186 709438
rect 386422 709202 386604 709438
rect 386004 709118 386604 709202
rect 386004 708882 386186 709118
rect 386422 708882 386604 709118
rect 382404 707598 383004 707620
rect 382404 707362 382586 707598
rect 382822 707362 383004 707598
rect 382404 707278 383004 707362
rect 382404 707042 382586 707278
rect 382822 707042 383004 707278
rect 371604 697018 371786 697254
rect 372022 697018 372204 697254
rect 371604 696934 372204 697018
rect 371604 696698 371786 696934
rect 372022 696698 372204 696934
rect 371604 661254 372204 696698
rect 371604 661018 371786 661254
rect 372022 661018 372204 661254
rect 371604 660934 372204 661018
rect 371604 660698 371786 660934
rect 372022 660698 372204 660934
rect 371604 625254 372204 660698
rect 371604 625018 371786 625254
rect 372022 625018 372204 625254
rect 371604 624934 372204 625018
rect 371604 624698 371786 624934
rect 372022 624698 372204 624934
rect 371604 589254 372204 624698
rect 371604 589018 371786 589254
rect 372022 589018 372204 589254
rect 371604 588934 372204 589018
rect 371604 588698 371786 588934
rect 372022 588698 372204 588934
rect 369350 562670 370366 562730
rect 369350 562138 369410 562670
rect 368004 549418 368186 549654
rect 368422 549418 368604 549654
rect 368004 549334 368604 549418
rect 368004 549098 368186 549334
rect 368422 549098 368604 549334
rect 368004 513654 368604 549098
rect 368004 513418 368186 513654
rect 368422 513418 368604 513654
rect 368004 513334 368604 513418
rect 368004 513098 368186 513334
rect 368422 513098 368604 513334
rect 368004 477654 368604 513098
rect 368004 477418 368186 477654
rect 368422 477418 368604 477654
rect 368004 477334 368604 477418
rect 368004 477098 368186 477334
rect 368422 477098 368604 477334
rect 368004 441654 368604 477098
rect 368004 441418 368186 441654
rect 368422 441418 368604 441654
rect 368004 441334 368604 441418
rect 368004 441098 368186 441334
rect 368422 441098 368604 441334
rect 368004 405654 368604 441098
rect 368004 405418 368186 405654
rect 368422 405418 368604 405654
rect 368004 405334 368604 405418
rect 368004 405098 368186 405334
rect 368422 405098 368604 405334
rect 368004 369654 368604 405098
rect 368004 369418 368186 369654
rect 368422 369418 368604 369654
rect 368004 369334 368604 369418
rect 368004 369098 368186 369334
rect 368422 369098 368604 369334
rect 368004 333654 368604 369098
rect 368004 333418 368186 333654
rect 368422 333418 368604 333654
rect 368004 333334 368604 333418
rect 368004 333098 368186 333334
rect 368422 333098 368604 333334
rect 368004 297654 368604 333098
rect 368004 297418 368186 297654
rect 368422 297418 368604 297654
rect 368004 297334 368604 297418
rect 368004 297098 368186 297334
rect 368422 297098 368604 297334
rect 368004 261654 368604 297098
rect 368004 261418 368186 261654
rect 368422 261418 368604 261654
rect 368004 261334 368604 261418
rect 368004 261098 368186 261334
rect 368422 261098 368604 261334
rect 368004 225654 368604 261098
rect 368004 225418 368186 225654
rect 368422 225418 368604 225654
rect 368004 225334 368604 225418
rect 368004 225098 368186 225334
rect 368422 225098 368604 225334
rect 368004 189654 368604 225098
rect 368004 189418 368186 189654
rect 368422 189418 368604 189654
rect 368004 189334 368604 189418
rect 368004 189098 368186 189334
rect 368422 189098 368604 189334
rect 368004 153654 368604 189098
rect 368004 153418 368186 153654
rect 368422 153418 368604 153654
rect 368004 153334 368604 153418
rect 368004 153098 368186 153334
rect 368422 153098 368604 153334
rect 368004 117654 368604 153098
rect 368004 117418 368186 117654
rect 368422 117418 368604 117654
rect 368004 117334 368604 117418
rect 368004 117098 368186 117334
rect 368422 117098 368604 117334
rect 366955 87412 367021 87413
rect 366955 87348 366956 87412
rect 367020 87348 367021 87412
rect 366955 87347 367021 87348
rect 366958 87005 367018 87347
rect 366955 87004 367021 87005
rect 366955 86940 366956 87004
rect 367020 86940 367021 87004
rect 366955 86939 367021 86940
rect 364404 77818 364586 78054
rect 364822 77818 365004 78054
rect 364404 77734 365004 77818
rect 364404 77498 364586 77734
rect 364822 77498 365004 77734
rect 364404 42054 365004 77498
rect 364404 41818 364586 42054
rect 364822 41818 365004 42054
rect 364404 41734 365004 41818
rect 364404 41498 364586 41734
rect 364822 41498 365004 41734
rect 364404 6054 365004 41498
rect 368004 81654 368604 117098
rect 368004 81418 368186 81654
rect 368422 81418 368604 81654
rect 368004 81334 368604 81418
rect 368004 81098 368186 81334
rect 368422 81098 368604 81334
rect 368004 45654 368604 81098
rect 368004 45418 368186 45654
rect 368422 45418 368604 45654
rect 368004 45334 368604 45418
rect 368004 45098 368186 45334
rect 368422 45098 368604 45334
rect 366955 29340 367021 29341
rect 366955 29276 366956 29340
rect 367020 29276 367021 29340
rect 366955 29275 367021 29276
rect 366958 29069 367018 29275
rect 366955 29068 367021 29069
rect 366955 29004 366956 29068
rect 367020 29004 367021 29068
rect 366955 29003 367021 29004
rect 364404 5818 364586 6054
rect 364822 5818 365004 6054
rect 364404 5734 365004 5818
rect 364404 5498 364586 5734
rect 364822 5498 365004 5734
rect 364404 -2186 365004 5498
rect 364404 -2422 364586 -2186
rect 364822 -2422 365004 -2186
rect 364404 -2506 365004 -2422
rect 364404 -2742 364586 -2506
rect 364822 -2742 365004 -2506
rect 364404 -3684 365004 -2742
rect 368004 9654 368604 45098
rect 368004 9418 368186 9654
rect 368422 9418 368604 9654
rect 368004 9334 368604 9418
rect 368004 9098 368186 9334
rect 368422 9098 368604 9334
rect 368004 -4026 368604 9098
rect 368004 -4262 368186 -4026
rect 368422 -4262 368604 -4026
rect 368004 -4346 368604 -4262
rect 368004 -4582 368186 -4346
rect 368422 -4582 368604 -4346
rect 368004 -5524 368604 -4582
rect 371604 553254 372204 588698
rect 378804 705758 379404 705780
rect 378804 705522 378986 705758
rect 379222 705522 379404 705758
rect 378804 705438 379404 705522
rect 378804 705202 378986 705438
rect 379222 705202 379404 705438
rect 378804 668454 379404 705202
rect 378804 668218 378986 668454
rect 379222 668218 379404 668454
rect 378804 668134 379404 668218
rect 378804 667898 378986 668134
rect 379222 667898 379404 668134
rect 378804 632454 379404 667898
rect 378804 632218 378986 632454
rect 379222 632218 379404 632454
rect 378804 632134 379404 632218
rect 378804 631898 378986 632134
rect 379222 631898 379404 632134
rect 378804 596454 379404 631898
rect 378804 596218 378986 596454
rect 379222 596218 379404 596454
rect 378804 596134 379404 596218
rect 378804 595898 378986 596134
rect 379222 595898 379404 596134
rect 376707 560964 376773 560965
rect 376707 560900 376708 560964
rect 376772 560900 376773 560964
rect 376707 560899 376773 560900
rect 376710 560557 376770 560899
rect 376707 560556 376773 560557
rect 376707 560492 376708 560556
rect 376772 560492 376773 560556
rect 376707 560491 376773 560492
rect 371604 553018 371786 553254
rect 372022 553018 372204 553254
rect 371604 552934 372204 553018
rect 371604 552698 371786 552934
rect 372022 552698 372204 552934
rect 371604 517254 372204 552698
rect 371604 517018 371786 517254
rect 372022 517018 372204 517254
rect 371604 516934 372204 517018
rect 371604 516698 371786 516934
rect 372022 516698 372204 516934
rect 371604 481254 372204 516698
rect 371604 481018 371786 481254
rect 372022 481018 372204 481254
rect 371604 480934 372204 481018
rect 371604 480698 371786 480934
rect 372022 480698 372204 480934
rect 371604 445254 372204 480698
rect 371604 445018 371786 445254
rect 372022 445018 372204 445254
rect 371604 444934 372204 445018
rect 371604 444698 371786 444934
rect 372022 444698 372204 444934
rect 371604 409254 372204 444698
rect 371604 409018 371786 409254
rect 372022 409018 372204 409254
rect 371604 408934 372204 409018
rect 371604 408698 371786 408934
rect 372022 408698 372204 408934
rect 371604 373254 372204 408698
rect 371604 373018 371786 373254
rect 372022 373018 372204 373254
rect 371604 372934 372204 373018
rect 371604 372698 371786 372934
rect 372022 372698 372204 372934
rect 371604 337254 372204 372698
rect 371604 337018 371786 337254
rect 372022 337018 372204 337254
rect 371604 336934 372204 337018
rect 371604 336698 371786 336934
rect 372022 336698 372204 336934
rect 371604 301254 372204 336698
rect 371604 301018 371786 301254
rect 372022 301018 372204 301254
rect 371604 300934 372204 301018
rect 371604 300698 371786 300934
rect 372022 300698 372204 300934
rect 371604 265254 372204 300698
rect 371604 265018 371786 265254
rect 372022 265018 372204 265254
rect 371604 264934 372204 265018
rect 371604 264698 371786 264934
rect 372022 264698 372204 264934
rect 371604 229254 372204 264698
rect 371604 229018 371786 229254
rect 372022 229018 372204 229254
rect 371604 228934 372204 229018
rect 371604 228698 371786 228934
rect 372022 228698 372204 228934
rect 371604 193254 372204 228698
rect 371604 193018 371786 193254
rect 372022 193018 372204 193254
rect 371604 192934 372204 193018
rect 371604 192698 371786 192934
rect 372022 192698 372204 192934
rect 371604 157254 372204 192698
rect 371604 157018 371786 157254
rect 372022 157018 372204 157254
rect 371604 156934 372204 157018
rect 371604 156698 371786 156934
rect 372022 156698 372204 156934
rect 371604 121254 372204 156698
rect 371604 121018 371786 121254
rect 372022 121018 372204 121254
rect 371604 120934 372204 121018
rect 371604 120698 371786 120934
rect 372022 120698 372204 120934
rect 371604 85254 372204 120698
rect 371604 85018 371786 85254
rect 372022 85018 372204 85254
rect 371604 84934 372204 85018
rect 371604 84698 371786 84934
rect 372022 84698 372204 84934
rect 371604 49254 372204 84698
rect 371604 49018 371786 49254
rect 372022 49018 372204 49254
rect 371604 48934 372204 49018
rect 371604 48698 371786 48934
rect 372022 48698 372204 48934
rect 371604 13254 372204 48698
rect 371604 13018 371786 13254
rect 372022 13018 372204 13254
rect 371604 12934 372204 13018
rect 371604 12698 371786 12934
rect 372022 12698 372204 12934
rect 353604 -7022 353786 -6786
rect 354022 -7022 354204 -6786
rect 353604 -7106 354204 -7022
rect 353604 -7342 353786 -7106
rect 354022 -7342 354204 -7106
rect 353604 -7364 354204 -7342
rect 371604 -5866 372204 12698
rect 378804 560454 379404 595898
rect 378804 560218 378986 560454
rect 379222 560218 379404 560454
rect 378804 560134 379404 560218
rect 378804 559898 378986 560134
rect 379222 559898 379404 560134
rect 378804 524454 379404 559898
rect 378804 524218 378986 524454
rect 379222 524218 379404 524454
rect 378804 524134 379404 524218
rect 378804 523898 378986 524134
rect 379222 523898 379404 524134
rect 378804 488454 379404 523898
rect 378804 488218 378986 488454
rect 379222 488218 379404 488454
rect 378804 488134 379404 488218
rect 378804 487898 378986 488134
rect 379222 487898 379404 488134
rect 378804 452454 379404 487898
rect 378804 452218 378986 452454
rect 379222 452218 379404 452454
rect 378804 452134 379404 452218
rect 378804 451898 378986 452134
rect 379222 451898 379404 452134
rect 378804 416454 379404 451898
rect 378804 416218 378986 416454
rect 379222 416218 379404 416454
rect 378804 416134 379404 416218
rect 378804 415898 378986 416134
rect 379222 415898 379404 416134
rect 378804 380454 379404 415898
rect 378804 380218 378986 380454
rect 379222 380218 379404 380454
rect 378804 380134 379404 380218
rect 378804 379898 378986 380134
rect 379222 379898 379404 380134
rect 378804 344454 379404 379898
rect 378804 344218 378986 344454
rect 379222 344218 379404 344454
rect 378804 344134 379404 344218
rect 378804 343898 378986 344134
rect 379222 343898 379404 344134
rect 378804 308454 379404 343898
rect 378804 308218 378986 308454
rect 379222 308218 379404 308454
rect 378804 308134 379404 308218
rect 378804 307898 378986 308134
rect 379222 307898 379404 308134
rect 378804 272454 379404 307898
rect 378804 272218 378986 272454
rect 379222 272218 379404 272454
rect 378804 272134 379404 272218
rect 378804 271898 378986 272134
rect 379222 271898 379404 272134
rect 378804 236454 379404 271898
rect 378804 236218 378986 236454
rect 379222 236218 379404 236454
rect 378804 236134 379404 236218
rect 378804 235898 378986 236134
rect 379222 235898 379404 236134
rect 378804 200454 379404 235898
rect 378804 200218 378986 200454
rect 379222 200218 379404 200454
rect 378804 200134 379404 200218
rect 378804 199898 378986 200134
rect 379222 199898 379404 200134
rect 378804 164454 379404 199898
rect 378804 164218 378986 164454
rect 379222 164218 379404 164454
rect 378804 164134 379404 164218
rect 378804 163898 378986 164134
rect 379222 163898 379404 164134
rect 378804 128454 379404 163898
rect 378804 128218 378986 128454
rect 379222 128218 379404 128454
rect 378804 128134 379404 128218
rect 378804 127898 378986 128134
rect 379222 127898 379404 128134
rect 378804 92454 379404 127898
rect 378804 92218 378986 92454
rect 379222 92218 379404 92454
rect 378804 92134 379404 92218
rect 378804 91898 378986 92134
rect 379222 91898 379404 92134
rect 378804 56454 379404 91898
rect 378804 56218 378986 56454
rect 379222 56218 379404 56454
rect 378804 56134 379404 56218
rect 378804 55898 378986 56134
rect 379222 55898 379404 56134
rect 378804 20454 379404 55898
rect 378804 20218 378986 20454
rect 379222 20218 379404 20454
rect 378804 20134 379404 20218
rect 378804 19898 378986 20134
rect 379222 19898 379404 20134
rect 378804 -1266 379404 19898
rect 378804 -1502 378986 -1266
rect 379222 -1502 379404 -1266
rect 378804 -1586 379404 -1502
rect 378804 -1822 378986 -1586
rect 379222 -1822 379404 -1586
rect 378804 -1844 379404 -1822
rect 382404 672054 383004 707042
rect 382404 671818 382586 672054
rect 382822 671818 383004 672054
rect 382404 671734 383004 671818
rect 382404 671498 382586 671734
rect 382822 671498 383004 671734
rect 382404 636054 383004 671498
rect 382404 635818 382586 636054
rect 382822 635818 383004 636054
rect 382404 635734 383004 635818
rect 382404 635498 382586 635734
rect 382822 635498 383004 635734
rect 382404 600054 383004 635498
rect 382404 599818 382586 600054
rect 382822 599818 383004 600054
rect 382404 599734 383004 599818
rect 382404 599498 382586 599734
rect 382822 599498 383004 599734
rect 382404 564054 383004 599498
rect 382404 563818 382586 564054
rect 382822 563818 383004 564054
rect 382404 563734 383004 563818
rect 382404 563498 382586 563734
rect 382822 563498 383004 563734
rect 382404 528054 383004 563498
rect 386004 675654 386604 708882
rect 386004 675418 386186 675654
rect 386422 675418 386604 675654
rect 386004 675334 386604 675418
rect 386004 675098 386186 675334
rect 386422 675098 386604 675334
rect 386004 639654 386604 675098
rect 386004 639418 386186 639654
rect 386422 639418 386604 639654
rect 386004 639334 386604 639418
rect 386004 639098 386186 639334
rect 386422 639098 386604 639334
rect 386004 603654 386604 639098
rect 386004 603418 386186 603654
rect 386422 603418 386604 603654
rect 386004 603334 386604 603418
rect 386004 603098 386186 603334
rect 386422 603098 386604 603334
rect 386004 567654 386604 603098
rect 386004 567418 386186 567654
rect 386422 567418 386604 567654
rect 386004 567334 386604 567418
rect 386004 567098 386186 567334
rect 386422 567098 386604 567334
rect 384067 559468 384133 559469
rect 384067 559404 384068 559468
rect 384132 559404 384133 559468
rect 384067 559403 384133 559404
rect 383147 559332 383213 559333
rect 383147 559268 383148 559332
rect 383212 559268 383213 559332
rect 383147 559267 383213 559268
rect 383150 558245 383210 559267
rect 384070 559197 384130 559403
rect 384067 559196 384133 559197
rect 384067 559132 384068 559196
rect 384132 559132 384133 559196
rect 384067 559131 384133 559132
rect 383147 558244 383213 558245
rect 383147 558180 383148 558244
rect 383212 558180 383213 558244
rect 383147 558179 383213 558180
rect 382404 527818 382586 528054
rect 382822 527818 383004 528054
rect 382404 527734 383004 527818
rect 382404 527498 382586 527734
rect 382822 527498 383004 527734
rect 382404 492054 383004 527498
rect 382404 491818 382586 492054
rect 382822 491818 383004 492054
rect 382404 491734 383004 491818
rect 382404 491498 382586 491734
rect 382822 491498 383004 491734
rect 382404 456054 383004 491498
rect 382404 455818 382586 456054
rect 382822 455818 383004 456054
rect 382404 455734 383004 455818
rect 382404 455498 382586 455734
rect 382822 455498 383004 455734
rect 382404 420054 383004 455498
rect 382404 419818 382586 420054
rect 382822 419818 383004 420054
rect 382404 419734 383004 419818
rect 382404 419498 382586 419734
rect 382822 419498 383004 419734
rect 382404 384054 383004 419498
rect 382404 383818 382586 384054
rect 382822 383818 383004 384054
rect 382404 383734 383004 383818
rect 382404 383498 382586 383734
rect 382822 383498 383004 383734
rect 382404 348054 383004 383498
rect 382404 347818 382586 348054
rect 382822 347818 383004 348054
rect 382404 347734 383004 347818
rect 382404 347498 382586 347734
rect 382822 347498 383004 347734
rect 382404 312054 383004 347498
rect 382404 311818 382586 312054
rect 382822 311818 383004 312054
rect 382404 311734 383004 311818
rect 382404 311498 382586 311734
rect 382822 311498 383004 311734
rect 382404 276054 383004 311498
rect 382404 275818 382586 276054
rect 382822 275818 383004 276054
rect 382404 275734 383004 275818
rect 382404 275498 382586 275734
rect 382822 275498 383004 275734
rect 382404 240054 383004 275498
rect 382404 239818 382586 240054
rect 382822 239818 383004 240054
rect 382404 239734 383004 239818
rect 382404 239498 382586 239734
rect 382822 239498 383004 239734
rect 382404 204054 383004 239498
rect 382404 203818 382586 204054
rect 382822 203818 383004 204054
rect 382404 203734 383004 203818
rect 382404 203498 382586 203734
rect 382822 203498 383004 203734
rect 382404 168054 383004 203498
rect 382404 167818 382586 168054
rect 382822 167818 383004 168054
rect 382404 167734 383004 167818
rect 382404 167498 382586 167734
rect 382822 167498 383004 167734
rect 382404 132054 383004 167498
rect 382404 131818 382586 132054
rect 382822 131818 383004 132054
rect 382404 131734 383004 131818
rect 382404 131498 382586 131734
rect 382822 131498 383004 131734
rect 382404 96054 383004 131498
rect 382404 95818 382586 96054
rect 382822 95818 383004 96054
rect 382404 95734 383004 95818
rect 382404 95498 382586 95734
rect 382822 95498 383004 95734
rect 382404 60054 383004 95498
rect 382404 59818 382586 60054
rect 382822 59818 383004 60054
rect 382404 59734 383004 59818
rect 382404 59498 382586 59734
rect 382822 59498 383004 59734
rect 382404 24054 383004 59498
rect 382404 23818 382586 24054
rect 382822 23818 383004 24054
rect 382404 23734 383004 23818
rect 382404 23498 382586 23734
rect 382822 23498 383004 23734
rect 382404 -3106 383004 23498
rect 382404 -3342 382586 -3106
rect 382822 -3342 383004 -3106
rect 382404 -3426 383004 -3342
rect 382404 -3662 382586 -3426
rect 382822 -3662 383004 -3426
rect 382404 -3684 383004 -3662
rect 386004 531654 386604 567098
rect 386004 531418 386186 531654
rect 386422 531418 386604 531654
rect 386004 531334 386604 531418
rect 386004 531098 386186 531334
rect 386422 531098 386604 531334
rect 386004 495654 386604 531098
rect 386004 495418 386186 495654
rect 386422 495418 386604 495654
rect 386004 495334 386604 495418
rect 386004 495098 386186 495334
rect 386422 495098 386604 495334
rect 386004 459654 386604 495098
rect 386004 459418 386186 459654
rect 386422 459418 386604 459654
rect 386004 459334 386604 459418
rect 386004 459098 386186 459334
rect 386422 459098 386604 459334
rect 386004 423654 386604 459098
rect 386004 423418 386186 423654
rect 386422 423418 386604 423654
rect 386004 423334 386604 423418
rect 386004 423098 386186 423334
rect 386422 423098 386604 423334
rect 386004 387654 386604 423098
rect 386004 387418 386186 387654
rect 386422 387418 386604 387654
rect 386004 387334 386604 387418
rect 386004 387098 386186 387334
rect 386422 387098 386604 387334
rect 386004 351654 386604 387098
rect 386004 351418 386186 351654
rect 386422 351418 386604 351654
rect 386004 351334 386604 351418
rect 386004 351098 386186 351334
rect 386422 351098 386604 351334
rect 386004 315654 386604 351098
rect 386004 315418 386186 315654
rect 386422 315418 386604 315654
rect 386004 315334 386604 315418
rect 386004 315098 386186 315334
rect 386422 315098 386604 315334
rect 386004 279654 386604 315098
rect 386004 279418 386186 279654
rect 386422 279418 386604 279654
rect 386004 279334 386604 279418
rect 386004 279098 386186 279334
rect 386422 279098 386604 279334
rect 386004 243654 386604 279098
rect 386004 243418 386186 243654
rect 386422 243418 386604 243654
rect 386004 243334 386604 243418
rect 386004 243098 386186 243334
rect 386422 243098 386604 243334
rect 386004 207654 386604 243098
rect 386004 207418 386186 207654
rect 386422 207418 386604 207654
rect 386004 207334 386604 207418
rect 386004 207098 386186 207334
rect 386422 207098 386604 207334
rect 386004 171654 386604 207098
rect 386004 171418 386186 171654
rect 386422 171418 386604 171654
rect 386004 171334 386604 171418
rect 386004 171098 386186 171334
rect 386422 171098 386604 171334
rect 386004 135654 386604 171098
rect 386004 135418 386186 135654
rect 386422 135418 386604 135654
rect 386004 135334 386604 135418
rect 386004 135098 386186 135334
rect 386422 135098 386604 135334
rect 386004 99654 386604 135098
rect 386004 99418 386186 99654
rect 386422 99418 386604 99654
rect 386004 99334 386604 99418
rect 386004 99098 386186 99334
rect 386422 99098 386604 99334
rect 386004 63654 386604 99098
rect 386004 63418 386186 63654
rect 386422 63418 386604 63654
rect 386004 63334 386604 63418
rect 386004 63098 386186 63334
rect 386422 63098 386604 63334
rect 386004 27654 386604 63098
rect 386004 27418 386186 27654
rect 386422 27418 386604 27654
rect 386004 27334 386604 27418
rect 386004 27098 386186 27334
rect 386422 27098 386604 27334
rect 386004 -4946 386604 27098
rect 386004 -5182 386186 -4946
rect 386422 -5182 386604 -4946
rect 386004 -5266 386604 -5182
rect 386004 -5502 386186 -5266
rect 386422 -5502 386604 -5266
rect 386004 -5524 386604 -5502
rect 389604 679254 390204 710722
rect 407604 710358 408204 711300
rect 407604 710122 407786 710358
rect 408022 710122 408204 710358
rect 407604 710038 408204 710122
rect 407604 709802 407786 710038
rect 408022 709802 408204 710038
rect 404004 708518 404604 709460
rect 404004 708282 404186 708518
rect 404422 708282 404604 708518
rect 404004 708198 404604 708282
rect 404004 707962 404186 708198
rect 404422 707962 404604 708198
rect 400404 706678 401004 707620
rect 400404 706442 400586 706678
rect 400822 706442 401004 706678
rect 400404 706358 401004 706442
rect 400404 706122 400586 706358
rect 400822 706122 401004 706358
rect 389604 679018 389786 679254
rect 390022 679018 390204 679254
rect 389604 678934 390204 679018
rect 389604 678698 389786 678934
rect 390022 678698 390204 678934
rect 389604 643254 390204 678698
rect 389604 643018 389786 643254
rect 390022 643018 390204 643254
rect 389604 642934 390204 643018
rect 389604 642698 389786 642934
rect 390022 642698 390204 642934
rect 389604 607254 390204 642698
rect 389604 607018 389786 607254
rect 390022 607018 390204 607254
rect 389604 606934 390204 607018
rect 389604 606698 389786 606934
rect 390022 606698 390204 606934
rect 389604 571254 390204 606698
rect 389604 571018 389786 571254
rect 390022 571018 390204 571254
rect 389604 570934 390204 571018
rect 389604 570698 389786 570934
rect 390022 570698 390204 570934
rect 389604 535254 390204 570698
rect 396804 704838 397404 705780
rect 396804 704602 396986 704838
rect 397222 704602 397404 704838
rect 396804 704518 397404 704602
rect 396804 704282 396986 704518
rect 397222 704282 397404 704518
rect 396804 686454 397404 704282
rect 396804 686218 396986 686454
rect 397222 686218 397404 686454
rect 396804 686134 397404 686218
rect 396804 685898 396986 686134
rect 397222 685898 397404 686134
rect 396804 650454 397404 685898
rect 396804 650218 396986 650454
rect 397222 650218 397404 650454
rect 396804 650134 397404 650218
rect 396804 649898 396986 650134
rect 397222 649898 397404 650134
rect 396804 614454 397404 649898
rect 396804 614218 396986 614454
rect 397222 614218 397404 614454
rect 396804 614134 397404 614218
rect 396804 613898 396986 614134
rect 397222 613898 397404 614134
rect 396804 578454 397404 613898
rect 396804 578218 396986 578454
rect 397222 578218 397404 578454
rect 396804 578134 397404 578218
rect 396804 577898 396986 578134
rect 397222 577898 397404 578134
rect 393270 561373 393330 562582
rect 393267 561372 393333 561373
rect 393267 561308 393268 561372
rect 393332 561308 393333 561372
rect 393267 561307 393333 561308
rect 396027 559332 396093 559333
rect 396027 559268 396028 559332
rect 396092 559268 396093 559332
rect 396027 559267 396093 559268
rect 396030 559061 396090 559267
rect 396027 559060 396093 559061
rect 396027 558996 396028 559060
rect 396092 558996 396093 559060
rect 396027 558995 396093 558996
rect 389604 535018 389786 535254
rect 390022 535018 390204 535254
rect 389604 534934 390204 535018
rect 389604 534698 389786 534934
rect 390022 534698 390204 534934
rect 389604 499254 390204 534698
rect 389604 499018 389786 499254
rect 390022 499018 390204 499254
rect 389604 498934 390204 499018
rect 389604 498698 389786 498934
rect 390022 498698 390204 498934
rect 389604 463254 390204 498698
rect 389604 463018 389786 463254
rect 390022 463018 390204 463254
rect 389604 462934 390204 463018
rect 389604 462698 389786 462934
rect 390022 462698 390204 462934
rect 389604 427254 390204 462698
rect 389604 427018 389786 427254
rect 390022 427018 390204 427254
rect 389604 426934 390204 427018
rect 389604 426698 389786 426934
rect 390022 426698 390204 426934
rect 389604 391254 390204 426698
rect 389604 391018 389786 391254
rect 390022 391018 390204 391254
rect 389604 390934 390204 391018
rect 389604 390698 389786 390934
rect 390022 390698 390204 390934
rect 389604 355254 390204 390698
rect 389604 355018 389786 355254
rect 390022 355018 390204 355254
rect 389604 354934 390204 355018
rect 389604 354698 389786 354934
rect 390022 354698 390204 354934
rect 389604 319254 390204 354698
rect 389604 319018 389786 319254
rect 390022 319018 390204 319254
rect 389604 318934 390204 319018
rect 389604 318698 389786 318934
rect 390022 318698 390204 318934
rect 389604 283254 390204 318698
rect 389604 283018 389786 283254
rect 390022 283018 390204 283254
rect 389604 282934 390204 283018
rect 389604 282698 389786 282934
rect 390022 282698 390204 282934
rect 389604 247254 390204 282698
rect 389604 247018 389786 247254
rect 390022 247018 390204 247254
rect 389604 246934 390204 247018
rect 389604 246698 389786 246934
rect 390022 246698 390204 246934
rect 389604 211254 390204 246698
rect 389604 211018 389786 211254
rect 390022 211018 390204 211254
rect 389604 210934 390204 211018
rect 389604 210698 389786 210934
rect 390022 210698 390204 210934
rect 389604 175254 390204 210698
rect 389604 175018 389786 175254
rect 390022 175018 390204 175254
rect 389604 174934 390204 175018
rect 389604 174698 389786 174934
rect 390022 174698 390204 174934
rect 389604 139254 390204 174698
rect 389604 139018 389786 139254
rect 390022 139018 390204 139254
rect 389604 138934 390204 139018
rect 389604 138698 389786 138934
rect 390022 138698 390204 138934
rect 389604 103254 390204 138698
rect 389604 103018 389786 103254
rect 390022 103018 390204 103254
rect 389604 102934 390204 103018
rect 389604 102698 389786 102934
rect 390022 102698 390204 102934
rect 389604 67254 390204 102698
rect 389604 67018 389786 67254
rect 390022 67018 390204 67254
rect 389604 66934 390204 67018
rect 389604 66698 389786 66934
rect 390022 66698 390204 66934
rect 389604 31254 390204 66698
rect 389604 31018 389786 31254
rect 390022 31018 390204 31254
rect 389604 30934 390204 31018
rect 389604 30698 389786 30934
rect 390022 30698 390204 30934
rect 371604 -6102 371786 -5866
rect 372022 -6102 372204 -5866
rect 371604 -6186 372204 -6102
rect 371604 -6422 371786 -6186
rect 372022 -6422 372204 -6186
rect 371604 -7364 372204 -6422
rect 389604 -6786 390204 30698
rect 396804 542454 397404 577898
rect 396804 542218 396986 542454
rect 397222 542218 397404 542454
rect 396804 542134 397404 542218
rect 396804 541898 396986 542134
rect 397222 541898 397404 542134
rect 396804 506454 397404 541898
rect 396804 506218 396986 506454
rect 397222 506218 397404 506454
rect 396804 506134 397404 506218
rect 396804 505898 396986 506134
rect 397222 505898 397404 506134
rect 396804 470454 397404 505898
rect 396804 470218 396986 470454
rect 397222 470218 397404 470454
rect 396804 470134 397404 470218
rect 396804 469898 396986 470134
rect 397222 469898 397404 470134
rect 396804 434454 397404 469898
rect 396804 434218 396986 434454
rect 397222 434218 397404 434454
rect 396804 434134 397404 434218
rect 396804 433898 396986 434134
rect 397222 433898 397404 434134
rect 396804 398454 397404 433898
rect 396804 398218 396986 398454
rect 397222 398218 397404 398454
rect 396804 398134 397404 398218
rect 396804 397898 396986 398134
rect 397222 397898 397404 398134
rect 396804 362454 397404 397898
rect 396804 362218 396986 362454
rect 397222 362218 397404 362454
rect 396804 362134 397404 362218
rect 396804 361898 396986 362134
rect 397222 361898 397404 362134
rect 396804 326454 397404 361898
rect 396804 326218 396986 326454
rect 397222 326218 397404 326454
rect 396804 326134 397404 326218
rect 396804 325898 396986 326134
rect 397222 325898 397404 326134
rect 396804 290454 397404 325898
rect 396804 290218 396986 290454
rect 397222 290218 397404 290454
rect 396804 290134 397404 290218
rect 396804 289898 396986 290134
rect 397222 289898 397404 290134
rect 396804 254454 397404 289898
rect 396804 254218 396986 254454
rect 397222 254218 397404 254454
rect 396804 254134 397404 254218
rect 396804 253898 396986 254134
rect 397222 253898 397404 254134
rect 396804 218454 397404 253898
rect 396804 218218 396986 218454
rect 397222 218218 397404 218454
rect 396804 218134 397404 218218
rect 396804 217898 396986 218134
rect 397222 217898 397404 218134
rect 396804 182454 397404 217898
rect 396804 182218 396986 182454
rect 397222 182218 397404 182454
rect 396804 182134 397404 182218
rect 396804 181898 396986 182134
rect 397222 181898 397404 182134
rect 396804 146454 397404 181898
rect 396804 146218 396986 146454
rect 397222 146218 397404 146454
rect 396804 146134 397404 146218
rect 396804 145898 396986 146134
rect 397222 145898 397404 146134
rect 396804 110454 397404 145898
rect 396804 110218 396986 110454
rect 397222 110218 397404 110454
rect 396804 110134 397404 110218
rect 396804 109898 396986 110134
rect 397222 109898 397404 110134
rect 396804 74454 397404 109898
rect 396804 74218 396986 74454
rect 397222 74218 397404 74454
rect 396804 74134 397404 74218
rect 396804 73898 396986 74134
rect 397222 73898 397404 74134
rect 396804 38454 397404 73898
rect 396804 38218 396986 38454
rect 397222 38218 397404 38454
rect 396804 38134 397404 38218
rect 396804 37898 396986 38134
rect 397222 37898 397404 38134
rect 396804 2454 397404 37898
rect 396804 2218 396986 2454
rect 397222 2218 397404 2454
rect 396804 2134 397404 2218
rect 396804 1898 396986 2134
rect 397222 1898 397404 2134
rect 396804 -346 397404 1898
rect 396804 -582 396986 -346
rect 397222 -582 397404 -346
rect 396804 -666 397404 -582
rect 396804 -902 396986 -666
rect 397222 -902 397404 -666
rect 396804 -1844 397404 -902
rect 400404 690054 401004 706122
rect 400404 689818 400586 690054
rect 400822 689818 401004 690054
rect 400404 689734 401004 689818
rect 400404 689498 400586 689734
rect 400822 689498 401004 689734
rect 400404 654054 401004 689498
rect 400404 653818 400586 654054
rect 400822 653818 401004 654054
rect 400404 653734 401004 653818
rect 400404 653498 400586 653734
rect 400822 653498 401004 653734
rect 400404 618054 401004 653498
rect 400404 617818 400586 618054
rect 400822 617818 401004 618054
rect 400404 617734 401004 617818
rect 400404 617498 400586 617734
rect 400822 617498 401004 617734
rect 400404 582054 401004 617498
rect 400404 581818 400586 582054
rect 400822 581818 401004 582054
rect 400404 581734 401004 581818
rect 400404 581498 400586 581734
rect 400822 581498 401004 581734
rect 400404 546054 401004 581498
rect 400404 545818 400586 546054
rect 400822 545818 401004 546054
rect 400404 545734 401004 545818
rect 400404 545498 400586 545734
rect 400822 545498 401004 545734
rect 400404 510054 401004 545498
rect 400404 509818 400586 510054
rect 400822 509818 401004 510054
rect 400404 509734 401004 509818
rect 400404 509498 400586 509734
rect 400822 509498 401004 509734
rect 400404 474054 401004 509498
rect 400404 473818 400586 474054
rect 400822 473818 401004 474054
rect 400404 473734 401004 473818
rect 400404 473498 400586 473734
rect 400822 473498 401004 473734
rect 400404 438054 401004 473498
rect 400404 437818 400586 438054
rect 400822 437818 401004 438054
rect 400404 437734 401004 437818
rect 400404 437498 400586 437734
rect 400822 437498 401004 437734
rect 400404 402054 401004 437498
rect 400404 401818 400586 402054
rect 400822 401818 401004 402054
rect 400404 401734 401004 401818
rect 400404 401498 400586 401734
rect 400822 401498 401004 401734
rect 400404 366054 401004 401498
rect 400404 365818 400586 366054
rect 400822 365818 401004 366054
rect 400404 365734 401004 365818
rect 400404 365498 400586 365734
rect 400822 365498 401004 365734
rect 400404 330054 401004 365498
rect 400404 329818 400586 330054
rect 400822 329818 401004 330054
rect 400404 329734 401004 329818
rect 400404 329498 400586 329734
rect 400822 329498 401004 329734
rect 400404 294054 401004 329498
rect 400404 293818 400586 294054
rect 400822 293818 401004 294054
rect 400404 293734 401004 293818
rect 400404 293498 400586 293734
rect 400822 293498 401004 293734
rect 400404 258054 401004 293498
rect 400404 257818 400586 258054
rect 400822 257818 401004 258054
rect 400404 257734 401004 257818
rect 400404 257498 400586 257734
rect 400822 257498 401004 257734
rect 400404 222054 401004 257498
rect 400404 221818 400586 222054
rect 400822 221818 401004 222054
rect 400404 221734 401004 221818
rect 400404 221498 400586 221734
rect 400822 221498 401004 221734
rect 400404 186054 401004 221498
rect 400404 185818 400586 186054
rect 400822 185818 401004 186054
rect 400404 185734 401004 185818
rect 400404 185498 400586 185734
rect 400822 185498 401004 185734
rect 400404 150054 401004 185498
rect 400404 149818 400586 150054
rect 400822 149818 401004 150054
rect 400404 149734 401004 149818
rect 400404 149498 400586 149734
rect 400822 149498 401004 149734
rect 400404 114054 401004 149498
rect 400404 113818 400586 114054
rect 400822 113818 401004 114054
rect 400404 113734 401004 113818
rect 400404 113498 400586 113734
rect 400822 113498 401004 113734
rect 400404 78054 401004 113498
rect 400404 77818 400586 78054
rect 400822 77818 401004 78054
rect 400404 77734 401004 77818
rect 400404 77498 400586 77734
rect 400822 77498 401004 77734
rect 400404 42054 401004 77498
rect 400404 41818 400586 42054
rect 400822 41818 401004 42054
rect 400404 41734 401004 41818
rect 400404 41498 400586 41734
rect 400822 41498 401004 41734
rect 400404 6054 401004 41498
rect 400404 5818 400586 6054
rect 400822 5818 401004 6054
rect 400404 5734 401004 5818
rect 400404 5498 400586 5734
rect 400822 5498 401004 5734
rect 400404 -2186 401004 5498
rect 400404 -2422 400586 -2186
rect 400822 -2422 401004 -2186
rect 400404 -2506 401004 -2422
rect 400404 -2742 400586 -2506
rect 400822 -2742 401004 -2506
rect 400404 -3684 401004 -2742
rect 404004 693654 404604 707962
rect 404004 693418 404186 693654
rect 404422 693418 404604 693654
rect 404004 693334 404604 693418
rect 404004 693098 404186 693334
rect 404422 693098 404604 693334
rect 404004 657654 404604 693098
rect 404004 657418 404186 657654
rect 404422 657418 404604 657654
rect 404004 657334 404604 657418
rect 404004 657098 404186 657334
rect 404422 657098 404604 657334
rect 404004 621654 404604 657098
rect 404004 621418 404186 621654
rect 404422 621418 404604 621654
rect 404004 621334 404604 621418
rect 404004 621098 404186 621334
rect 404422 621098 404604 621334
rect 404004 585654 404604 621098
rect 404004 585418 404186 585654
rect 404422 585418 404604 585654
rect 404004 585334 404604 585418
rect 404004 585098 404186 585334
rect 404422 585098 404604 585334
rect 404004 549654 404604 585098
rect 407604 697254 408204 709802
rect 425604 711278 426204 711300
rect 425604 711042 425786 711278
rect 426022 711042 426204 711278
rect 425604 710958 426204 711042
rect 425604 710722 425786 710958
rect 426022 710722 426204 710958
rect 422004 709438 422604 709460
rect 422004 709202 422186 709438
rect 422422 709202 422604 709438
rect 422004 709118 422604 709202
rect 422004 708882 422186 709118
rect 422422 708882 422604 709118
rect 418404 707598 419004 707620
rect 418404 707362 418586 707598
rect 418822 707362 419004 707598
rect 418404 707278 419004 707362
rect 418404 707042 418586 707278
rect 418822 707042 419004 707278
rect 407604 697018 407786 697254
rect 408022 697018 408204 697254
rect 407604 696934 408204 697018
rect 407604 696698 407786 696934
rect 408022 696698 408204 696934
rect 407604 661254 408204 696698
rect 407604 661018 407786 661254
rect 408022 661018 408204 661254
rect 407604 660934 408204 661018
rect 407604 660698 407786 660934
rect 408022 660698 408204 660934
rect 407604 625254 408204 660698
rect 407604 625018 407786 625254
rect 408022 625018 408204 625254
rect 407604 624934 408204 625018
rect 407604 624698 407786 624934
rect 408022 624698 408204 624934
rect 407604 589254 408204 624698
rect 407604 589018 407786 589254
rect 408022 589018 408204 589254
rect 407604 588934 408204 589018
rect 407604 588698 407786 588934
rect 408022 588698 408204 588934
rect 406334 561373 406394 561902
rect 406331 561372 406397 561373
rect 406331 561308 406332 561372
rect 406396 561308 406397 561372
rect 406331 561307 406397 561308
rect 404004 549418 404186 549654
rect 404422 549418 404604 549654
rect 404004 549334 404604 549418
rect 404004 549098 404186 549334
rect 404422 549098 404604 549334
rect 404004 513654 404604 549098
rect 404004 513418 404186 513654
rect 404422 513418 404604 513654
rect 404004 513334 404604 513418
rect 404004 513098 404186 513334
rect 404422 513098 404604 513334
rect 404004 477654 404604 513098
rect 404004 477418 404186 477654
rect 404422 477418 404604 477654
rect 404004 477334 404604 477418
rect 404004 477098 404186 477334
rect 404422 477098 404604 477334
rect 404004 441654 404604 477098
rect 404004 441418 404186 441654
rect 404422 441418 404604 441654
rect 404004 441334 404604 441418
rect 404004 441098 404186 441334
rect 404422 441098 404604 441334
rect 404004 405654 404604 441098
rect 404004 405418 404186 405654
rect 404422 405418 404604 405654
rect 404004 405334 404604 405418
rect 404004 405098 404186 405334
rect 404422 405098 404604 405334
rect 404004 369654 404604 405098
rect 404004 369418 404186 369654
rect 404422 369418 404604 369654
rect 404004 369334 404604 369418
rect 404004 369098 404186 369334
rect 404422 369098 404604 369334
rect 404004 333654 404604 369098
rect 404004 333418 404186 333654
rect 404422 333418 404604 333654
rect 404004 333334 404604 333418
rect 404004 333098 404186 333334
rect 404422 333098 404604 333334
rect 404004 297654 404604 333098
rect 404004 297418 404186 297654
rect 404422 297418 404604 297654
rect 404004 297334 404604 297418
rect 404004 297098 404186 297334
rect 404422 297098 404604 297334
rect 404004 261654 404604 297098
rect 404004 261418 404186 261654
rect 404422 261418 404604 261654
rect 404004 261334 404604 261418
rect 404004 261098 404186 261334
rect 404422 261098 404604 261334
rect 404004 225654 404604 261098
rect 404004 225418 404186 225654
rect 404422 225418 404604 225654
rect 404004 225334 404604 225418
rect 404004 225098 404186 225334
rect 404422 225098 404604 225334
rect 404004 189654 404604 225098
rect 404004 189418 404186 189654
rect 404422 189418 404604 189654
rect 404004 189334 404604 189418
rect 404004 189098 404186 189334
rect 404422 189098 404604 189334
rect 404004 153654 404604 189098
rect 404004 153418 404186 153654
rect 404422 153418 404604 153654
rect 404004 153334 404604 153418
rect 404004 153098 404186 153334
rect 404422 153098 404604 153334
rect 404004 117654 404604 153098
rect 404004 117418 404186 117654
rect 404422 117418 404604 117654
rect 404004 117334 404604 117418
rect 404004 117098 404186 117334
rect 404422 117098 404604 117334
rect 404004 81654 404604 117098
rect 404004 81418 404186 81654
rect 404422 81418 404604 81654
rect 404004 81334 404604 81418
rect 404004 81098 404186 81334
rect 404422 81098 404604 81334
rect 404004 45654 404604 81098
rect 404004 45418 404186 45654
rect 404422 45418 404604 45654
rect 404004 45334 404604 45418
rect 404004 45098 404186 45334
rect 404422 45098 404604 45334
rect 404004 9654 404604 45098
rect 404004 9418 404186 9654
rect 404422 9418 404604 9654
rect 404004 9334 404604 9418
rect 404004 9098 404186 9334
rect 404422 9098 404604 9334
rect 404004 -4026 404604 9098
rect 404004 -4262 404186 -4026
rect 404422 -4262 404604 -4026
rect 404004 -4346 404604 -4262
rect 404004 -4582 404186 -4346
rect 404422 -4582 404604 -4346
rect 404004 -5524 404604 -4582
rect 407604 553254 408204 588698
rect 414804 705758 415404 705780
rect 414804 705522 414986 705758
rect 415222 705522 415404 705758
rect 414804 705438 415404 705522
rect 414804 705202 414986 705438
rect 415222 705202 415404 705438
rect 414804 668454 415404 705202
rect 414804 668218 414986 668454
rect 415222 668218 415404 668454
rect 414804 668134 415404 668218
rect 414804 667898 414986 668134
rect 415222 667898 415404 668134
rect 414804 632454 415404 667898
rect 414804 632218 414986 632454
rect 415222 632218 415404 632454
rect 414804 632134 415404 632218
rect 414804 631898 414986 632134
rect 415222 631898 415404 632134
rect 414804 596454 415404 631898
rect 414804 596218 414986 596454
rect 415222 596218 415404 596454
rect 414804 596134 415404 596218
rect 414804 595898 414986 596134
rect 415222 595898 415404 596134
rect 414804 560454 415404 595898
rect 414804 560218 414986 560454
rect 415222 560218 415404 560454
rect 414804 560134 415404 560218
rect 414804 559898 414986 560134
rect 415222 559898 415404 560134
rect 409091 559468 409157 559469
rect 409091 559404 409092 559468
rect 409156 559404 409157 559468
rect 409091 559403 409157 559404
rect 409094 559061 409154 559403
rect 409091 559060 409157 559061
rect 409091 558996 409092 559060
rect 409156 558996 409157 559060
rect 409091 558995 409157 558996
rect 407604 553018 407786 553254
rect 408022 553018 408204 553254
rect 407604 552934 408204 553018
rect 407604 552698 407786 552934
rect 408022 552698 408204 552934
rect 407604 517254 408204 552698
rect 407604 517018 407786 517254
rect 408022 517018 408204 517254
rect 407604 516934 408204 517018
rect 407604 516698 407786 516934
rect 408022 516698 408204 516934
rect 407604 481254 408204 516698
rect 407604 481018 407786 481254
rect 408022 481018 408204 481254
rect 407604 480934 408204 481018
rect 407604 480698 407786 480934
rect 408022 480698 408204 480934
rect 407604 445254 408204 480698
rect 407604 445018 407786 445254
rect 408022 445018 408204 445254
rect 407604 444934 408204 445018
rect 407604 444698 407786 444934
rect 408022 444698 408204 444934
rect 407604 409254 408204 444698
rect 407604 409018 407786 409254
rect 408022 409018 408204 409254
rect 407604 408934 408204 409018
rect 407604 408698 407786 408934
rect 408022 408698 408204 408934
rect 407604 373254 408204 408698
rect 407604 373018 407786 373254
rect 408022 373018 408204 373254
rect 407604 372934 408204 373018
rect 407604 372698 407786 372934
rect 408022 372698 408204 372934
rect 407604 337254 408204 372698
rect 407604 337018 407786 337254
rect 408022 337018 408204 337254
rect 407604 336934 408204 337018
rect 407604 336698 407786 336934
rect 408022 336698 408204 336934
rect 407604 301254 408204 336698
rect 407604 301018 407786 301254
rect 408022 301018 408204 301254
rect 407604 300934 408204 301018
rect 407604 300698 407786 300934
rect 408022 300698 408204 300934
rect 407604 265254 408204 300698
rect 407604 265018 407786 265254
rect 408022 265018 408204 265254
rect 407604 264934 408204 265018
rect 407604 264698 407786 264934
rect 408022 264698 408204 264934
rect 407604 229254 408204 264698
rect 407604 229018 407786 229254
rect 408022 229018 408204 229254
rect 407604 228934 408204 229018
rect 407604 228698 407786 228934
rect 408022 228698 408204 228934
rect 407604 193254 408204 228698
rect 407604 193018 407786 193254
rect 408022 193018 408204 193254
rect 407604 192934 408204 193018
rect 407604 192698 407786 192934
rect 408022 192698 408204 192934
rect 407604 157254 408204 192698
rect 407604 157018 407786 157254
rect 408022 157018 408204 157254
rect 407604 156934 408204 157018
rect 407604 156698 407786 156934
rect 408022 156698 408204 156934
rect 407604 121254 408204 156698
rect 407604 121018 407786 121254
rect 408022 121018 408204 121254
rect 407604 120934 408204 121018
rect 407604 120698 407786 120934
rect 408022 120698 408204 120934
rect 407604 85254 408204 120698
rect 407604 85018 407786 85254
rect 408022 85018 408204 85254
rect 407604 84934 408204 85018
rect 407604 84698 407786 84934
rect 408022 84698 408204 84934
rect 407604 49254 408204 84698
rect 407604 49018 407786 49254
rect 408022 49018 408204 49254
rect 407604 48934 408204 49018
rect 407604 48698 407786 48934
rect 408022 48698 408204 48934
rect 407604 13254 408204 48698
rect 407604 13018 407786 13254
rect 408022 13018 408204 13254
rect 407604 12934 408204 13018
rect 407604 12698 407786 12934
rect 408022 12698 408204 12934
rect 389604 -7022 389786 -6786
rect 390022 -7022 390204 -6786
rect 389604 -7106 390204 -7022
rect 389604 -7342 389786 -7106
rect 390022 -7342 390204 -7106
rect 389604 -7364 390204 -7342
rect 407604 -5866 408204 12698
rect 414804 524454 415404 559898
rect 414804 524218 414986 524454
rect 415222 524218 415404 524454
rect 414804 524134 415404 524218
rect 414804 523898 414986 524134
rect 415222 523898 415404 524134
rect 414804 488454 415404 523898
rect 414804 488218 414986 488454
rect 415222 488218 415404 488454
rect 414804 488134 415404 488218
rect 414804 487898 414986 488134
rect 415222 487898 415404 488134
rect 414804 452454 415404 487898
rect 414804 452218 414986 452454
rect 415222 452218 415404 452454
rect 414804 452134 415404 452218
rect 414804 451898 414986 452134
rect 415222 451898 415404 452134
rect 414804 416454 415404 451898
rect 414804 416218 414986 416454
rect 415222 416218 415404 416454
rect 414804 416134 415404 416218
rect 414804 415898 414986 416134
rect 415222 415898 415404 416134
rect 414804 380454 415404 415898
rect 414804 380218 414986 380454
rect 415222 380218 415404 380454
rect 414804 380134 415404 380218
rect 414804 379898 414986 380134
rect 415222 379898 415404 380134
rect 414804 344454 415404 379898
rect 414804 344218 414986 344454
rect 415222 344218 415404 344454
rect 414804 344134 415404 344218
rect 414804 343898 414986 344134
rect 415222 343898 415404 344134
rect 414804 308454 415404 343898
rect 414804 308218 414986 308454
rect 415222 308218 415404 308454
rect 414804 308134 415404 308218
rect 414804 307898 414986 308134
rect 415222 307898 415404 308134
rect 414804 272454 415404 307898
rect 414804 272218 414986 272454
rect 415222 272218 415404 272454
rect 414804 272134 415404 272218
rect 414804 271898 414986 272134
rect 415222 271898 415404 272134
rect 414804 236454 415404 271898
rect 414804 236218 414986 236454
rect 415222 236218 415404 236454
rect 414804 236134 415404 236218
rect 414804 235898 414986 236134
rect 415222 235898 415404 236134
rect 414804 200454 415404 235898
rect 414804 200218 414986 200454
rect 415222 200218 415404 200454
rect 414804 200134 415404 200218
rect 414804 199898 414986 200134
rect 415222 199898 415404 200134
rect 414804 164454 415404 199898
rect 414804 164218 414986 164454
rect 415222 164218 415404 164454
rect 414804 164134 415404 164218
rect 414804 163898 414986 164134
rect 415222 163898 415404 164134
rect 414804 128454 415404 163898
rect 414804 128218 414986 128454
rect 415222 128218 415404 128454
rect 414804 128134 415404 128218
rect 414804 127898 414986 128134
rect 415222 127898 415404 128134
rect 414804 92454 415404 127898
rect 414804 92218 414986 92454
rect 415222 92218 415404 92454
rect 414804 92134 415404 92218
rect 414804 91898 414986 92134
rect 415222 91898 415404 92134
rect 414804 56454 415404 91898
rect 414804 56218 414986 56454
rect 415222 56218 415404 56454
rect 414804 56134 415404 56218
rect 414804 55898 414986 56134
rect 415222 55898 415404 56134
rect 414804 20454 415404 55898
rect 414804 20218 414986 20454
rect 415222 20218 415404 20454
rect 414804 20134 415404 20218
rect 414804 19898 414986 20134
rect 415222 19898 415404 20134
rect 414804 -1266 415404 19898
rect 414804 -1502 414986 -1266
rect 415222 -1502 415404 -1266
rect 414804 -1586 415404 -1502
rect 414804 -1822 414986 -1586
rect 415222 -1822 415404 -1586
rect 414804 -1844 415404 -1822
rect 418404 672054 419004 707042
rect 418404 671818 418586 672054
rect 418822 671818 419004 672054
rect 418404 671734 419004 671818
rect 418404 671498 418586 671734
rect 418822 671498 419004 671734
rect 418404 636054 419004 671498
rect 418404 635818 418586 636054
rect 418822 635818 419004 636054
rect 418404 635734 419004 635818
rect 418404 635498 418586 635734
rect 418822 635498 419004 635734
rect 418404 600054 419004 635498
rect 418404 599818 418586 600054
rect 418822 599818 419004 600054
rect 418404 599734 419004 599818
rect 418404 599498 418586 599734
rect 418822 599498 419004 599734
rect 418404 564054 419004 599498
rect 418404 563818 418586 564054
rect 418822 563818 419004 564054
rect 418404 563734 419004 563818
rect 418404 563498 418586 563734
rect 418822 563498 419004 563734
rect 418404 528054 419004 563498
rect 418404 527818 418586 528054
rect 418822 527818 419004 528054
rect 418404 527734 419004 527818
rect 418404 527498 418586 527734
rect 418822 527498 419004 527734
rect 418404 492054 419004 527498
rect 418404 491818 418586 492054
rect 418822 491818 419004 492054
rect 418404 491734 419004 491818
rect 418404 491498 418586 491734
rect 418822 491498 419004 491734
rect 418404 456054 419004 491498
rect 418404 455818 418586 456054
rect 418822 455818 419004 456054
rect 418404 455734 419004 455818
rect 418404 455498 418586 455734
rect 418822 455498 419004 455734
rect 418404 420054 419004 455498
rect 418404 419818 418586 420054
rect 418822 419818 419004 420054
rect 418404 419734 419004 419818
rect 418404 419498 418586 419734
rect 418822 419498 419004 419734
rect 418404 384054 419004 419498
rect 418404 383818 418586 384054
rect 418822 383818 419004 384054
rect 418404 383734 419004 383818
rect 418404 383498 418586 383734
rect 418822 383498 419004 383734
rect 418404 348054 419004 383498
rect 418404 347818 418586 348054
rect 418822 347818 419004 348054
rect 418404 347734 419004 347818
rect 418404 347498 418586 347734
rect 418822 347498 419004 347734
rect 418404 312054 419004 347498
rect 418404 311818 418586 312054
rect 418822 311818 419004 312054
rect 418404 311734 419004 311818
rect 418404 311498 418586 311734
rect 418822 311498 419004 311734
rect 418404 276054 419004 311498
rect 418404 275818 418586 276054
rect 418822 275818 419004 276054
rect 418404 275734 419004 275818
rect 418404 275498 418586 275734
rect 418822 275498 419004 275734
rect 418404 240054 419004 275498
rect 418404 239818 418586 240054
rect 418822 239818 419004 240054
rect 418404 239734 419004 239818
rect 418404 239498 418586 239734
rect 418822 239498 419004 239734
rect 418404 204054 419004 239498
rect 418404 203818 418586 204054
rect 418822 203818 419004 204054
rect 418404 203734 419004 203818
rect 418404 203498 418586 203734
rect 418822 203498 419004 203734
rect 418404 168054 419004 203498
rect 418404 167818 418586 168054
rect 418822 167818 419004 168054
rect 418404 167734 419004 167818
rect 418404 167498 418586 167734
rect 418822 167498 419004 167734
rect 418404 132054 419004 167498
rect 418404 131818 418586 132054
rect 418822 131818 419004 132054
rect 418404 131734 419004 131818
rect 418404 131498 418586 131734
rect 418822 131498 419004 131734
rect 418404 96054 419004 131498
rect 418404 95818 418586 96054
rect 418822 95818 419004 96054
rect 418404 95734 419004 95818
rect 418404 95498 418586 95734
rect 418822 95498 419004 95734
rect 418404 60054 419004 95498
rect 418404 59818 418586 60054
rect 418822 59818 419004 60054
rect 418404 59734 419004 59818
rect 418404 59498 418586 59734
rect 418822 59498 419004 59734
rect 418404 24054 419004 59498
rect 418404 23818 418586 24054
rect 418822 23818 419004 24054
rect 418404 23734 419004 23818
rect 418404 23498 418586 23734
rect 418822 23498 419004 23734
rect 418404 -3106 419004 23498
rect 418404 -3342 418586 -3106
rect 418822 -3342 419004 -3106
rect 418404 -3426 419004 -3342
rect 418404 -3662 418586 -3426
rect 418822 -3662 419004 -3426
rect 418404 -3684 419004 -3662
rect 422004 675654 422604 708882
rect 422004 675418 422186 675654
rect 422422 675418 422604 675654
rect 422004 675334 422604 675418
rect 422004 675098 422186 675334
rect 422422 675098 422604 675334
rect 422004 639654 422604 675098
rect 422004 639418 422186 639654
rect 422422 639418 422604 639654
rect 422004 639334 422604 639418
rect 422004 639098 422186 639334
rect 422422 639098 422604 639334
rect 422004 603654 422604 639098
rect 422004 603418 422186 603654
rect 422422 603418 422604 603654
rect 422004 603334 422604 603418
rect 422004 603098 422186 603334
rect 422422 603098 422604 603334
rect 422004 567654 422604 603098
rect 422004 567418 422186 567654
rect 422422 567418 422604 567654
rect 422004 567334 422604 567418
rect 422004 567098 422186 567334
rect 422422 567098 422604 567334
rect 422004 531654 422604 567098
rect 425604 679254 426204 710722
rect 443604 710358 444204 711300
rect 443604 710122 443786 710358
rect 444022 710122 444204 710358
rect 443604 710038 444204 710122
rect 443604 709802 443786 710038
rect 444022 709802 444204 710038
rect 440004 708518 440604 709460
rect 440004 708282 440186 708518
rect 440422 708282 440604 708518
rect 440004 708198 440604 708282
rect 440004 707962 440186 708198
rect 440422 707962 440604 708198
rect 436404 706678 437004 707620
rect 436404 706442 436586 706678
rect 436822 706442 437004 706678
rect 436404 706358 437004 706442
rect 436404 706122 436586 706358
rect 436822 706122 437004 706358
rect 425604 679018 425786 679254
rect 426022 679018 426204 679254
rect 425604 678934 426204 679018
rect 425604 678698 425786 678934
rect 426022 678698 426204 678934
rect 425604 643254 426204 678698
rect 425604 643018 425786 643254
rect 426022 643018 426204 643254
rect 425604 642934 426204 643018
rect 425604 642698 425786 642934
rect 426022 642698 426204 642934
rect 425604 607254 426204 642698
rect 425604 607018 425786 607254
rect 426022 607018 426204 607254
rect 425604 606934 426204 607018
rect 425604 606698 425786 606934
rect 426022 606698 426204 606934
rect 425604 571254 426204 606698
rect 425604 571018 425786 571254
rect 426022 571018 426204 571254
rect 425604 570934 426204 571018
rect 425604 570698 425786 570934
rect 426022 570698 426204 570934
rect 422004 531418 422186 531654
rect 422422 531418 422604 531654
rect 422004 531334 422604 531418
rect 422004 531098 422186 531334
rect 422422 531098 422604 531334
rect 422004 495654 422604 531098
rect 422004 495418 422186 495654
rect 422422 495418 422604 495654
rect 422004 495334 422604 495418
rect 422004 495098 422186 495334
rect 422422 495098 422604 495334
rect 422004 459654 422604 495098
rect 422004 459418 422186 459654
rect 422422 459418 422604 459654
rect 422004 459334 422604 459418
rect 422004 459098 422186 459334
rect 422422 459098 422604 459334
rect 422004 423654 422604 459098
rect 422004 423418 422186 423654
rect 422422 423418 422604 423654
rect 422004 423334 422604 423418
rect 422004 423098 422186 423334
rect 422422 423098 422604 423334
rect 422004 387654 422604 423098
rect 422004 387418 422186 387654
rect 422422 387418 422604 387654
rect 422004 387334 422604 387418
rect 422004 387098 422186 387334
rect 422422 387098 422604 387334
rect 422004 351654 422604 387098
rect 422004 351418 422186 351654
rect 422422 351418 422604 351654
rect 422004 351334 422604 351418
rect 422004 351098 422186 351334
rect 422422 351098 422604 351334
rect 422004 315654 422604 351098
rect 422004 315418 422186 315654
rect 422422 315418 422604 315654
rect 422004 315334 422604 315418
rect 422004 315098 422186 315334
rect 422422 315098 422604 315334
rect 422004 279654 422604 315098
rect 422004 279418 422186 279654
rect 422422 279418 422604 279654
rect 422004 279334 422604 279418
rect 422004 279098 422186 279334
rect 422422 279098 422604 279334
rect 422004 243654 422604 279098
rect 422004 243418 422186 243654
rect 422422 243418 422604 243654
rect 422004 243334 422604 243418
rect 422004 243098 422186 243334
rect 422422 243098 422604 243334
rect 422004 207654 422604 243098
rect 422004 207418 422186 207654
rect 422422 207418 422604 207654
rect 422004 207334 422604 207418
rect 422004 207098 422186 207334
rect 422422 207098 422604 207334
rect 422004 171654 422604 207098
rect 422004 171418 422186 171654
rect 422422 171418 422604 171654
rect 422004 171334 422604 171418
rect 422004 171098 422186 171334
rect 422422 171098 422604 171334
rect 422004 135654 422604 171098
rect 422004 135418 422186 135654
rect 422422 135418 422604 135654
rect 422004 135334 422604 135418
rect 422004 135098 422186 135334
rect 422422 135098 422604 135334
rect 422004 99654 422604 135098
rect 422004 99418 422186 99654
rect 422422 99418 422604 99654
rect 422004 99334 422604 99418
rect 422004 99098 422186 99334
rect 422422 99098 422604 99334
rect 422004 63654 422604 99098
rect 422004 63418 422186 63654
rect 422422 63418 422604 63654
rect 422004 63334 422604 63418
rect 422004 63098 422186 63334
rect 422422 63098 422604 63334
rect 422004 27654 422604 63098
rect 422004 27418 422186 27654
rect 422422 27418 422604 27654
rect 422004 27334 422604 27418
rect 422004 27098 422186 27334
rect 422422 27098 422604 27334
rect 422004 -4946 422604 27098
rect 422004 -5182 422186 -4946
rect 422422 -5182 422604 -4946
rect 422004 -5266 422604 -5182
rect 422004 -5502 422186 -5266
rect 422422 -5502 422604 -5266
rect 422004 -5524 422604 -5502
rect 425604 535254 426204 570698
rect 432804 704838 433404 705780
rect 432804 704602 432986 704838
rect 433222 704602 433404 704838
rect 432804 704518 433404 704602
rect 432804 704282 432986 704518
rect 433222 704282 433404 704518
rect 432804 686454 433404 704282
rect 432804 686218 432986 686454
rect 433222 686218 433404 686454
rect 432804 686134 433404 686218
rect 432804 685898 432986 686134
rect 433222 685898 433404 686134
rect 432804 650454 433404 685898
rect 432804 650218 432986 650454
rect 433222 650218 433404 650454
rect 432804 650134 433404 650218
rect 432804 649898 432986 650134
rect 433222 649898 433404 650134
rect 432804 614454 433404 649898
rect 432804 614218 432986 614454
rect 433222 614218 433404 614454
rect 432804 614134 433404 614218
rect 432804 613898 432986 614134
rect 433222 613898 433404 614134
rect 432804 578454 433404 613898
rect 432804 578218 432986 578454
rect 433222 578218 433404 578454
rect 432804 578134 433404 578218
rect 432804 577898 432986 578134
rect 433222 577898 433404 578134
rect 425604 535018 425786 535254
rect 426022 535018 426204 535254
rect 425604 534934 426204 535018
rect 425604 534698 425786 534934
rect 426022 534698 426204 534934
rect 425604 499254 426204 534698
rect 425604 499018 425786 499254
rect 426022 499018 426204 499254
rect 425604 498934 426204 499018
rect 425604 498698 425786 498934
rect 426022 498698 426204 498934
rect 425604 463254 426204 498698
rect 425604 463018 425786 463254
rect 426022 463018 426204 463254
rect 425604 462934 426204 463018
rect 425604 462698 425786 462934
rect 426022 462698 426204 462934
rect 425604 427254 426204 462698
rect 425604 427018 425786 427254
rect 426022 427018 426204 427254
rect 425604 426934 426204 427018
rect 425604 426698 425786 426934
rect 426022 426698 426204 426934
rect 425604 391254 426204 426698
rect 425604 391018 425786 391254
rect 426022 391018 426204 391254
rect 425604 390934 426204 391018
rect 425604 390698 425786 390934
rect 426022 390698 426204 390934
rect 425604 355254 426204 390698
rect 425604 355018 425786 355254
rect 426022 355018 426204 355254
rect 425604 354934 426204 355018
rect 425604 354698 425786 354934
rect 426022 354698 426204 354934
rect 425604 319254 426204 354698
rect 425604 319018 425786 319254
rect 426022 319018 426204 319254
rect 425604 318934 426204 319018
rect 425604 318698 425786 318934
rect 426022 318698 426204 318934
rect 425604 283254 426204 318698
rect 425604 283018 425786 283254
rect 426022 283018 426204 283254
rect 425604 282934 426204 283018
rect 425604 282698 425786 282934
rect 426022 282698 426204 282934
rect 425604 247254 426204 282698
rect 425604 247018 425786 247254
rect 426022 247018 426204 247254
rect 425604 246934 426204 247018
rect 425604 246698 425786 246934
rect 426022 246698 426204 246934
rect 425604 211254 426204 246698
rect 425604 211018 425786 211254
rect 426022 211018 426204 211254
rect 425604 210934 426204 211018
rect 425604 210698 425786 210934
rect 426022 210698 426204 210934
rect 425604 175254 426204 210698
rect 425604 175018 425786 175254
rect 426022 175018 426204 175254
rect 425604 174934 426204 175018
rect 425604 174698 425786 174934
rect 426022 174698 426204 174934
rect 425604 139254 426204 174698
rect 425604 139018 425786 139254
rect 426022 139018 426204 139254
rect 425604 138934 426204 139018
rect 425604 138698 425786 138934
rect 426022 138698 426204 138934
rect 425604 103254 426204 138698
rect 425604 103018 425786 103254
rect 426022 103018 426204 103254
rect 425604 102934 426204 103018
rect 425604 102698 425786 102934
rect 426022 102698 426204 102934
rect 425604 67254 426204 102698
rect 425604 67018 425786 67254
rect 426022 67018 426204 67254
rect 425604 66934 426204 67018
rect 425604 66698 425786 66934
rect 426022 66698 426204 66934
rect 425604 31254 426204 66698
rect 425604 31018 425786 31254
rect 426022 31018 426204 31254
rect 425604 30934 426204 31018
rect 425604 30698 425786 30934
rect 426022 30698 426204 30934
rect 407604 -6102 407786 -5866
rect 408022 -6102 408204 -5866
rect 407604 -6186 408204 -6102
rect 407604 -6422 407786 -6186
rect 408022 -6422 408204 -6186
rect 407604 -7364 408204 -6422
rect 425604 -6786 426204 30698
rect 432804 542454 433404 577898
rect 436404 690054 437004 706122
rect 436404 689818 436586 690054
rect 436822 689818 437004 690054
rect 436404 689734 437004 689818
rect 436404 689498 436586 689734
rect 436822 689498 437004 689734
rect 436404 654054 437004 689498
rect 436404 653818 436586 654054
rect 436822 653818 437004 654054
rect 436404 653734 437004 653818
rect 436404 653498 436586 653734
rect 436822 653498 437004 653734
rect 436404 618054 437004 653498
rect 436404 617818 436586 618054
rect 436822 617818 437004 618054
rect 436404 617734 437004 617818
rect 436404 617498 436586 617734
rect 436822 617498 437004 617734
rect 436404 582054 437004 617498
rect 436404 581818 436586 582054
rect 436822 581818 437004 582054
rect 436404 581734 437004 581818
rect 436404 581498 436586 581734
rect 436822 581498 437004 581734
rect 432804 542218 432986 542454
rect 433222 542218 433404 542454
rect 432804 542134 433404 542218
rect 432804 541898 432986 542134
rect 433222 541898 433404 542134
rect 432804 506454 433404 541898
rect 432804 506218 432986 506454
rect 433222 506218 433404 506454
rect 432804 506134 433404 506218
rect 432804 505898 432986 506134
rect 433222 505898 433404 506134
rect 432804 470454 433404 505898
rect 432804 470218 432986 470454
rect 433222 470218 433404 470454
rect 432804 470134 433404 470218
rect 432804 469898 432986 470134
rect 433222 469898 433404 470134
rect 432804 434454 433404 469898
rect 432804 434218 432986 434454
rect 433222 434218 433404 434454
rect 432804 434134 433404 434218
rect 432804 433898 432986 434134
rect 433222 433898 433404 434134
rect 432804 398454 433404 433898
rect 432804 398218 432986 398454
rect 433222 398218 433404 398454
rect 432804 398134 433404 398218
rect 432804 397898 432986 398134
rect 433222 397898 433404 398134
rect 432804 362454 433404 397898
rect 432804 362218 432986 362454
rect 433222 362218 433404 362454
rect 432804 362134 433404 362218
rect 432804 361898 432986 362134
rect 433222 361898 433404 362134
rect 432804 326454 433404 361898
rect 432804 326218 432986 326454
rect 433222 326218 433404 326454
rect 432804 326134 433404 326218
rect 432804 325898 432986 326134
rect 433222 325898 433404 326134
rect 432804 290454 433404 325898
rect 436404 546054 437004 581498
rect 436404 545818 436586 546054
rect 436822 545818 437004 546054
rect 436404 545734 437004 545818
rect 436404 545498 436586 545734
rect 436822 545498 437004 545734
rect 436404 510054 437004 545498
rect 436404 509818 436586 510054
rect 436822 509818 437004 510054
rect 436404 509734 437004 509818
rect 436404 509498 436586 509734
rect 436822 509498 437004 509734
rect 436404 474054 437004 509498
rect 436404 473818 436586 474054
rect 436822 473818 437004 474054
rect 436404 473734 437004 473818
rect 436404 473498 436586 473734
rect 436822 473498 437004 473734
rect 436404 438054 437004 473498
rect 436404 437818 436586 438054
rect 436822 437818 437004 438054
rect 436404 437734 437004 437818
rect 436404 437498 436586 437734
rect 436822 437498 437004 437734
rect 436404 402054 437004 437498
rect 436404 401818 436586 402054
rect 436822 401818 437004 402054
rect 436404 401734 437004 401818
rect 436404 401498 436586 401734
rect 436822 401498 437004 401734
rect 436404 366054 437004 401498
rect 436404 365818 436586 366054
rect 436822 365818 437004 366054
rect 436404 365734 437004 365818
rect 436404 365498 436586 365734
rect 436822 365498 437004 365734
rect 436404 330054 437004 365498
rect 436404 329818 436586 330054
rect 436822 329818 437004 330054
rect 436404 329734 437004 329818
rect 436404 329498 436586 329734
rect 436822 329498 437004 329734
rect 434483 299436 434549 299437
rect 434483 299372 434484 299436
rect 434548 299372 434549 299436
rect 434483 299371 434549 299372
rect 432804 290218 432986 290454
rect 433222 290218 433404 290454
rect 432804 290134 433404 290218
rect 432804 289898 432986 290134
rect 433222 289898 433404 290134
rect 434486 289917 434546 299371
rect 436404 294054 437004 329498
rect 436404 293818 436586 294054
rect 436822 293818 437004 294054
rect 436404 293734 437004 293818
rect 436404 293498 436586 293734
rect 436822 293498 437004 293734
rect 432804 254454 433404 289898
rect 434483 289916 434549 289917
rect 434483 289852 434484 289916
rect 434548 289852 434549 289916
rect 434483 289851 434549 289852
rect 434483 280124 434549 280125
rect 434483 280060 434484 280124
rect 434548 280060 434549 280124
rect 434483 280059 434549 280060
rect 434486 270605 434546 280059
rect 434483 270604 434549 270605
rect 434483 270540 434484 270604
rect 434548 270540 434549 270604
rect 434483 270539 434549 270540
rect 434483 260812 434549 260813
rect 434483 260748 434484 260812
rect 434548 260748 434549 260812
rect 434483 260747 434549 260748
rect 432804 254218 432986 254454
rect 433222 254218 433404 254454
rect 432804 254134 433404 254218
rect 432804 253898 432986 254134
rect 433222 253898 433404 254134
rect 432804 218454 433404 253898
rect 434486 251293 434546 260747
rect 436404 258054 437004 293498
rect 436404 257818 436586 258054
rect 436822 257818 437004 258054
rect 436404 257734 437004 257818
rect 436404 257498 436586 257734
rect 436822 257498 437004 257734
rect 434483 251292 434549 251293
rect 434483 251228 434484 251292
rect 434548 251228 434549 251292
rect 434483 251227 434549 251228
rect 432804 218218 432986 218454
rect 433222 218218 433404 218454
rect 432804 218134 433404 218218
rect 432804 217898 432986 218134
rect 433222 217898 433404 218134
rect 432804 182454 433404 217898
rect 432804 182218 432986 182454
rect 433222 182218 433404 182454
rect 432804 182134 433404 182218
rect 432804 181898 432986 182134
rect 433222 181898 433404 182134
rect 432804 146454 433404 181898
rect 436404 222054 437004 257498
rect 436404 221818 436586 222054
rect 436822 221818 437004 222054
rect 436404 221734 437004 221818
rect 436404 221498 436586 221734
rect 436822 221498 437004 221734
rect 436404 186054 437004 221498
rect 436404 185818 436586 186054
rect 436822 185818 437004 186054
rect 436404 185734 437004 185818
rect 436404 185498 436586 185734
rect 436822 185498 437004 185734
rect 434299 173908 434365 173909
rect 434299 173844 434300 173908
rect 434364 173844 434365 173908
rect 434299 173843 434365 173844
rect 434302 164253 434362 173843
rect 434299 164252 434365 164253
rect 434299 164188 434300 164252
rect 434364 164188 434365 164252
rect 434299 164187 434365 164188
rect 432804 146218 432986 146454
rect 433222 146218 433404 146454
rect 432804 146134 433404 146218
rect 432804 145898 432986 146134
rect 433222 145898 433404 146134
rect 432804 110454 433404 145898
rect 432804 110218 432986 110454
rect 433222 110218 433404 110454
rect 432804 110134 433404 110218
rect 432804 109898 432986 110134
rect 433222 109898 433404 110134
rect 432804 74454 433404 109898
rect 432804 74218 432986 74454
rect 433222 74218 433404 74454
rect 432804 74134 433404 74218
rect 432804 73898 432986 74134
rect 433222 73898 433404 74134
rect 432804 38454 433404 73898
rect 436404 150054 437004 185498
rect 436404 149818 436586 150054
rect 436822 149818 437004 150054
rect 436404 149734 437004 149818
rect 436404 149498 436586 149734
rect 436822 149498 437004 149734
rect 436404 114054 437004 149498
rect 436404 113818 436586 114054
rect 436822 113818 437004 114054
rect 436404 113734 437004 113818
rect 436404 113498 436586 113734
rect 436822 113498 437004 113734
rect 436404 78054 437004 113498
rect 436404 77818 436586 78054
rect 436822 77818 437004 78054
rect 436404 77734 437004 77818
rect 436404 77498 436586 77734
rect 436822 77498 437004 77734
rect 434299 48244 434365 48245
rect 434299 48180 434300 48244
rect 434364 48180 434365 48244
rect 434299 48179 434365 48180
rect 434302 41309 434362 48179
rect 436404 42054 437004 77498
rect 436404 41818 436586 42054
rect 436822 41818 437004 42054
rect 436404 41734 437004 41818
rect 436404 41498 436586 41734
rect 436822 41498 437004 41734
rect 434299 41308 434365 41309
rect 434299 41244 434300 41308
rect 434364 41244 434365 41308
rect 434299 41243 434365 41244
rect 432804 38218 432986 38454
rect 433222 38218 433404 38454
rect 432804 38134 433404 38218
rect 432804 37898 432986 38134
rect 433222 37898 433404 38134
rect 432804 2454 433404 37898
rect 432804 2218 432986 2454
rect 433222 2218 433404 2454
rect 432804 2134 433404 2218
rect 432804 1898 432986 2134
rect 433222 1898 433404 2134
rect 432804 -346 433404 1898
rect 432804 -582 432986 -346
rect 433222 -582 433404 -346
rect 432804 -666 433404 -582
rect 432804 -902 432986 -666
rect 433222 -902 433404 -666
rect 432804 -1844 433404 -902
rect 436404 6054 437004 41498
rect 436404 5818 436586 6054
rect 436822 5818 437004 6054
rect 436404 5734 437004 5818
rect 436404 5498 436586 5734
rect 436822 5498 437004 5734
rect 436404 -2186 437004 5498
rect 436404 -2422 436586 -2186
rect 436822 -2422 437004 -2186
rect 436404 -2506 437004 -2422
rect 436404 -2742 436586 -2506
rect 436822 -2742 437004 -2506
rect 436404 -3684 437004 -2742
rect 440004 693654 440604 707962
rect 440004 693418 440186 693654
rect 440422 693418 440604 693654
rect 440004 693334 440604 693418
rect 440004 693098 440186 693334
rect 440422 693098 440604 693334
rect 440004 657654 440604 693098
rect 440004 657418 440186 657654
rect 440422 657418 440604 657654
rect 440004 657334 440604 657418
rect 440004 657098 440186 657334
rect 440422 657098 440604 657334
rect 440004 621654 440604 657098
rect 440004 621418 440186 621654
rect 440422 621418 440604 621654
rect 440004 621334 440604 621418
rect 440004 621098 440186 621334
rect 440422 621098 440604 621334
rect 440004 585654 440604 621098
rect 440004 585418 440186 585654
rect 440422 585418 440604 585654
rect 440004 585334 440604 585418
rect 440004 585098 440186 585334
rect 440422 585098 440604 585334
rect 440004 549654 440604 585098
rect 440004 549418 440186 549654
rect 440422 549418 440604 549654
rect 440004 549334 440604 549418
rect 440004 549098 440186 549334
rect 440422 549098 440604 549334
rect 440004 513654 440604 549098
rect 440004 513418 440186 513654
rect 440422 513418 440604 513654
rect 440004 513334 440604 513418
rect 440004 513098 440186 513334
rect 440422 513098 440604 513334
rect 440004 477654 440604 513098
rect 440004 477418 440186 477654
rect 440422 477418 440604 477654
rect 440004 477334 440604 477418
rect 440004 477098 440186 477334
rect 440422 477098 440604 477334
rect 440004 441654 440604 477098
rect 440004 441418 440186 441654
rect 440422 441418 440604 441654
rect 440004 441334 440604 441418
rect 440004 441098 440186 441334
rect 440422 441098 440604 441334
rect 440004 405654 440604 441098
rect 440004 405418 440186 405654
rect 440422 405418 440604 405654
rect 440004 405334 440604 405418
rect 440004 405098 440186 405334
rect 440422 405098 440604 405334
rect 440004 369654 440604 405098
rect 440004 369418 440186 369654
rect 440422 369418 440604 369654
rect 440004 369334 440604 369418
rect 440004 369098 440186 369334
rect 440422 369098 440604 369334
rect 440004 333654 440604 369098
rect 440004 333418 440186 333654
rect 440422 333418 440604 333654
rect 440004 333334 440604 333418
rect 440004 333098 440186 333334
rect 440422 333098 440604 333334
rect 440004 297654 440604 333098
rect 440004 297418 440186 297654
rect 440422 297418 440604 297654
rect 440004 297334 440604 297418
rect 440004 297098 440186 297334
rect 440422 297098 440604 297334
rect 440004 261654 440604 297098
rect 440004 261418 440186 261654
rect 440422 261418 440604 261654
rect 440004 261334 440604 261418
rect 440004 261098 440186 261334
rect 440422 261098 440604 261334
rect 440004 225654 440604 261098
rect 440004 225418 440186 225654
rect 440422 225418 440604 225654
rect 440004 225334 440604 225418
rect 440004 225098 440186 225334
rect 440422 225098 440604 225334
rect 440004 189654 440604 225098
rect 440004 189418 440186 189654
rect 440422 189418 440604 189654
rect 440004 189334 440604 189418
rect 440004 189098 440186 189334
rect 440422 189098 440604 189334
rect 440004 153654 440604 189098
rect 440004 153418 440186 153654
rect 440422 153418 440604 153654
rect 440004 153334 440604 153418
rect 440004 153098 440186 153334
rect 440422 153098 440604 153334
rect 440004 117654 440604 153098
rect 440004 117418 440186 117654
rect 440422 117418 440604 117654
rect 440004 117334 440604 117418
rect 440004 117098 440186 117334
rect 440422 117098 440604 117334
rect 440004 81654 440604 117098
rect 440004 81418 440186 81654
rect 440422 81418 440604 81654
rect 440004 81334 440604 81418
rect 440004 81098 440186 81334
rect 440422 81098 440604 81334
rect 440004 45654 440604 81098
rect 440004 45418 440186 45654
rect 440422 45418 440604 45654
rect 440004 45334 440604 45418
rect 440004 45098 440186 45334
rect 440422 45098 440604 45334
rect 440004 9654 440604 45098
rect 440004 9418 440186 9654
rect 440422 9418 440604 9654
rect 440004 9334 440604 9418
rect 440004 9098 440186 9334
rect 440422 9098 440604 9334
rect 440004 -4026 440604 9098
rect 440004 -4262 440186 -4026
rect 440422 -4262 440604 -4026
rect 440004 -4346 440604 -4262
rect 440004 -4582 440186 -4346
rect 440422 -4582 440604 -4346
rect 440004 -5524 440604 -4582
rect 443604 697254 444204 709802
rect 461604 711278 462204 711300
rect 461604 711042 461786 711278
rect 462022 711042 462204 711278
rect 461604 710958 462204 711042
rect 461604 710722 461786 710958
rect 462022 710722 462204 710958
rect 458004 709438 458604 709460
rect 458004 709202 458186 709438
rect 458422 709202 458604 709438
rect 458004 709118 458604 709202
rect 458004 708882 458186 709118
rect 458422 708882 458604 709118
rect 454404 707598 455004 707620
rect 454404 707362 454586 707598
rect 454822 707362 455004 707598
rect 454404 707278 455004 707362
rect 454404 707042 454586 707278
rect 454822 707042 455004 707278
rect 443604 697018 443786 697254
rect 444022 697018 444204 697254
rect 443604 696934 444204 697018
rect 443604 696698 443786 696934
rect 444022 696698 444204 696934
rect 443604 661254 444204 696698
rect 443604 661018 443786 661254
rect 444022 661018 444204 661254
rect 443604 660934 444204 661018
rect 443604 660698 443786 660934
rect 444022 660698 444204 660934
rect 443604 625254 444204 660698
rect 443604 625018 443786 625254
rect 444022 625018 444204 625254
rect 443604 624934 444204 625018
rect 443604 624698 443786 624934
rect 444022 624698 444204 624934
rect 443604 589254 444204 624698
rect 443604 589018 443786 589254
rect 444022 589018 444204 589254
rect 443604 588934 444204 589018
rect 443604 588698 443786 588934
rect 444022 588698 444204 588934
rect 443604 553254 444204 588698
rect 450804 705758 451404 705780
rect 450804 705522 450986 705758
rect 451222 705522 451404 705758
rect 450804 705438 451404 705522
rect 450804 705202 450986 705438
rect 451222 705202 451404 705438
rect 450804 668454 451404 705202
rect 450804 668218 450986 668454
rect 451222 668218 451404 668454
rect 450804 668134 451404 668218
rect 450804 667898 450986 668134
rect 451222 667898 451404 668134
rect 450804 632454 451404 667898
rect 450804 632218 450986 632454
rect 451222 632218 451404 632454
rect 450804 632134 451404 632218
rect 450804 631898 450986 632134
rect 451222 631898 451404 632134
rect 450804 596454 451404 631898
rect 450804 596218 450986 596454
rect 451222 596218 451404 596454
rect 450804 596134 451404 596218
rect 450804 595898 450986 596134
rect 451222 595898 451404 596134
rect 446259 563004 446325 563005
rect 446259 562940 446260 563004
rect 446324 562940 446325 563004
rect 446259 562939 446325 562940
rect 444419 559332 444485 559333
rect 444419 559268 444420 559332
rect 444484 559268 444485 559332
rect 444419 559267 444485 559268
rect 445707 559332 445773 559333
rect 445707 559268 445708 559332
rect 445772 559268 445773 559332
rect 445707 559267 445773 559268
rect 443604 553018 443786 553254
rect 444022 553018 444204 553254
rect 443604 552934 444204 553018
rect 443604 552698 443786 552934
rect 444022 552698 444204 552934
rect 443604 517254 444204 552698
rect 443604 517018 443786 517254
rect 444022 517018 444204 517254
rect 443604 516934 444204 517018
rect 443604 516698 443786 516934
rect 444022 516698 444204 516934
rect 443604 481254 444204 516698
rect 443604 481018 443786 481254
rect 444022 481018 444204 481254
rect 443604 480934 444204 481018
rect 443604 480698 443786 480934
rect 444022 480698 444204 480934
rect 443604 445254 444204 480698
rect 443604 445018 443786 445254
rect 444022 445018 444204 445254
rect 443604 444934 444204 445018
rect 443604 444698 443786 444934
rect 444022 444698 444204 444934
rect 443604 409254 444204 444698
rect 443604 409018 443786 409254
rect 444022 409018 444204 409254
rect 443604 408934 444204 409018
rect 443604 408698 443786 408934
rect 444022 408698 444204 408934
rect 443604 373254 444204 408698
rect 443604 373018 443786 373254
rect 444022 373018 444204 373254
rect 443604 372934 444204 373018
rect 443604 372698 443786 372934
rect 444022 372698 444204 372934
rect 443604 337254 444204 372698
rect 443604 337018 443786 337254
rect 444022 337018 444204 337254
rect 443604 336934 444204 337018
rect 443604 336698 443786 336934
rect 444022 336698 444204 336934
rect 443604 301254 444204 336698
rect 443604 301018 443786 301254
rect 444022 301018 444204 301254
rect 443604 300934 444204 301018
rect 443604 300698 443786 300934
rect 444022 300698 444204 300934
rect 443604 265254 444204 300698
rect 443604 265018 443786 265254
rect 444022 265018 444204 265254
rect 443604 264934 444204 265018
rect 443604 264698 443786 264934
rect 444022 264698 444204 264934
rect 443604 229254 444204 264698
rect 443604 229018 443786 229254
rect 444022 229018 444204 229254
rect 443604 228934 444204 229018
rect 443604 228698 443786 228934
rect 444022 228698 444204 228934
rect 443604 193254 444204 228698
rect 443604 193018 443786 193254
rect 444022 193018 444204 193254
rect 443604 192934 444204 193018
rect 443604 192698 443786 192934
rect 444022 192698 444204 192934
rect 443604 157254 444204 192698
rect 443604 157018 443786 157254
rect 444022 157018 444204 157254
rect 443604 156934 444204 157018
rect 443604 156698 443786 156934
rect 444022 156698 444204 156934
rect 443604 121254 444204 156698
rect 443604 121018 443786 121254
rect 444022 121018 444204 121254
rect 443604 120934 444204 121018
rect 443604 120698 443786 120934
rect 444022 120698 444204 120934
rect 443604 85254 444204 120698
rect 443604 85018 443786 85254
rect 444022 85018 444204 85254
rect 443604 84934 444204 85018
rect 443604 84698 443786 84934
rect 444022 84698 444204 84934
rect 443604 49254 444204 84698
rect 443604 49018 443786 49254
rect 444022 49018 444204 49254
rect 443604 48934 444204 49018
rect 443604 48698 443786 48934
rect 444022 48698 444204 48934
rect 443604 13254 444204 48698
rect 444422 35869 444482 559267
rect 444419 35868 444485 35869
rect 444419 35804 444420 35868
rect 444484 35804 444485 35868
rect 444419 35803 444485 35804
rect 443604 13018 443786 13254
rect 444022 13018 444204 13254
rect 443604 12934 444204 13018
rect 443604 12698 443786 12934
rect 444022 12698 444204 12934
rect 425604 -7022 425786 -6786
rect 426022 -7022 426204 -6786
rect 425604 -7106 426204 -7022
rect 425604 -7342 425786 -7106
rect 426022 -7342 426204 -7106
rect 425604 -7364 426204 -7342
rect 443604 -5866 444204 12698
rect 445710 8261 445770 559267
rect 446262 486165 446322 562939
rect 450804 560454 451404 595898
rect 447731 560284 447797 560285
rect 447731 560220 447732 560284
rect 447796 560220 447797 560284
rect 447731 560219 447797 560220
rect 446259 486164 446325 486165
rect 446259 486100 446260 486164
rect 446324 486100 446325 486164
rect 446259 486099 446325 486100
rect 447734 204645 447794 560219
rect 450804 560218 450986 560454
rect 451222 560218 451404 560454
rect 450804 560134 451404 560218
rect 450804 559898 450986 560134
rect 451222 559898 451404 560134
rect 448467 559332 448533 559333
rect 448467 559268 448468 559332
rect 448532 559268 448533 559332
rect 448467 559267 448533 559268
rect 447731 204644 447797 204645
rect 447731 204580 447732 204644
rect 447796 204580 447797 204644
rect 447731 204579 447797 204580
rect 448470 21997 448530 559267
rect 450804 524454 451404 559898
rect 450804 524218 450986 524454
rect 451222 524218 451404 524454
rect 450804 524134 451404 524218
rect 450804 523898 450986 524134
rect 451222 523898 451404 524134
rect 450804 488454 451404 523898
rect 450804 488218 450986 488454
rect 451222 488218 451404 488454
rect 450804 488134 451404 488218
rect 450804 487898 450986 488134
rect 451222 487898 451404 488134
rect 450804 452454 451404 487898
rect 450804 452218 450986 452454
rect 451222 452218 451404 452454
rect 450804 452134 451404 452218
rect 450804 451898 450986 452134
rect 451222 451898 451404 452134
rect 450804 416454 451404 451898
rect 450804 416218 450986 416454
rect 451222 416218 451404 416454
rect 450804 416134 451404 416218
rect 450804 415898 450986 416134
rect 451222 415898 451404 416134
rect 450804 380454 451404 415898
rect 450804 380218 450986 380454
rect 451222 380218 451404 380454
rect 450804 380134 451404 380218
rect 450804 379898 450986 380134
rect 451222 379898 451404 380134
rect 450804 344454 451404 379898
rect 450804 344218 450986 344454
rect 451222 344218 451404 344454
rect 450804 344134 451404 344218
rect 450804 343898 450986 344134
rect 451222 343898 451404 344134
rect 450804 308454 451404 343898
rect 450804 308218 450986 308454
rect 451222 308218 451404 308454
rect 450804 308134 451404 308218
rect 450804 307898 450986 308134
rect 451222 307898 451404 308134
rect 450804 272454 451404 307898
rect 450804 272218 450986 272454
rect 451222 272218 451404 272454
rect 450804 272134 451404 272218
rect 450804 271898 450986 272134
rect 451222 271898 451404 272134
rect 450804 236454 451404 271898
rect 450804 236218 450986 236454
rect 451222 236218 451404 236454
rect 450804 236134 451404 236218
rect 450804 235898 450986 236134
rect 451222 235898 451404 236134
rect 450804 200454 451404 235898
rect 450804 200218 450986 200454
rect 451222 200218 451404 200454
rect 450804 200134 451404 200218
rect 450804 199898 450986 200134
rect 451222 199898 451404 200134
rect 450804 164454 451404 199898
rect 450804 164218 450986 164454
rect 451222 164218 451404 164454
rect 450804 164134 451404 164218
rect 450804 163898 450986 164134
rect 451222 163898 451404 164134
rect 450804 128454 451404 163898
rect 454404 672054 455004 707042
rect 454404 671818 454586 672054
rect 454822 671818 455004 672054
rect 454404 671734 455004 671818
rect 454404 671498 454586 671734
rect 454822 671498 455004 671734
rect 454404 636054 455004 671498
rect 454404 635818 454586 636054
rect 454822 635818 455004 636054
rect 454404 635734 455004 635818
rect 454404 635498 454586 635734
rect 454822 635498 455004 635734
rect 454404 600054 455004 635498
rect 454404 599818 454586 600054
rect 454822 599818 455004 600054
rect 454404 599734 455004 599818
rect 454404 599498 454586 599734
rect 454822 599498 455004 599734
rect 454404 564054 455004 599498
rect 454404 563818 454586 564054
rect 454822 563818 455004 564054
rect 454404 563734 455004 563818
rect 454404 563498 454586 563734
rect 454822 563498 455004 563734
rect 454404 528054 455004 563498
rect 454404 527818 454586 528054
rect 454822 527818 455004 528054
rect 454404 527734 455004 527818
rect 454404 527498 454586 527734
rect 454822 527498 455004 527734
rect 454404 492054 455004 527498
rect 454404 491818 454586 492054
rect 454822 491818 455004 492054
rect 454404 491734 455004 491818
rect 454404 491498 454586 491734
rect 454822 491498 455004 491734
rect 454404 456054 455004 491498
rect 454404 455818 454586 456054
rect 454822 455818 455004 456054
rect 454404 455734 455004 455818
rect 454404 455498 454586 455734
rect 454822 455498 455004 455734
rect 454404 420054 455004 455498
rect 454404 419818 454586 420054
rect 454822 419818 455004 420054
rect 454404 419734 455004 419818
rect 454404 419498 454586 419734
rect 454822 419498 455004 419734
rect 454404 384054 455004 419498
rect 454404 383818 454586 384054
rect 454822 383818 455004 384054
rect 454404 383734 455004 383818
rect 454404 383498 454586 383734
rect 454822 383498 455004 383734
rect 454404 348054 455004 383498
rect 454404 347818 454586 348054
rect 454822 347818 455004 348054
rect 454404 347734 455004 347818
rect 454404 347498 454586 347734
rect 454822 347498 455004 347734
rect 454404 312054 455004 347498
rect 454404 311818 454586 312054
rect 454822 311818 455004 312054
rect 454404 311734 455004 311818
rect 454404 311498 454586 311734
rect 454822 311498 455004 311734
rect 454404 276054 455004 311498
rect 454404 275818 454586 276054
rect 454822 275818 455004 276054
rect 454404 275734 455004 275818
rect 454404 275498 454586 275734
rect 454822 275498 455004 275734
rect 454404 240054 455004 275498
rect 454404 239818 454586 240054
rect 454822 239818 455004 240054
rect 454404 239734 455004 239818
rect 454404 239498 454586 239734
rect 454822 239498 455004 239734
rect 454404 204054 455004 239498
rect 454404 203818 454586 204054
rect 454822 203818 455004 204054
rect 454404 203734 455004 203818
rect 454404 203498 454586 203734
rect 454822 203498 455004 203734
rect 454404 168054 455004 203498
rect 454404 167818 454586 168054
rect 454822 167818 455004 168054
rect 454404 167734 455004 167818
rect 454404 167498 454586 167734
rect 454822 167498 455004 167734
rect 453987 134604 454053 134605
rect 453987 134540 453988 134604
rect 454052 134540 454053 134604
rect 453987 134539 454053 134540
rect 453990 134333 454050 134539
rect 453987 134332 454053 134333
rect 453987 134268 453988 134332
rect 454052 134268 454053 134332
rect 453987 134267 454053 134268
rect 450804 128218 450986 128454
rect 451222 128218 451404 128454
rect 450804 128134 451404 128218
rect 450804 127898 450986 128134
rect 451222 127898 451404 128134
rect 450804 92454 451404 127898
rect 450804 92218 450986 92454
rect 451222 92218 451404 92454
rect 450804 92134 451404 92218
rect 450804 91898 450986 92134
rect 451222 91898 451404 92134
rect 450804 56454 451404 91898
rect 454404 132054 455004 167498
rect 454404 131818 454586 132054
rect 454822 131818 455004 132054
rect 454404 131734 455004 131818
rect 454404 131498 454586 131734
rect 454822 131498 455004 131734
rect 454404 96054 455004 131498
rect 454404 95818 454586 96054
rect 454822 95818 455004 96054
rect 454404 95734 455004 95818
rect 454404 95498 454586 95734
rect 454822 95498 455004 95734
rect 453987 87548 454053 87549
rect 453987 87484 453988 87548
rect 454052 87484 454053 87548
rect 453987 87483 454053 87484
rect 453990 87277 454050 87483
rect 453987 87276 454053 87277
rect 453987 87212 453988 87276
rect 454052 87212 454053 87276
rect 453987 87211 454053 87212
rect 453987 64292 454053 64293
rect 453987 64228 453988 64292
rect 454052 64228 454053 64292
rect 453987 64227 454053 64228
rect 453990 64021 454050 64227
rect 453987 64020 454053 64021
rect 453987 63956 453988 64020
rect 454052 63956 454053 64020
rect 453987 63955 454053 63956
rect 450804 56218 450986 56454
rect 451222 56218 451404 56454
rect 450804 56134 451404 56218
rect 450804 55898 450986 56134
rect 451222 55898 451404 56134
rect 448467 21996 448533 21997
rect 448467 21932 448468 21996
rect 448532 21932 448533 21996
rect 448467 21931 448533 21932
rect 450804 20454 451404 55898
rect 454404 60054 455004 95498
rect 454404 59818 454586 60054
rect 454822 59818 455004 60054
rect 454404 59734 455004 59818
rect 454404 59498 454586 59734
rect 454822 59498 455004 59734
rect 453987 40764 454053 40765
rect 453987 40700 453988 40764
rect 454052 40700 454053 40764
rect 453987 40699 454053 40700
rect 453990 40493 454050 40699
rect 453987 40492 454053 40493
rect 453987 40428 453988 40492
rect 454052 40428 454053 40492
rect 453987 40427 454053 40428
rect 450804 20218 450986 20454
rect 451222 20218 451404 20454
rect 450804 20134 451404 20218
rect 450804 19898 450986 20134
rect 451222 19898 451404 20134
rect 445707 8260 445773 8261
rect 445707 8196 445708 8260
rect 445772 8196 445773 8260
rect 445707 8195 445773 8196
rect 450804 -1266 451404 19898
rect 450804 -1502 450986 -1266
rect 451222 -1502 451404 -1266
rect 450804 -1586 451404 -1502
rect 450804 -1822 450986 -1586
rect 451222 -1822 451404 -1586
rect 450804 -1844 451404 -1822
rect 454404 24054 455004 59498
rect 454404 23818 454586 24054
rect 454822 23818 455004 24054
rect 454404 23734 455004 23818
rect 454404 23498 454586 23734
rect 454822 23498 455004 23734
rect 454404 -3106 455004 23498
rect 454404 -3342 454586 -3106
rect 454822 -3342 455004 -3106
rect 454404 -3426 455004 -3342
rect 454404 -3662 454586 -3426
rect 454822 -3662 455004 -3426
rect 454404 -3684 455004 -3662
rect 458004 675654 458604 708882
rect 458004 675418 458186 675654
rect 458422 675418 458604 675654
rect 458004 675334 458604 675418
rect 458004 675098 458186 675334
rect 458422 675098 458604 675334
rect 458004 639654 458604 675098
rect 458004 639418 458186 639654
rect 458422 639418 458604 639654
rect 458004 639334 458604 639418
rect 458004 639098 458186 639334
rect 458422 639098 458604 639334
rect 458004 603654 458604 639098
rect 458004 603418 458186 603654
rect 458422 603418 458604 603654
rect 458004 603334 458604 603418
rect 458004 603098 458186 603334
rect 458422 603098 458604 603334
rect 458004 567654 458604 603098
rect 458004 567418 458186 567654
rect 458422 567418 458604 567654
rect 458004 567334 458604 567418
rect 458004 567098 458186 567334
rect 458422 567098 458604 567334
rect 458004 531654 458604 567098
rect 458004 531418 458186 531654
rect 458422 531418 458604 531654
rect 458004 531334 458604 531418
rect 458004 531098 458186 531334
rect 458422 531098 458604 531334
rect 458004 495654 458604 531098
rect 458004 495418 458186 495654
rect 458422 495418 458604 495654
rect 458004 495334 458604 495418
rect 458004 495098 458186 495334
rect 458422 495098 458604 495334
rect 458004 459654 458604 495098
rect 458004 459418 458186 459654
rect 458422 459418 458604 459654
rect 458004 459334 458604 459418
rect 458004 459098 458186 459334
rect 458422 459098 458604 459334
rect 458004 423654 458604 459098
rect 458004 423418 458186 423654
rect 458422 423418 458604 423654
rect 458004 423334 458604 423418
rect 458004 423098 458186 423334
rect 458422 423098 458604 423334
rect 458004 387654 458604 423098
rect 458004 387418 458186 387654
rect 458422 387418 458604 387654
rect 458004 387334 458604 387418
rect 458004 387098 458186 387334
rect 458422 387098 458604 387334
rect 458004 351654 458604 387098
rect 458004 351418 458186 351654
rect 458422 351418 458604 351654
rect 458004 351334 458604 351418
rect 458004 351098 458186 351334
rect 458422 351098 458604 351334
rect 458004 315654 458604 351098
rect 458004 315418 458186 315654
rect 458422 315418 458604 315654
rect 458004 315334 458604 315418
rect 458004 315098 458186 315334
rect 458422 315098 458604 315334
rect 458004 279654 458604 315098
rect 458004 279418 458186 279654
rect 458422 279418 458604 279654
rect 458004 279334 458604 279418
rect 458004 279098 458186 279334
rect 458422 279098 458604 279334
rect 458004 243654 458604 279098
rect 458004 243418 458186 243654
rect 458422 243418 458604 243654
rect 458004 243334 458604 243418
rect 458004 243098 458186 243334
rect 458422 243098 458604 243334
rect 458004 207654 458604 243098
rect 458004 207418 458186 207654
rect 458422 207418 458604 207654
rect 458004 207334 458604 207418
rect 458004 207098 458186 207334
rect 458422 207098 458604 207334
rect 458004 171654 458604 207098
rect 458004 171418 458186 171654
rect 458422 171418 458604 171654
rect 458004 171334 458604 171418
rect 458004 171098 458186 171334
rect 458422 171098 458604 171334
rect 458004 135654 458604 171098
rect 458004 135418 458186 135654
rect 458422 135418 458604 135654
rect 458004 135334 458604 135418
rect 458004 135098 458186 135334
rect 458422 135098 458604 135334
rect 458004 99654 458604 135098
rect 458004 99418 458186 99654
rect 458422 99418 458604 99654
rect 458004 99334 458604 99418
rect 458004 99098 458186 99334
rect 458422 99098 458604 99334
rect 458004 63654 458604 99098
rect 458004 63418 458186 63654
rect 458422 63418 458604 63654
rect 458004 63334 458604 63418
rect 458004 63098 458186 63334
rect 458422 63098 458604 63334
rect 458004 27654 458604 63098
rect 458004 27418 458186 27654
rect 458422 27418 458604 27654
rect 458004 27334 458604 27418
rect 458004 27098 458186 27334
rect 458422 27098 458604 27334
rect 458004 -4946 458604 27098
rect 458004 -5182 458186 -4946
rect 458422 -5182 458604 -4946
rect 458004 -5266 458604 -5182
rect 458004 -5502 458186 -5266
rect 458422 -5502 458604 -5266
rect 458004 -5524 458604 -5502
rect 461604 679254 462204 710722
rect 479604 710358 480204 711300
rect 479604 710122 479786 710358
rect 480022 710122 480204 710358
rect 479604 710038 480204 710122
rect 479604 709802 479786 710038
rect 480022 709802 480204 710038
rect 476004 708518 476604 709460
rect 476004 708282 476186 708518
rect 476422 708282 476604 708518
rect 476004 708198 476604 708282
rect 476004 707962 476186 708198
rect 476422 707962 476604 708198
rect 472404 706678 473004 707620
rect 472404 706442 472586 706678
rect 472822 706442 473004 706678
rect 472404 706358 473004 706442
rect 472404 706122 472586 706358
rect 472822 706122 473004 706358
rect 461604 679018 461786 679254
rect 462022 679018 462204 679254
rect 461604 678934 462204 679018
rect 461604 678698 461786 678934
rect 462022 678698 462204 678934
rect 461604 643254 462204 678698
rect 461604 643018 461786 643254
rect 462022 643018 462204 643254
rect 461604 642934 462204 643018
rect 461604 642698 461786 642934
rect 462022 642698 462204 642934
rect 461604 607254 462204 642698
rect 461604 607018 461786 607254
rect 462022 607018 462204 607254
rect 461604 606934 462204 607018
rect 461604 606698 461786 606934
rect 462022 606698 462204 606934
rect 461604 571254 462204 606698
rect 461604 571018 461786 571254
rect 462022 571018 462204 571254
rect 461604 570934 462204 571018
rect 461604 570698 461786 570934
rect 462022 570698 462204 570934
rect 461604 535254 462204 570698
rect 461604 535018 461786 535254
rect 462022 535018 462204 535254
rect 461604 534934 462204 535018
rect 461604 534698 461786 534934
rect 462022 534698 462204 534934
rect 461604 499254 462204 534698
rect 461604 499018 461786 499254
rect 462022 499018 462204 499254
rect 461604 498934 462204 499018
rect 461604 498698 461786 498934
rect 462022 498698 462204 498934
rect 461604 463254 462204 498698
rect 461604 463018 461786 463254
rect 462022 463018 462204 463254
rect 461604 462934 462204 463018
rect 461604 462698 461786 462934
rect 462022 462698 462204 462934
rect 461604 427254 462204 462698
rect 461604 427018 461786 427254
rect 462022 427018 462204 427254
rect 461604 426934 462204 427018
rect 461604 426698 461786 426934
rect 462022 426698 462204 426934
rect 461604 391254 462204 426698
rect 461604 391018 461786 391254
rect 462022 391018 462204 391254
rect 461604 390934 462204 391018
rect 461604 390698 461786 390934
rect 462022 390698 462204 390934
rect 461604 355254 462204 390698
rect 461604 355018 461786 355254
rect 462022 355018 462204 355254
rect 461604 354934 462204 355018
rect 461604 354698 461786 354934
rect 462022 354698 462204 354934
rect 461604 319254 462204 354698
rect 461604 319018 461786 319254
rect 462022 319018 462204 319254
rect 461604 318934 462204 319018
rect 461604 318698 461786 318934
rect 462022 318698 462204 318934
rect 461604 283254 462204 318698
rect 461604 283018 461786 283254
rect 462022 283018 462204 283254
rect 461604 282934 462204 283018
rect 461604 282698 461786 282934
rect 462022 282698 462204 282934
rect 461604 247254 462204 282698
rect 461604 247018 461786 247254
rect 462022 247018 462204 247254
rect 461604 246934 462204 247018
rect 461604 246698 461786 246934
rect 462022 246698 462204 246934
rect 461604 211254 462204 246698
rect 461604 211018 461786 211254
rect 462022 211018 462204 211254
rect 461604 210934 462204 211018
rect 461604 210698 461786 210934
rect 462022 210698 462204 210934
rect 461604 175254 462204 210698
rect 461604 175018 461786 175254
rect 462022 175018 462204 175254
rect 461604 174934 462204 175018
rect 461604 174698 461786 174934
rect 462022 174698 462204 174934
rect 461604 139254 462204 174698
rect 461604 139018 461786 139254
rect 462022 139018 462204 139254
rect 461604 138934 462204 139018
rect 461604 138698 461786 138934
rect 462022 138698 462204 138934
rect 461604 103254 462204 138698
rect 461604 103018 461786 103254
rect 462022 103018 462204 103254
rect 461604 102934 462204 103018
rect 461604 102698 461786 102934
rect 462022 102698 462204 102934
rect 461604 67254 462204 102698
rect 461604 67018 461786 67254
rect 462022 67018 462204 67254
rect 461604 66934 462204 67018
rect 461604 66698 461786 66934
rect 462022 66698 462204 66934
rect 461604 31254 462204 66698
rect 461604 31018 461786 31254
rect 462022 31018 462204 31254
rect 461604 30934 462204 31018
rect 461604 30698 461786 30934
rect 462022 30698 462204 30934
rect 443604 -6102 443786 -5866
rect 444022 -6102 444204 -5866
rect 443604 -6186 444204 -6102
rect 443604 -6422 443786 -6186
rect 444022 -6422 444204 -6186
rect 443604 -7364 444204 -6422
rect 461604 -6786 462204 30698
rect 468804 704838 469404 705780
rect 468804 704602 468986 704838
rect 469222 704602 469404 704838
rect 468804 704518 469404 704602
rect 468804 704282 468986 704518
rect 469222 704282 469404 704518
rect 468804 686454 469404 704282
rect 468804 686218 468986 686454
rect 469222 686218 469404 686454
rect 468804 686134 469404 686218
rect 468804 685898 468986 686134
rect 469222 685898 469404 686134
rect 468804 650454 469404 685898
rect 468804 650218 468986 650454
rect 469222 650218 469404 650454
rect 468804 650134 469404 650218
rect 468804 649898 468986 650134
rect 469222 649898 469404 650134
rect 468804 614454 469404 649898
rect 468804 614218 468986 614454
rect 469222 614218 469404 614454
rect 468804 614134 469404 614218
rect 468804 613898 468986 614134
rect 469222 613898 469404 614134
rect 468804 578454 469404 613898
rect 468804 578218 468986 578454
rect 469222 578218 469404 578454
rect 468804 578134 469404 578218
rect 468804 577898 468986 578134
rect 469222 577898 469404 578134
rect 468804 542454 469404 577898
rect 468804 542218 468986 542454
rect 469222 542218 469404 542454
rect 468804 542134 469404 542218
rect 468804 541898 468986 542134
rect 469222 541898 469404 542134
rect 468804 506454 469404 541898
rect 468804 506218 468986 506454
rect 469222 506218 469404 506454
rect 468804 506134 469404 506218
rect 468804 505898 468986 506134
rect 469222 505898 469404 506134
rect 468804 470454 469404 505898
rect 468804 470218 468986 470454
rect 469222 470218 469404 470454
rect 468804 470134 469404 470218
rect 468804 469898 468986 470134
rect 469222 469898 469404 470134
rect 468804 434454 469404 469898
rect 468804 434218 468986 434454
rect 469222 434218 469404 434454
rect 468804 434134 469404 434218
rect 468804 433898 468986 434134
rect 469222 433898 469404 434134
rect 468804 398454 469404 433898
rect 468804 398218 468986 398454
rect 469222 398218 469404 398454
rect 468804 398134 469404 398218
rect 468804 397898 468986 398134
rect 469222 397898 469404 398134
rect 468804 362454 469404 397898
rect 468804 362218 468986 362454
rect 469222 362218 469404 362454
rect 468804 362134 469404 362218
rect 468804 361898 468986 362134
rect 469222 361898 469404 362134
rect 468804 326454 469404 361898
rect 468804 326218 468986 326454
rect 469222 326218 469404 326454
rect 468804 326134 469404 326218
rect 468804 325898 468986 326134
rect 469222 325898 469404 326134
rect 468804 290454 469404 325898
rect 468804 290218 468986 290454
rect 469222 290218 469404 290454
rect 468804 290134 469404 290218
rect 468804 289898 468986 290134
rect 469222 289898 469404 290134
rect 468804 254454 469404 289898
rect 468804 254218 468986 254454
rect 469222 254218 469404 254454
rect 468804 254134 469404 254218
rect 468804 253898 468986 254134
rect 469222 253898 469404 254134
rect 468804 218454 469404 253898
rect 468804 218218 468986 218454
rect 469222 218218 469404 218454
rect 468804 218134 469404 218218
rect 468804 217898 468986 218134
rect 469222 217898 469404 218134
rect 468804 182454 469404 217898
rect 468804 182218 468986 182454
rect 469222 182218 469404 182454
rect 468804 182134 469404 182218
rect 468804 181898 468986 182134
rect 469222 181898 469404 182134
rect 468804 146454 469404 181898
rect 468804 146218 468986 146454
rect 469222 146218 469404 146454
rect 468804 146134 469404 146218
rect 468804 145898 468986 146134
rect 469222 145898 469404 146134
rect 468804 110454 469404 145898
rect 468804 110218 468986 110454
rect 469222 110218 469404 110454
rect 468804 110134 469404 110218
rect 468804 109898 468986 110134
rect 469222 109898 469404 110134
rect 468804 74454 469404 109898
rect 468804 74218 468986 74454
rect 469222 74218 469404 74454
rect 468804 74134 469404 74218
rect 468804 73898 468986 74134
rect 469222 73898 469404 74134
rect 468804 38454 469404 73898
rect 468804 38218 468986 38454
rect 469222 38218 469404 38454
rect 468804 38134 469404 38218
rect 468804 37898 468986 38134
rect 469222 37898 469404 38134
rect 462267 29476 462333 29477
rect 462267 29412 462268 29476
rect 462332 29412 462333 29476
rect 462267 29411 462333 29412
rect 462270 29205 462330 29411
rect 462267 29204 462333 29205
rect 462267 29140 462268 29204
rect 462332 29140 462333 29204
rect 462267 29139 462333 29140
rect 462267 17100 462333 17101
rect 462267 17036 462268 17100
rect 462332 17036 462333 17100
rect 462267 17035 462333 17036
rect 462270 16829 462330 17035
rect 462267 16828 462333 16829
rect 462267 16764 462268 16828
rect 462332 16764 462333 16828
rect 462267 16763 462333 16764
rect 468804 2454 469404 37898
rect 468804 2218 468986 2454
rect 469222 2218 469404 2454
rect 468804 2134 469404 2218
rect 468804 1898 468986 2134
rect 469222 1898 469404 2134
rect 468804 -346 469404 1898
rect 468804 -582 468986 -346
rect 469222 -582 469404 -346
rect 468804 -666 469404 -582
rect 468804 -902 468986 -666
rect 469222 -902 469404 -666
rect 468804 -1844 469404 -902
rect 472404 690054 473004 706122
rect 472404 689818 472586 690054
rect 472822 689818 473004 690054
rect 472404 689734 473004 689818
rect 472404 689498 472586 689734
rect 472822 689498 473004 689734
rect 472404 654054 473004 689498
rect 472404 653818 472586 654054
rect 472822 653818 473004 654054
rect 472404 653734 473004 653818
rect 472404 653498 472586 653734
rect 472822 653498 473004 653734
rect 472404 618054 473004 653498
rect 472404 617818 472586 618054
rect 472822 617818 473004 618054
rect 472404 617734 473004 617818
rect 472404 617498 472586 617734
rect 472822 617498 473004 617734
rect 472404 582054 473004 617498
rect 472404 581818 472586 582054
rect 472822 581818 473004 582054
rect 472404 581734 473004 581818
rect 472404 581498 472586 581734
rect 472822 581498 473004 581734
rect 472404 546054 473004 581498
rect 472404 545818 472586 546054
rect 472822 545818 473004 546054
rect 472404 545734 473004 545818
rect 472404 545498 472586 545734
rect 472822 545498 473004 545734
rect 472404 510054 473004 545498
rect 472404 509818 472586 510054
rect 472822 509818 473004 510054
rect 472404 509734 473004 509818
rect 472404 509498 472586 509734
rect 472822 509498 473004 509734
rect 472404 474054 473004 509498
rect 472404 473818 472586 474054
rect 472822 473818 473004 474054
rect 472404 473734 473004 473818
rect 472404 473498 472586 473734
rect 472822 473498 473004 473734
rect 472404 438054 473004 473498
rect 472404 437818 472586 438054
rect 472822 437818 473004 438054
rect 472404 437734 473004 437818
rect 472404 437498 472586 437734
rect 472822 437498 473004 437734
rect 472404 402054 473004 437498
rect 472404 401818 472586 402054
rect 472822 401818 473004 402054
rect 472404 401734 473004 401818
rect 472404 401498 472586 401734
rect 472822 401498 473004 401734
rect 472404 366054 473004 401498
rect 472404 365818 472586 366054
rect 472822 365818 473004 366054
rect 472404 365734 473004 365818
rect 472404 365498 472586 365734
rect 472822 365498 473004 365734
rect 472404 330054 473004 365498
rect 472404 329818 472586 330054
rect 472822 329818 473004 330054
rect 472404 329734 473004 329818
rect 472404 329498 472586 329734
rect 472822 329498 473004 329734
rect 472404 294054 473004 329498
rect 472404 293818 472586 294054
rect 472822 293818 473004 294054
rect 472404 293734 473004 293818
rect 472404 293498 472586 293734
rect 472822 293498 473004 293734
rect 472404 258054 473004 293498
rect 472404 257818 472586 258054
rect 472822 257818 473004 258054
rect 472404 257734 473004 257818
rect 472404 257498 472586 257734
rect 472822 257498 473004 257734
rect 472404 222054 473004 257498
rect 472404 221818 472586 222054
rect 472822 221818 473004 222054
rect 472404 221734 473004 221818
rect 472404 221498 472586 221734
rect 472822 221498 473004 221734
rect 472404 186054 473004 221498
rect 472404 185818 472586 186054
rect 472822 185818 473004 186054
rect 472404 185734 473004 185818
rect 472404 185498 472586 185734
rect 472822 185498 473004 185734
rect 472404 150054 473004 185498
rect 472404 149818 472586 150054
rect 472822 149818 473004 150054
rect 472404 149734 473004 149818
rect 472404 149498 472586 149734
rect 472822 149498 473004 149734
rect 472404 114054 473004 149498
rect 472404 113818 472586 114054
rect 472822 113818 473004 114054
rect 472404 113734 473004 113818
rect 472404 113498 472586 113734
rect 472822 113498 473004 113734
rect 472404 78054 473004 113498
rect 476004 693654 476604 707962
rect 476004 693418 476186 693654
rect 476422 693418 476604 693654
rect 476004 693334 476604 693418
rect 476004 693098 476186 693334
rect 476422 693098 476604 693334
rect 476004 657654 476604 693098
rect 476004 657418 476186 657654
rect 476422 657418 476604 657654
rect 476004 657334 476604 657418
rect 476004 657098 476186 657334
rect 476422 657098 476604 657334
rect 476004 621654 476604 657098
rect 476004 621418 476186 621654
rect 476422 621418 476604 621654
rect 476004 621334 476604 621418
rect 476004 621098 476186 621334
rect 476422 621098 476604 621334
rect 476004 585654 476604 621098
rect 476004 585418 476186 585654
rect 476422 585418 476604 585654
rect 476004 585334 476604 585418
rect 476004 585098 476186 585334
rect 476422 585098 476604 585334
rect 476004 549654 476604 585098
rect 476004 549418 476186 549654
rect 476422 549418 476604 549654
rect 476004 549334 476604 549418
rect 476004 549098 476186 549334
rect 476422 549098 476604 549334
rect 476004 513654 476604 549098
rect 476004 513418 476186 513654
rect 476422 513418 476604 513654
rect 476004 513334 476604 513418
rect 476004 513098 476186 513334
rect 476422 513098 476604 513334
rect 476004 477654 476604 513098
rect 476004 477418 476186 477654
rect 476422 477418 476604 477654
rect 476004 477334 476604 477418
rect 476004 477098 476186 477334
rect 476422 477098 476604 477334
rect 476004 441654 476604 477098
rect 476004 441418 476186 441654
rect 476422 441418 476604 441654
rect 476004 441334 476604 441418
rect 476004 441098 476186 441334
rect 476422 441098 476604 441334
rect 476004 405654 476604 441098
rect 476004 405418 476186 405654
rect 476422 405418 476604 405654
rect 476004 405334 476604 405418
rect 476004 405098 476186 405334
rect 476422 405098 476604 405334
rect 476004 369654 476604 405098
rect 476004 369418 476186 369654
rect 476422 369418 476604 369654
rect 476004 369334 476604 369418
rect 476004 369098 476186 369334
rect 476422 369098 476604 369334
rect 476004 333654 476604 369098
rect 476004 333418 476186 333654
rect 476422 333418 476604 333654
rect 476004 333334 476604 333418
rect 476004 333098 476186 333334
rect 476422 333098 476604 333334
rect 476004 297654 476604 333098
rect 476004 297418 476186 297654
rect 476422 297418 476604 297654
rect 476004 297334 476604 297418
rect 476004 297098 476186 297334
rect 476422 297098 476604 297334
rect 476004 261654 476604 297098
rect 476004 261418 476186 261654
rect 476422 261418 476604 261654
rect 476004 261334 476604 261418
rect 476004 261098 476186 261334
rect 476422 261098 476604 261334
rect 476004 225654 476604 261098
rect 476004 225418 476186 225654
rect 476422 225418 476604 225654
rect 476004 225334 476604 225418
rect 476004 225098 476186 225334
rect 476422 225098 476604 225334
rect 476004 189654 476604 225098
rect 476004 189418 476186 189654
rect 476422 189418 476604 189654
rect 476004 189334 476604 189418
rect 476004 189098 476186 189334
rect 476422 189098 476604 189334
rect 476004 153654 476604 189098
rect 476004 153418 476186 153654
rect 476422 153418 476604 153654
rect 476004 153334 476604 153418
rect 476004 153098 476186 153334
rect 476422 153098 476604 153334
rect 476004 117654 476604 153098
rect 476004 117418 476186 117654
rect 476422 117418 476604 117654
rect 476004 117334 476604 117418
rect 476004 117098 476186 117334
rect 476422 117098 476604 117334
rect 473307 87276 473373 87277
rect 473307 87212 473308 87276
rect 473372 87212 473373 87276
rect 473307 87211 473373 87212
rect 473310 87005 473370 87211
rect 473307 87004 473373 87005
rect 473307 86940 473308 87004
rect 473372 86940 473373 87004
rect 473307 86939 473373 86940
rect 472404 77818 472586 78054
rect 472822 77818 473004 78054
rect 472404 77734 473004 77818
rect 472404 77498 472586 77734
rect 472822 77498 473004 77734
rect 472404 42054 473004 77498
rect 472404 41818 472586 42054
rect 472822 41818 473004 42054
rect 472404 41734 473004 41818
rect 472404 41498 472586 41734
rect 472822 41498 473004 41734
rect 472404 6054 473004 41498
rect 472404 5818 472586 6054
rect 472822 5818 473004 6054
rect 472404 5734 473004 5818
rect 472404 5498 472586 5734
rect 472822 5498 473004 5734
rect 472404 -2186 473004 5498
rect 472404 -2422 472586 -2186
rect 472822 -2422 473004 -2186
rect 472404 -2506 473004 -2422
rect 472404 -2742 472586 -2506
rect 472822 -2742 473004 -2506
rect 472404 -3684 473004 -2742
rect 476004 81654 476604 117098
rect 476004 81418 476186 81654
rect 476422 81418 476604 81654
rect 476004 81334 476604 81418
rect 476004 81098 476186 81334
rect 476422 81098 476604 81334
rect 476004 45654 476604 81098
rect 476004 45418 476186 45654
rect 476422 45418 476604 45654
rect 476004 45334 476604 45418
rect 476004 45098 476186 45334
rect 476422 45098 476604 45334
rect 476004 9654 476604 45098
rect 476004 9418 476186 9654
rect 476422 9418 476604 9654
rect 476004 9334 476604 9418
rect 476004 9098 476186 9334
rect 476422 9098 476604 9334
rect 476004 -4026 476604 9098
rect 476004 -4262 476186 -4026
rect 476422 -4262 476604 -4026
rect 476004 -4346 476604 -4262
rect 476004 -4582 476186 -4346
rect 476422 -4582 476604 -4346
rect 476004 -5524 476604 -4582
rect 479604 697254 480204 709802
rect 497604 711278 498204 711300
rect 497604 711042 497786 711278
rect 498022 711042 498204 711278
rect 497604 710958 498204 711042
rect 497604 710722 497786 710958
rect 498022 710722 498204 710958
rect 494004 709438 494604 709460
rect 494004 709202 494186 709438
rect 494422 709202 494604 709438
rect 494004 709118 494604 709202
rect 494004 708882 494186 709118
rect 494422 708882 494604 709118
rect 490404 707598 491004 707620
rect 490404 707362 490586 707598
rect 490822 707362 491004 707598
rect 490404 707278 491004 707362
rect 490404 707042 490586 707278
rect 490822 707042 491004 707278
rect 479604 697018 479786 697254
rect 480022 697018 480204 697254
rect 479604 696934 480204 697018
rect 479604 696698 479786 696934
rect 480022 696698 480204 696934
rect 479604 661254 480204 696698
rect 479604 661018 479786 661254
rect 480022 661018 480204 661254
rect 479604 660934 480204 661018
rect 479604 660698 479786 660934
rect 480022 660698 480204 660934
rect 479604 625254 480204 660698
rect 479604 625018 479786 625254
rect 480022 625018 480204 625254
rect 479604 624934 480204 625018
rect 479604 624698 479786 624934
rect 480022 624698 480204 624934
rect 479604 589254 480204 624698
rect 479604 589018 479786 589254
rect 480022 589018 480204 589254
rect 479604 588934 480204 589018
rect 479604 588698 479786 588934
rect 480022 588698 480204 588934
rect 479604 553254 480204 588698
rect 479604 553018 479786 553254
rect 480022 553018 480204 553254
rect 479604 552934 480204 553018
rect 479604 552698 479786 552934
rect 480022 552698 480204 552934
rect 479604 517254 480204 552698
rect 479604 517018 479786 517254
rect 480022 517018 480204 517254
rect 479604 516934 480204 517018
rect 479604 516698 479786 516934
rect 480022 516698 480204 516934
rect 479604 481254 480204 516698
rect 479604 481018 479786 481254
rect 480022 481018 480204 481254
rect 479604 480934 480204 481018
rect 479604 480698 479786 480934
rect 480022 480698 480204 480934
rect 479604 445254 480204 480698
rect 479604 445018 479786 445254
rect 480022 445018 480204 445254
rect 479604 444934 480204 445018
rect 479604 444698 479786 444934
rect 480022 444698 480204 444934
rect 479604 409254 480204 444698
rect 479604 409018 479786 409254
rect 480022 409018 480204 409254
rect 479604 408934 480204 409018
rect 479604 408698 479786 408934
rect 480022 408698 480204 408934
rect 479604 373254 480204 408698
rect 479604 373018 479786 373254
rect 480022 373018 480204 373254
rect 479604 372934 480204 373018
rect 479604 372698 479786 372934
rect 480022 372698 480204 372934
rect 479604 337254 480204 372698
rect 479604 337018 479786 337254
rect 480022 337018 480204 337254
rect 479604 336934 480204 337018
rect 479604 336698 479786 336934
rect 480022 336698 480204 336934
rect 479604 301254 480204 336698
rect 479604 301018 479786 301254
rect 480022 301018 480204 301254
rect 479604 300934 480204 301018
rect 479604 300698 479786 300934
rect 480022 300698 480204 300934
rect 479604 265254 480204 300698
rect 479604 265018 479786 265254
rect 480022 265018 480204 265254
rect 479604 264934 480204 265018
rect 479604 264698 479786 264934
rect 480022 264698 480204 264934
rect 479604 229254 480204 264698
rect 479604 229018 479786 229254
rect 480022 229018 480204 229254
rect 479604 228934 480204 229018
rect 479604 228698 479786 228934
rect 480022 228698 480204 228934
rect 479604 193254 480204 228698
rect 479604 193018 479786 193254
rect 480022 193018 480204 193254
rect 479604 192934 480204 193018
rect 479604 192698 479786 192934
rect 480022 192698 480204 192934
rect 479604 157254 480204 192698
rect 479604 157018 479786 157254
rect 480022 157018 480204 157254
rect 479604 156934 480204 157018
rect 479604 156698 479786 156934
rect 480022 156698 480204 156934
rect 479604 121254 480204 156698
rect 479604 121018 479786 121254
rect 480022 121018 480204 121254
rect 479604 120934 480204 121018
rect 479604 120698 479786 120934
rect 480022 120698 480204 120934
rect 479604 85254 480204 120698
rect 479604 85018 479786 85254
rect 480022 85018 480204 85254
rect 479604 84934 480204 85018
rect 479604 84698 479786 84934
rect 480022 84698 480204 84934
rect 479604 49254 480204 84698
rect 479604 49018 479786 49254
rect 480022 49018 480204 49254
rect 479604 48934 480204 49018
rect 479604 48698 479786 48934
rect 480022 48698 480204 48934
rect 479604 13254 480204 48698
rect 479604 13018 479786 13254
rect 480022 13018 480204 13254
rect 479604 12934 480204 13018
rect 479604 12698 479786 12934
rect 480022 12698 480204 12934
rect 461604 -7022 461786 -6786
rect 462022 -7022 462204 -6786
rect 461604 -7106 462204 -7022
rect 461604 -7342 461786 -7106
rect 462022 -7342 462204 -7106
rect 461604 -7364 462204 -7342
rect 479604 -5866 480204 12698
rect 486804 705758 487404 705780
rect 486804 705522 486986 705758
rect 487222 705522 487404 705758
rect 486804 705438 487404 705522
rect 486804 705202 486986 705438
rect 487222 705202 487404 705438
rect 486804 668454 487404 705202
rect 486804 668218 486986 668454
rect 487222 668218 487404 668454
rect 486804 668134 487404 668218
rect 486804 667898 486986 668134
rect 487222 667898 487404 668134
rect 486804 632454 487404 667898
rect 486804 632218 486986 632454
rect 487222 632218 487404 632454
rect 486804 632134 487404 632218
rect 486804 631898 486986 632134
rect 487222 631898 487404 632134
rect 486804 596454 487404 631898
rect 486804 596218 486986 596454
rect 487222 596218 487404 596454
rect 486804 596134 487404 596218
rect 486804 595898 486986 596134
rect 487222 595898 487404 596134
rect 486804 560454 487404 595898
rect 486804 560218 486986 560454
rect 487222 560218 487404 560454
rect 486804 560134 487404 560218
rect 486804 559898 486986 560134
rect 487222 559898 487404 560134
rect 486804 524454 487404 559898
rect 486804 524218 486986 524454
rect 487222 524218 487404 524454
rect 486804 524134 487404 524218
rect 486804 523898 486986 524134
rect 487222 523898 487404 524134
rect 486804 488454 487404 523898
rect 486804 488218 486986 488454
rect 487222 488218 487404 488454
rect 486804 488134 487404 488218
rect 486804 487898 486986 488134
rect 487222 487898 487404 488134
rect 486804 452454 487404 487898
rect 486804 452218 486986 452454
rect 487222 452218 487404 452454
rect 486804 452134 487404 452218
rect 486804 451898 486986 452134
rect 487222 451898 487404 452134
rect 486804 416454 487404 451898
rect 486804 416218 486986 416454
rect 487222 416218 487404 416454
rect 486804 416134 487404 416218
rect 486804 415898 486986 416134
rect 487222 415898 487404 416134
rect 486804 380454 487404 415898
rect 486804 380218 486986 380454
rect 487222 380218 487404 380454
rect 486804 380134 487404 380218
rect 486804 379898 486986 380134
rect 487222 379898 487404 380134
rect 486804 344454 487404 379898
rect 486804 344218 486986 344454
rect 487222 344218 487404 344454
rect 486804 344134 487404 344218
rect 486804 343898 486986 344134
rect 487222 343898 487404 344134
rect 486804 308454 487404 343898
rect 486804 308218 486986 308454
rect 487222 308218 487404 308454
rect 486804 308134 487404 308218
rect 486804 307898 486986 308134
rect 487222 307898 487404 308134
rect 486804 272454 487404 307898
rect 486804 272218 486986 272454
rect 487222 272218 487404 272454
rect 486804 272134 487404 272218
rect 486804 271898 486986 272134
rect 487222 271898 487404 272134
rect 486804 236454 487404 271898
rect 486804 236218 486986 236454
rect 487222 236218 487404 236454
rect 486804 236134 487404 236218
rect 486804 235898 486986 236134
rect 487222 235898 487404 236134
rect 486804 200454 487404 235898
rect 486804 200218 486986 200454
rect 487222 200218 487404 200454
rect 486804 200134 487404 200218
rect 486804 199898 486986 200134
rect 487222 199898 487404 200134
rect 486804 164454 487404 199898
rect 486804 164218 486986 164454
rect 487222 164218 487404 164454
rect 486804 164134 487404 164218
rect 486804 163898 486986 164134
rect 487222 163898 487404 164134
rect 486804 128454 487404 163898
rect 486804 128218 486986 128454
rect 487222 128218 487404 128454
rect 486804 128134 487404 128218
rect 486804 127898 486986 128134
rect 487222 127898 487404 128134
rect 486804 92454 487404 127898
rect 486804 92218 486986 92454
rect 487222 92218 487404 92454
rect 486804 92134 487404 92218
rect 486804 91898 486986 92134
rect 487222 91898 487404 92134
rect 486804 56454 487404 91898
rect 486804 56218 486986 56454
rect 487222 56218 487404 56454
rect 486804 56134 487404 56218
rect 486804 55898 486986 56134
rect 487222 55898 487404 56134
rect 486804 20454 487404 55898
rect 486804 20218 486986 20454
rect 487222 20218 487404 20454
rect 486804 20134 487404 20218
rect 486804 19898 486986 20134
rect 487222 19898 487404 20134
rect 486804 -1266 487404 19898
rect 486804 -1502 486986 -1266
rect 487222 -1502 487404 -1266
rect 486804 -1586 487404 -1502
rect 486804 -1822 486986 -1586
rect 487222 -1822 487404 -1586
rect 486804 -1844 487404 -1822
rect 490404 672054 491004 707042
rect 490404 671818 490586 672054
rect 490822 671818 491004 672054
rect 490404 671734 491004 671818
rect 490404 671498 490586 671734
rect 490822 671498 491004 671734
rect 490404 636054 491004 671498
rect 490404 635818 490586 636054
rect 490822 635818 491004 636054
rect 490404 635734 491004 635818
rect 490404 635498 490586 635734
rect 490822 635498 491004 635734
rect 490404 600054 491004 635498
rect 490404 599818 490586 600054
rect 490822 599818 491004 600054
rect 490404 599734 491004 599818
rect 490404 599498 490586 599734
rect 490822 599498 491004 599734
rect 490404 564054 491004 599498
rect 490404 563818 490586 564054
rect 490822 563818 491004 564054
rect 490404 563734 491004 563818
rect 490404 563498 490586 563734
rect 490822 563498 491004 563734
rect 490404 528054 491004 563498
rect 490404 527818 490586 528054
rect 490822 527818 491004 528054
rect 490404 527734 491004 527818
rect 490404 527498 490586 527734
rect 490822 527498 491004 527734
rect 490404 492054 491004 527498
rect 490404 491818 490586 492054
rect 490822 491818 491004 492054
rect 490404 491734 491004 491818
rect 490404 491498 490586 491734
rect 490822 491498 491004 491734
rect 490404 456054 491004 491498
rect 490404 455818 490586 456054
rect 490822 455818 491004 456054
rect 490404 455734 491004 455818
rect 490404 455498 490586 455734
rect 490822 455498 491004 455734
rect 490404 420054 491004 455498
rect 490404 419818 490586 420054
rect 490822 419818 491004 420054
rect 490404 419734 491004 419818
rect 490404 419498 490586 419734
rect 490822 419498 491004 419734
rect 490404 384054 491004 419498
rect 490404 383818 490586 384054
rect 490822 383818 491004 384054
rect 490404 383734 491004 383818
rect 490404 383498 490586 383734
rect 490822 383498 491004 383734
rect 490404 348054 491004 383498
rect 490404 347818 490586 348054
rect 490822 347818 491004 348054
rect 490404 347734 491004 347818
rect 490404 347498 490586 347734
rect 490822 347498 491004 347734
rect 490404 312054 491004 347498
rect 490404 311818 490586 312054
rect 490822 311818 491004 312054
rect 490404 311734 491004 311818
rect 490404 311498 490586 311734
rect 490822 311498 491004 311734
rect 490404 276054 491004 311498
rect 490404 275818 490586 276054
rect 490822 275818 491004 276054
rect 490404 275734 491004 275818
rect 490404 275498 490586 275734
rect 490822 275498 491004 275734
rect 490404 240054 491004 275498
rect 490404 239818 490586 240054
rect 490822 239818 491004 240054
rect 490404 239734 491004 239818
rect 490404 239498 490586 239734
rect 490822 239498 491004 239734
rect 490404 204054 491004 239498
rect 490404 203818 490586 204054
rect 490822 203818 491004 204054
rect 490404 203734 491004 203818
rect 490404 203498 490586 203734
rect 490822 203498 491004 203734
rect 490404 168054 491004 203498
rect 490404 167818 490586 168054
rect 490822 167818 491004 168054
rect 490404 167734 491004 167818
rect 490404 167498 490586 167734
rect 490822 167498 491004 167734
rect 490404 132054 491004 167498
rect 490404 131818 490586 132054
rect 490822 131818 491004 132054
rect 490404 131734 491004 131818
rect 490404 131498 490586 131734
rect 490822 131498 491004 131734
rect 490404 96054 491004 131498
rect 490404 95818 490586 96054
rect 490822 95818 491004 96054
rect 490404 95734 491004 95818
rect 490404 95498 490586 95734
rect 490822 95498 491004 95734
rect 490404 60054 491004 95498
rect 490404 59818 490586 60054
rect 490822 59818 491004 60054
rect 490404 59734 491004 59818
rect 490404 59498 490586 59734
rect 490822 59498 491004 59734
rect 490404 24054 491004 59498
rect 490404 23818 490586 24054
rect 490822 23818 491004 24054
rect 490404 23734 491004 23818
rect 490404 23498 490586 23734
rect 490822 23498 491004 23734
rect 490404 -3106 491004 23498
rect 490404 -3342 490586 -3106
rect 490822 -3342 491004 -3106
rect 490404 -3426 491004 -3342
rect 490404 -3662 490586 -3426
rect 490822 -3662 491004 -3426
rect 490404 -3684 491004 -3662
rect 494004 675654 494604 708882
rect 494004 675418 494186 675654
rect 494422 675418 494604 675654
rect 494004 675334 494604 675418
rect 494004 675098 494186 675334
rect 494422 675098 494604 675334
rect 494004 639654 494604 675098
rect 494004 639418 494186 639654
rect 494422 639418 494604 639654
rect 494004 639334 494604 639418
rect 494004 639098 494186 639334
rect 494422 639098 494604 639334
rect 494004 603654 494604 639098
rect 494004 603418 494186 603654
rect 494422 603418 494604 603654
rect 494004 603334 494604 603418
rect 494004 603098 494186 603334
rect 494422 603098 494604 603334
rect 494004 567654 494604 603098
rect 494004 567418 494186 567654
rect 494422 567418 494604 567654
rect 494004 567334 494604 567418
rect 494004 567098 494186 567334
rect 494422 567098 494604 567334
rect 494004 531654 494604 567098
rect 494004 531418 494186 531654
rect 494422 531418 494604 531654
rect 494004 531334 494604 531418
rect 494004 531098 494186 531334
rect 494422 531098 494604 531334
rect 494004 495654 494604 531098
rect 494004 495418 494186 495654
rect 494422 495418 494604 495654
rect 494004 495334 494604 495418
rect 494004 495098 494186 495334
rect 494422 495098 494604 495334
rect 494004 459654 494604 495098
rect 494004 459418 494186 459654
rect 494422 459418 494604 459654
rect 494004 459334 494604 459418
rect 494004 459098 494186 459334
rect 494422 459098 494604 459334
rect 494004 423654 494604 459098
rect 494004 423418 494186 423654
rect 494422 423418 494604 423654
rect 494004 423334 494604 423418
rect 494004 423098 494186 423334
rect 494422 423098 494604 423334
rect 494004 387654 494604 423098
rect 494004 387418 494186 387654
rect 494422 387418 494604 387654
rect 494004 387334 494604 387418
rect 494004 387098 494186 387334
rect 494422 387098 494604 387334
rect 494004 351654 494604 387098
rect 494004 351418 494186 351654
rect 494422 351418 494604 351654
rect 494004 351334 494604 351418
rect 494004 351098 494186 351334
rect 494422 351098 494604 351334
rect 494004 315654 494604 351098
rect 494004 315418 494186 315654
rect 494422 315418 494604 315654
rect 494004 315334 494604 315418
rect 494004 315098 494186 315334
rect 494422 315098 494604 315334
rect 494004 279654 494604 315098
rect 494004 279418 494186 279654
rect 494422 279418 494604 279654
rect 494004 279334 494604 279418
rect 494004 279098 494186 279334
rect 494422 279098 494604 279334
rect 494004 243654 494604 279098
rect 494004 243418 494186 243654
rect 494422 243418 494604 243654
rect 494004 243334 494604 243418
rect 494004 243098 494186 243334
rect 494422 243098 494604 243334
rect 494004 207654 494604 243098
rect 494004 207418 494186 207654
rect 494422 207418 494604 207654
rect 494004 207334 494604 207418
rect 494004 207098 494186 207334
rect 494422 207098 494604 207334
rect 494004 171654 494604 207098
rect 494004 171418 494186 171654
rect 494422 171418 494604 171654
rect 494004 171334 494604 171418
rect 494004 171098 494186 171334
rect 494422 171098 494604 171334
rect 494004 135654 494604 171098
rect 494004 135418 494186 135654
rect 494422 135418 494604 135654
rect 494004 135334 494604 135418
rect 494004 135098 494186 135334
rect 494422 135098 494604 135334
rect 494004 99654 494604 135098
rect 494004 99418 494186 99654
rect 494422 99418 494604 99654
rect 494004 99334 494604 99418
rect 494004 99098 494186 99334
rect 494422 99098 494604 99334
rect 494004 63654 494604 99098
rect 494004 63418 494186 63654
rect 494422 63418 494604 63654
rect 494004 63334 494604 63418
rect 494004 63098 494186 63334
rect 494422 63098 494604 63334
rect 494004 27654 494604 63098
rect 494004 27418 494186 27654
rect 494422 27418 494604 27654
rect 494004 27334 494604 27418
rect 494004 27098 494186 27334
rect 494422 27098 494604 27334
rect 494004 -4946 494604 27098
rect 494004 -5182 494186 -4946
rect 494422 -5182 494604 -4946
rect 494004 -5266 494604 -5182
rect 494004 -5502 494186 -5266
rect 494422 -5502 494604 -5266
rect 494004 -5524 494604 -5502
rect 497604 679254 498204 710722
rect 515604 710358 516204 711300
rect 515604 710122 515786 710358
rect 516022 710122 516204 710358
rect 515604 710038 516204 710122
rect 515604 709802 515786 710038
rect 516022 709802 516204 710038
rect 512004 708518 512604 709460
rect 512004 708282 512186 708518
rect 512422 708282 512604 708518
rect 512004 708198 512604 708282
rect 512004 707962 512186 708198
rect 512422 707962 512604 708198
rect 508404 706678 509004 707620
rect 508404 706442 508586 706678
rect 508822 706442 509004 706678
rect 508404 706358 509004 706442
rect 508404 706122 508586 706358
rect 508822 706122 509004 706358
rect 497604 679018 497786 679254
rect 498022 679018 498204 679254
rect 497604 678934 498204 679018
rect 497604 678698 497786 678934
rect 498022 678698 498204 678934
rect 497604 643254 498204 678698
rect 497604 643018 497786 643254
rect 498022 643018 498204 643254
rect 497604 642934 498204 643018
rect 497604 642698 497786 642934
rect 498022 642698 498204 642934
rect 497604 607254 498204 642698
rect 497604 607018 497786 607254
rect 498022 607018 498204 607254
rect 497604 606934 498204 607018
rect 497604 606698 497786 606934
rect 498022 606698 498204 606934
rect 497604 571254 498204 606698
rect 497604 571018 497786 571254
rect 498022 571018 498204 571254
rect 497604 570934 498204 571018
rect 497604 570698 497786 570934
rect 498022 570698 498204 570934
rect 497604 535254 498204 570698
rect 497604 535018 497786 535254
rect 498022 535018 498204 535254
rect 497604 534934 498204 535018
rect 497604 534698 497786 534934
rect 498022 534698 498204 534934
rect 497604 499254 498204 534698
rect 497604 499018 497786 499254
rect 498022 499018 498204 499254
rect 497604 498934 498204 499018
rect 497604 498698 497786 498934
rect 498022 498698 498204 498934
rect 497604 463254 498204 498698
rect 497604 463018 497786 463254
rect 498022 463018 498204 463254
rect 497604 462934 498204 463018
rect 497604 462698 497786 462934
rect 498022 462698 498204 462934
rect 497604 427254 498204 462698
rect 497604 427018 497786 427254
rect 498022 427018 498204 427254
rect 497604 426934 498204 427018
rect 497604 426698 497786 426934
rect 498022 426698 498204 426934
rect 497604 391254 498204 426698
rect 497604 391018 497786 391254
rect 498022 391018 498204 391254
rect 497604 390934 498204 391018
rect 497604 390698 497786 390934
rect 498022 390698 498204 390934
rect 497604 355254 498204 390698
rect 497604 355018 497786 355254
rect 498022 355018 498204 355254
rect 497604 354934 498204 355018
rect 497604 354698 497786 354934
rect 498022 354698 498204 354934
rect 497604 319254 498204 354698
rect 497604 319018 497786 319254
rect 498022 319018 498204 319254
rect 497604 318934 498204 319018
rect 497604 318698 497786 318934
rect 498022 318698 498204 318934
rect 497604 283254 498204 318698
rect 497604 283018 497786 283254
rect 498022 283018 498204 283254
rect 497604 282934 498204 283018
rect 497604 282698 497786 282934
rect 498022 282698 498204 282934
rect 497604 247254 498204 282698
rect 497604 247018 497786 247254
rect 498022 247018 498204 247254
rect 497604 246934 498204 247018
rect 497604 246698 497786 246934
rect 498022 246698 498204 246934
rect 497604 211254 498204 246698
rect 497604 211018 497786 211254
rect 498022 211018 498204 211254
rect 497604 210934 498204 211018
rect 497604 210698 497786 210934
rect 498022 210698 498204 210934
rect 497604 175254 498204 210698
rect 497604 175018 497786 175254
rect 498022 175018 498204 175254
rect 497604 174934 498204 175018
rect 497604 174698 497786 174934
rect 498022 174698 498204 174934
rect 497604 139254 498204 174698
rect 497604 139018 497786 139254
rect 498022 139018 498204 139254
rect 497604 138934 498204 139018
rect 497604 138698 497786 138934
rect 498022 138698 498204 138934
rect 497604 103254 498204 138698
rect 497604 103018 497786 103254
rect 498022 103018 498204 103254
rect 497604 102934 498204 103018
rect 497604 102698 497786 102934
rect 498022 102698 498204 102934
rect 497604 67254 498204 102698
rect 497604 67018 497786 67254
rect 498022 67018 498204 67254
rect 497604 66934 498204 67018
rect 497604 66698 497786 66934
rect 498022 66698 498204 66934
rect 497604 31254 498204 66698
rect 497604 31018 497786 31254
rect 498022 31018 498204 31254
rect 497604 30934 498204 31018
rect 497604 30698 497786 30934
rect 498022 30698 498204 30934
rect 479604 -6102 479786 -5866
rect 480022 -6102 480204 -5866
rect 479604 -6186 480204 -6102
rect 479604 -6422 479786 -6186
rect 480022 -6422 480204 -6186
rect 479604 -7364 480204 -6422
rect 497604 -6786 498204 30698
rect 504804 704838 505404 705780
rect 504804 704602 504986 704838
rect 505222 704602 505404 704838
rect 504804 704518 505404 704602
rect 504804 704282 504986 704518
rect 505222 704282 505404 704518
rect 504804 686454 505404 704282
rect 504804 686218 504986 686454
rect 505222 686218 505404 686454
rect 504804 686134 505404 686218
rect 504804 685898 504986 686134
rect 505222 685898 505404 686134
rect 504804 650454 505404 685898
rect 504804 650218 504986 650454
rect 505222 650218 505404 650454
rect 504804 650134 505404 650218
rect 504804 649898 504986 650134
rect 505222 649898 505404 650134
rect 504804 614454 505404 649898
rect 504804 614218 504986 614454
rect 505222 614218 505404 614454
rect 504804 614134 505404 614218
rect 504804 613898 504986 614134
rect 505222 613898 505404 614134
rect 504804 578454 505404 613898
rect 504804 578218 504986 578454
rect 505222 578218 505404 578454
rect 504804 578134 505404 578218
rect 504804 577898 504986 578134
rect 505222 577898 505404 578134
rect 504804 542454 505404 577898
rect 504804 542218 504986 542454
rect 505222 542218 505404 542454
rect 504804 542134 505404 542218
rect 504804 541898 504986 542134
rect 505222 541898 505404 542134
rect 504804 506454 505404 541898
rect 504804 506218 504986 506454
rect 505222 506218 505404 506454
rect 504804 506134 505404 506218
rect 504804 505898 504986 506134
rect 505222 505898 505404 506134
rect 504804 470454 505404 505898
rect 504804 470218 504986 470454
rect 505222 470218 505404 470454
rect 504804 470134 505404 470218
rect 504804 469898 504986 470134
rect 505222 469898 505404 470134
rect 504804 434454 505404 469898
rect 504804 434218 504986 434454
rect 505222 434218 505404 434454
rect 504804 434134 505404 434218
rect 504804 433898 504986 434134
rect 505222 433898 505404 434134
rect 504804 398454 505404 433898
rect 504804 398218 504986 398454
rect 505222 398218 505404 398454
rect 504804 398134 505404 398218
rect 504804 397898 504986 398134
rect 505222 397898 505404 398134
rect 504804 362454 505404 397898
rect 504804 362218 504986 362454
rect 505222 362218 505404 362454
rect 504804 362134 505404 362218
rect 504804 361898 504986 362134
rect 505222 361898 505404 362134
rect 504804 326454 505404 361898
rect 504804 326218 504986 326454
rect 505222 326218 505404 326454
rect 504804 326134 505404 326218
rect 504804 325898 504986 326134
rect 505222 325898 505404 326134
rect 504804 290454 505404 325898
rect 504804 290218 504986 290454
rect 505222 290218 505404 290454
rect 504804 290134 505404 290218
rect 504804 289898 504986 290134
rect 505222 289898 505404 290134
rect 504804 254454 505404 289898
rect 504804 254218 504986 254454
rect 505222 254218 505404 254454
rect 504804 254134 505404 254218
rect 504804 253898 504986 254134
rect 505222 253898 505404 254134
rect 504804 218454 505404 253898
rect 504804 218218 504986 218454
rect 505222 218218 505404 218454
rect 504804 218134 505404 218218
rect 504804 217898 504986 218134
rect 505222 217898 505404 218134
rect 504804 182454 505404 217898
rect 504804 182218 504986 182454
rect 505222 182218 505404 182454
rect 504804 182134 505404 182218
rect 504804 181898 504986 182134
rect 505222 181898 505404 182134
rect 504804 146454 505404 181898
rect 504804 146218 504986 146454
rect 505222 146218 505404 146454
rect 504804 146134 505404 146218
rect 504804 145898 504986 146134
rect 505222 145898 505404 146134
rect 504804 110454 505404 145898
rect 504804 110218 504986 110454
rect 505222 110218 505404 110454
rect 504804 110134 505404 110218
rect 504804 109898 504986 110134
rect 505222 109898 505404 110134
rect 504804 74454 505404 109898
rect 504804 74218 504986 74454
rect 505222 74218 505404 74454
rect 504804 74134 505404 74218
rect 504804 73898 504986 74134
rect 505222 73898 505404 74134
rect 504804 38454 505404 73898
rect 504804 38218 504986 38454
rect 505222 38218 505404 38454
rect 504804 38134 505404 38218
rect 504804 37898 504986 38134
rect 505222 37898 505404 38134
rect 504804 2454 505404 37898
rect 504804 2218 504986 2454
rect 505222 2218 505404 2454
rect 504804 2134 505404 2218
rect 504804 1898 504986 2134
rect 505222 1898 505404 2134
rect 504804 -346 505404 1898
rect 504804 -582 504986 -346
rect 505222 -582 505404 -346
rect 504804 -666 505404 -582
rect 504804 -902 504986 -666
rect 505222 -902 505404 -666
rect 504804 -1844 505404 -902
rect 508404 690054 509004 706122
rect 508404 689818 508586 690054
rect 508822 689818 509004 690054
rect 508404 689734 509004 689818
rect 508404 689498 508586 689734
rect 508822 689498 509004 689734
rect 508404 654054 509004 689498
rect 508404 653818 508586 654054
rect 508822 653818 509004 654054
rect 508404 653734 509004 653818
rect 508404 653498 508586 653734
rect 508822 653498 509004 653734
rect 508404 618054 509004 653498
rect 508404 617818 508586 618054
rect 508822 617818 509004 618054
rect 508404 617734 509004 617818
rect 508404 617498 508586 617734
rect 508822 617498 509004 617734
rect 508404 582054 509004 617498
rect 508404 581818 508586 582054
rect 508822 581818 509004 582054
rect 508404 581734 509004 581818
rect 508404 581498 508586 581734
rect 508822 581498 509004 581734
rect 508404 546054 509004 581498
rect 508404 545818 508586 546054
rect 508822 545818 509004 546054
rect 508404 545734 509004 545818
rect 508404 545498 508586 545734
rect 508822 545498 509004 545734
rect 508404 510054 509004 545498
rect 508404 509818 508586 510054
rect 508822 509818 509004 510054
rect 508404 509734 509004 509818
rect 508404 509498 508586 509734
rect 508822 509498 509004 509734
rect 508404 474054 509004 509498
rect 508404 473818 508586 474054
rect 508822 473818 509004 474054
rect 508404 473734 509004 473818
rect 508404 473498 508586 473734
rect 508822 473498 509004 473734
rect 508404 438054 509004 473498
rect 508404 437818 508586 438054
rect 508822 437818 509004 438054
rect 508404 437734 509004 437818
rect 508404 437498 508586 437734
rect 508822 437498 509004 437734
rect 508404 402054 509004 437498
rect 508404 401818 508586 402054
rect 508822 401818 509004 402054
rect 508404 401734 509004 401818
rect 508404 401498 508586 401734
rect 508822 401498 509004 401734
rect 508404 366054 509004 401498
rect 508404 365818 508586 366054
rect 508822 365818 509004 366054
rect 508404 365734 509004 365818
rect 508404 365498 508586 365734
rect 508822 365498 509004 365734
rect 508404 330054 509004 365498
rect 508404 329818 508586 330054
rect 508822 329818 509004 330054
rect 508404 329734 509004 329818
rect 508404 329498 508586 329734
rect 508822 329498 509004 329734
rect 508404 294054 509004 329498
rect 508404 293818 508586 294054
rect 508822 293818 509004 294054
rect 508404 293734 509004 293818
rect 508404 293498 508586 293734
rect 508822 293498 509004 293734
rect 508404 258054 509004 293498
rect 508404 257818 508586 258054
rect 508822 257818 509004 258054
rect 508404 257734 509004 257818
rect 508404 257498 508586 257734
rect 508822 257498 509004 257734
rect 508404 222054 509004 257498
rect 508404 221818 508586 222054
rect 508822 221818 509004 222054
rect 508404 221734 509004 221818
rect 508404 221498 508586 221734
rect 508822 221498 509004 221734
rect 508404 186054 509004 221498
rect 508404 185818 508586 186054
rect 508822 185818 509004 186054
rect 508404 185734 509004 185818
rect 508404 185498 508586 185734
rect 508822 185498 509004 185734
rect 508404 150054 509004 185498
rect 508404 149818 508586 150054
rect 508822 149818 509004 150054
rect 508404 149734 509004 149818
rect 508404 149498 508586 149734
rect 508822 149498 509004 149734
rect 508404 114054 509004 149498
rect 508404 113818 508586 114054
rect 508822 113818 509004 114054
rect 508404 113734 509004 113818
rect 508404 113498 508586 113734
rect 508822 113498 509004 113734
rect 508404 78054 509004 113498
rect 508404 77818 508586 78054
rect 508822 77818 509004 78054
rect 508404 77734 509004 77818
rect 508404 77498 508586 77734
rect 508822 77498 509004 77734
rect 508404 42054 509004 77498
rect 508404 41818 508586 42054
rect 508822 41818 509004 42054
rect 508404 41734 509004 41818
rect 508404 41498 508586 41734
rect 508822 41498 509004 41734
rect 508404 6054 509004 41498
rect 508404 5818 508586 6054
rect 508822 5818 509004 6054
rect 508404 5734 509004 5818
rect 508404 5498 508586 5734
rect 508822 5498 509004 5734
rect 508404 -2186 509004 5498
rect 508404 -2422 508586 -2186
rect 508822 -2422 509004 -2186
rect 508404 -2506 509004 -2422
rect 508404 -2742 508586 -2506
rect 508822 -2742 509004 -2506
rect 508404 -3684 509004 -2742
rect 512004 693654 512604 707962
rect 512004 693418 512186 693654
rect 512422 693418 512604 693654
rect 512004 693334 512604 693418
rect 512004 693098 512186 693334
rect 512422 693098 512604 693334
rect 512004 657654 512604 693098
rect 512004 657418 512186 657654
rect 512422 657418 512604 657654
rect 512004 657334 512604 657418
rect 512004 657098 512186 657334
rect 512422 657098 512604 657334
rect 512004 621654 512604 657098
rect 512004 621418 512186 621654
rect 512422 621418 512604 621654
rect 512004 621334 512604 621418
rect 512004 621098 512186 621334
rect 512422 621098 512604 621334
rect 512004 585654 512604 621098
rect 512004 585418 512186 585654
rect 512422 585418 512604 585654
rect 512004 585334 512604 585418
rect 512004 585098 512186 585334
rect 512422 585098 512604 585334
rect 512004 549654 512604 585098
rect 512004 549418 512186 549654
rect 512422 549418 512604 549654
rect 512004 549334 512604 549418
rect 512004 549098 512186 549334
rect 512422 549098 512604 549334
rect 512004 513654 512604 549098
rect 512004 513418 512186 513654
rect 512422 513418 512604 513654
rect 512004 513334 512604 513418
rect 512004 513098 512186 513334
rect 512422 513098 512604 513334
rect 512004 477654 512604 513098
rect 512004 477418 512186 477654
rect 512422 477418 512604 477654
rect 512004 477334 512604 477418
rect 512004 477098 512186 477334
rect 512422 477098 512604 477334
rect 512004 441654 512604 477098
rect 512004 441418 512186 441654
rect 512422 441418 512604 441654
rect 512004 441334 512604 441418
rect 512004 441098 512186 441334
rect 512422 441098 512604 441334
rect 512004 405654 512604 441098
rect 512004 405418 512186 405654
rect 512422 405418 512604 405654
rect 512004 405334 512604 405418
rect 512004 405098 512186 405334
rect 512422 405098 512604 405334
rect 512004 369654 512604 405098
rect 512004 369418 512186 369654
rect 512422 369418 512604 369654
rect 512004 369334 512604 369418
rect 512004 369098 512186 369334
rect 512422 369098 512604 369334
rect 512004 333654 512604 369098
rect 512004 333418 512186 333654
rect 512422 333418 512604 333654
rect 512004 333334 512604 333418
rect 512004 333098 512186 333334
rect 512422 333098 512604 333334
rect 512004 297654 512604 333098
rect 512004 297418 512186 297654
rect 512422 297418 512604 297654
rect 512004 297334 512604 297418
rect 512004 297098 512186 297334
rect 512422 297098 512604 297334
rect 512004 261654 512604 297098
rect 512004 261418 512186 261654
rect 512422 261418 512604 261654
rect 512004 261334 512604 261418
rect 512004 261098 512186 261334
rect 512422 261098 512604 261334
rect 512004 225654 512604 261098
rect 512004 225418 512186 225654
rect 512422 225418 512604 225654
rect 512004 225334 512604 225418
rect 512004 225098 512186 225334
rect 512422 225098 512604 225334
rect 512004 189654 512604 225098
rect 512004 189418 512186 189654
rect 512422 189418 512604 189654
rect 512004 189334 512604 189418
rect 512004 189098 512186 189334
rect 512422 189098 512604 189334
rect 512004 153654 512604 189098
rect 512004 153418 512186 153654
rect 512422 153418 512604 153654
rect 512004 153334 512604 153418
rect 512004 153098 512186 153334
rect 512422 153098 512604 153334
rect 512004 117654 512604 153098
rect 512004 117418 512186 117654
rect 512422 117418 512604 117654
rect 512004 117334 512604 117418
rect 512004 117098 512186 117334
rect 512422 117098 512604 117334
rect 512004 81654 512604 117098
rect 512004 81418 512186 81654
rect 512422 81418 512604 81654
rect 512004 81334 512604 81418
rect 512004 81098 512186 81334
rect 512422 81098 512604 81334
rect 512004 45654 512604 81098
rect 512004 45418 512186 45654
rect 512422 45418 512604 45654
rect 512004 45334 512604 45418
rect 512004 45098 512186 45334
rect 512422 45098 512604 45334
rect 512004 9654 512604 45098
rect 512004 9418 512186 9654
rect 512422 9418 512604 9654
rect 512004 9334 512604 9418
rect 512004 9098 512186 9334
rect 512422 9098 512604 9334
rect 512004 -4026 512604 9098
rect 512004 -4262 512186 -4026
rect 512422 -4262 512604 -4026
rect 512004 -4346 512604 -4262
rect 512004 -4582 512186 -4346
rect 512422 -4582 512604 -4346
rect 512004 -5524 512604 -4582
rect 515604 697254 516204 709802
rect 533604 711278 534204 711300
rect 533604 711042 533786 711278
rect 534022 711042 534204 711278
rect 533604 710958 534204 711042
rect 533604 710722 533786 710958
rect 534022 710722 534204 710958
rect 530004 709438 530604 709460
rect 530004 709202 530186 709438
rect 530422 709202 530604 709438
rect 530004 709118 530604 709202
rect 530004 708882 530186 709118
rect 530422 708882 530604 709118
rect 526404 707598 527004 707620
rect 526404 707362 526586 707598
rect 526822 707362 527004 707598
rect 526404 707278 527004 707362
rect 526404 707042 526586 707278
rect 526822 707042 527004 707278
rect 515604 697018 515786 697254
rect 516022 697018 516204 697254
rect 515604 696934 516204 697018
rect 515604 696698 515786 696934
rect 516022 696698 516204 696934
rect 515604 661254 516204 696698
rect 515604 661018 515786 661254
rect 516022 661018 516204 661254
rect 515604 660934 516204 661018
rect 515604 660698 515786 660934
rect 516022 660698 516204 660934
rect 515604 625254 516204 660698
rect 515604 625018 515786 625254
rect 516022 625018 516204 625254
rect 515604 624934 516204 625018
rect 515604 624698 515786 624934
rect 516022 624698 516204 624934
rect 515604 589254 516204 624698
rect 515604 589018 515786 589254
rect 516022 589018 516204 589254
rect 515604 588934 516204 589018
rect 515604 588698 515786 588934
rect 516022 588698 516204 588934
rect 515604 553254 516204 588698
rect 515604 553018 515786 553254
rect 516022 553018 516204 553254
rect 515604 552934 516204 553018
rect 515604 552698 515786 552934
rect 516022 552698 516204 552934
rect 515604 517254 516204 552698
rect 515604 517018 515786 517254
rect 516022 517018 516204 517254
rect 515604 516934 516204 517018
rect 515604 516698 515786 516934
rect 516022 516698 516204 516934
rect 515604 481254 516204 516698
rect 515604 481018 515786 481254
rect 516022 481018 516204 481254
rect 515604 480934 516204 481018
rect 515604 480698 515786 480934
rect 516022 480698 516204 480934
rect 515604 445254 516204 480698
rect 515604 445018 515786 445254
rect 516022 445018 516204 445254
rect 515604 444934 516204 445018
rect 515604 444698 515786 444934
rect 516022 444698 516204 444934
rect 515604 409254 516204 444698
rect 515604 409018 515786 409254
rect 516022 409018 516204 409254
rect 515604 408934 516204 409018
rect 515604 408698 515786 408934
rect 516022 408698 516204 408934
rect 515604 373254 516204 408698
rect 515604 373018 515786 373254
rect 516022 373018 516204 373254
rect 515604 372934 516204 373018
rect 515604 372698 515786 372934
rect 516022 372698 516204 372934
rect 515604 337254 516204 372698
rect 515604 337018 515786 337254
rect 516022 337018 516204 337254
rect 515604 336934 516204 337018
rect 515604 336698 515786 336934
rect 516022 336698 516204 336934
rect 515604 301254 516204 336698
rect 515604 301018 515786 301254
rect 516022 301018 516204 301254
rect 515604 300934 516204 301018
rect 515604 300698 515786 300934
rect 516022 300698 516204 300934
rect 515604 265254 516204 300698
rect 515604 265018 515786 265254
rect 516022 265018 516204 265254
rect 515604 264934 516204 265018
rect 515604 264698 515786 264934
rect 516022 264698 516204 264934
rect 515604 229254 516204 264698
rect 515604 229018 515786 229254
rect 516022 229018 516204 229254
rect 515604 228934 516204 229018
rect 515604 228698 515786 228934
rect 516022 228698 516204 228934
rect 515604 193254 516204 228698
rect 515604 193018 515786 193254
rect 516022 193018 516204 193254
rect 515604 192934 516204 193018
rect 515604 192698 515786 192934
rect 516022 192698 516204 192934
rect 515604 157254 516204 192698
rect 515604 157018 515786 157254
rect 516022 157018 516204 157254
rect 515604 156934 516204 157018
rect 515604 156698 515786 156934
rect 516022 156698 516204 156934
rect 515604 121254 516204 156698
rect 515604 121018 515786 121254
rect 516022 121018 516204 121254
rect 515604 120934 516204 121018
rect 515604 120698 515786 120934
rect 516022 120698 516204 120934
rect 515604 85254 516204 120698
rect 515604 85018 515786 85254
rect 516022 85018 516204 85254
rect 515604 84934 516204 85018
rect 515604 84698 515786 84934
rect 516022 84698 516204 84934
rect 515604 49254 516204 84698
rect 515604 49018 515786 49254
rect 516022 49018 516204 49254
rect 515604 48934 516204 49018
rect 515604 48698 515786 48934
rect 516022 48698 516204 48934
rect 515604 13254 516204 48698
rect 515604 13018 515786 13254
rect 516022 13018 516204 13254
rect 515604 12934 516204 13018
rect 515604 12698 515786 12934
rect 516022 12698 516204 12934
rect 497604 -7022 497786 -6786
rect 498022 -7022 498204 -6786
rect 497604 -7106 498204 -7022
rect 497604 -7342 497786 -7106
rect 498022 -7342 498204 -7106
rect 497604 -7364 498204 -7342
rect 515604 -5866 516204 12698
rect 522804 705758 523404 705780
rect 522804 705522 522986 705758
rect 523222 705522 523404 705758
rect 522804 705438 523404 705522
rect 522804 705202 522986 705438
rect 523222 705202 523404 705438
rect 522804 668454 523404 705202
rect 522804 668218 522986 668454
rect 523222 668218 523404 668454
rect 522804 668134 523404 668218
rect 522804 667898 522986 668134
rect 523222 667898 523404 668134
rect 522804 632454 523404 667898
rect 522804 632218 522986 632454
rect 523222 632218 523404 632454
rect 522804 632134 523404 632218
rect 522804 631898 522986 632134
rect 523222 631898 523404 632134
rect 522804 596454 523404 631898
rect 522804 596218 522986 596454
rect 523222 596218 523404 596454
rect 522804 596134 523404 596218
rect 522804 595898 522986 596134
rect 523222 595898 523404 596134
rect 522804 560454 523404 595898
rect 522804 560218 522986 560454
rect 523222 560218 523404 560454
rect 522804 560134 523404 560218
rect 522804 559898 522986 560134
rect 523222 559898 523404 560134
rect 522804 524454 523404 559898
rect 522804 524218 522986 524454
rect 523222 524218 523404 524454
rect 522804 524134 523404 524218
rect 522804 523898 522986 524134
rect 523222 523898 523404 524134
rect 522804 488454 523404 523898
rect 522804 488218 522986 488454
rect 523222 488218 523404 488454
rect 522804 488134 523404 488218
rect 522804 487898 522986 488134
rect 523222 487898 523404 488134
rect 522804 452454 523404 487898
rect 522804 452218 522986 452454
rect 523222 452218 523404 452454
rect 522804 452134 523404 452218
rect 522804 451898 522986 452134
rect 523222 451898 523404 452134
rect 522804 416454 523404 451898
rect 522804 416218 522986 416454
rect 523222 416218 523404 416454
rect 522804 416134 523404 416218
rect 522804 415898 522986 416134
rect 523222 415898 523404 416134
rect 522804 380454 523404 415898
rect 522804 380218 522986 380454
rect 523222 380218 523404 380454
rect 522804 380134 523404 380218
rect 522804 379898 522986 380134
rect 523222 379898 523404 380134
rect 522804 344454 523404 379898
rect 522804 344218 522986 344454
rect 523222 344218 523404 344454
rect 522804 344134 523404 344218
rect 522804 343898 522986 344134
rect 523222 343898 523404 344134
rect 522804 308454 523404 343898
rect 522804 308218 522986 308454
rect 523222 308218 523404 308454
rect 522804 308134 523404 308218
rect 522804 307898 522986 308134
rect 523222 307898 523404 308134
rect 522804 272454 523404 307898
rect 522804 272218 522986 272454
rect 523222 272218 523404 272454
rect 522804 272134 523404 272218
rect 522804 271898 522986 272134
rect 523222 271898 523404 272134
rect 522804 236454 523404 271898
rect 522804 236218 522986 236454
rect 523222 236218 523404 236454
rect 522804 236134 523404 236218
rect 522804 235898 522986 236134
rect 523222 235898 523404 236134
rect 522804 200454 523404 235898
rect 522804 200218 522986 200454
rect 523222 200218 523404 200454
rect 522804 200134 523404 200218
rect 522804 199898 522986 200134
rect 523222 199898 523404 200134
rect 522804 164454 523404 199898
rect 522804 164218 522986 164454
rect 523222 164218 523404 164454
rect 522804 164134 523404 164218
rect 522804 163898 522986 164134
rect 523222 163898 523404 164134
rect 522804 128454 523404 163898
rect 522804 128218 522986 128454
rect 523222 128218 523404 128454
rect 522804 128134 523404 128218
rect 522804 127898 522986 128134
rect 523222 127898 523404 128134
rect 522804 92454 523404 127898
rect 522804 92218 522986 92454
rect 523222 92218 523404 92454
rect 522804 92134 523404 92218
rect 522804 91898 522986 92134
rect 523222 91898 523404 92134
rect 522804 56454 523404 91898
rect 522804 56218 522986 56454
rect 523222 56218 523404 56454
rect 522804 56134 523404 56218
rect 522804 55898 522986 56134
rect 523222 55898 523404 56134
rect 522804 20454 523404 55898
rect 522804 20218 522986 20454
rect 523222 20218 523404 20454
rect 522804 20134 523404 20218
rect 522804 19898 522986 20134
rect 523222 19898 523404 20134
rect 522804 -1266 523404 19898
rect 522804 -1502 522986 -1266
rect 523222 -1502 523404 -1266
rect 522804 -1586 523404 -1502
rect 522804 -1822 522986 -1586
rect 523222 -1822 523404 -1586
rect 522804 -1844 523404 -1822
rect 526404 672054 527004 707042
rect 526404 671818 526586 672054
rect 526822 671818 527004 672054
rect 526404 671734 527004 671818
rect 526404 671498 526586 671734
rect 526822 671498 527004 671734
rect 526404 636054 527004 671498
rect 526404 635818 526586 636054
rect 526822 635818 527004 636054
rect 526404 635734 527004 635818
rect 526404 635498 526586 635734
rect 526822 635498 527004 635734
rect 526404 600054 527004 635498
rect 526404 599818 526586 600054
rect 526822 599818 527004 600054
rect 526404 599734 527004 599818
rect 526404 599498 526586 599734
rect 526822 599498 527004 599734
rect 526404 564054 527004 599498
rect 526404 563818 526586 564054
rect 526822 563818 527004 564054
rect 526404 563734 527004 563818
rect 526404 563498 526586 563734
rect 526822 563498 527004 563734
rect 526404 528054 527004 563498
rect 526404 527818 526586 528054
rect 526822 527818 527004 528054
rect 526404 527734 527004 527818
rect 526404 527498 526586 527734
rect 526822 527498 527004 527734
rect 526404 492054 527004 527498
rect 526404 491818 526586 492054
rect 526822 491818 527004 492054
rect 526404 491734 527004 491818
rect 526404 491498 526586 491734
rect 526822 491498 527004 491734
rect 526404 456054 527004 491498
rect 526404 455818 526586 456054
rect 526822 455818 527004 456054
rect 526404 455734 527004 455818
rect 526404 455498 526586 455734
rect 526822 455498 527004 455734
rect 526404 420054 527004 455498
rect 526404 419818 526586 420054
rect 526822 419818 527004 420054
rect 526404 419734 527004 419818
rect 526404 419498 526586 419734
rect 526822 419498 527004 419734
rect 526404 384054 527004 419498
rect 526404 383818 526586 384054
rect 526822 383818 527004 384054
rect 526404 383734 527004 383818
rect 526404 383498 526586 383734
rect 526822 383498 527004 383734
rect 526404 348054 527004 383498
rect 526404 347818 526586 348054
rect 526822 347818 527004 348054
rect 526404 347734 527004 347818
rect 526404 347498 526586 347734
rect 526822 347498 527004 347734
rect 526404 312054 527004 347498
rect 526404 311818 526586 312054
rect 526822 311818 527004 312054
rect 526404 311734 527004 311818
rect 526404 311498 526586 311734
rect 526822 311498 527004 311734
rect 526404 276054 527004 311498
rect 526404 275818 526586 276054
rect 526822 275818 527004 276054
rect 526404 275734 527004 275818
rect 526404 275498 526586 275734
rect 526822 275498 527004 275734
rect 526404 240054 527004 275498
rect 526404 239818 526586 240054
rect 526822 239818 527004 240054
rect 526404 239734 527004 239818
rect 526404 239498 526586 239734
rect 526822 239498 527004 239734
rect 526404 204054 527004 239498
rect 526404 203818 526586 204054
rect 526822 203818 527004 204054
rect 526404 203734 527004 203818
rect 526404 203498 526586 203734
rect 526822 203498 527004 203734
rect 526404 168054 527004 203498
rect 526404 167818 526586 168054
rect 526822 167818 527004 168054
rect 526404 167734 527004 167818
rect 526404 167498 526586 167734
rect 526822 167498 527004 167734
rect 526404 132054 527004 167498
rect 526404 131818 526586 132054
rect 526822 131818 527004 132054
rect 526404 131734 527004 131818
rect 526404 131498 526586 131734
rect 526822 131498 527004 131734
rect 526404 96054 527004 131498
rect 526404 95818 526586 96054
rect 526822 95818 527004 96054
rect 526404 95734 527004 95818
rect 526404 95498 526586 95734
rect 526822 95498 527004 95734
rect 526404 60054 527004 95498
rect 526404 59818 526586 60054
rect 526822 59818 527004 60054
rect 526404 59734 527004 59818
rect 526404 59498 526586 59734
rect 526822 59498 527004 59734
rect 526404 24054 527004 59498
rect 526404 23818 526586 24054
rect 526822 23818 527004 24054
rect 526404 23734 527004 23818
rect 526404 23498 526586 23734
rect 526822 23498 527004 23734
rect 526404 -3106 527004 23498
rect 526404 -3342 526586 -3106
rect 526822 -3342 527004 -3106
rect 526404 -3426 527004 -3342
rect 526404 -3662 526586 -3426
rect 526822 -3662 527004 -3426
rect 526404 -3684 527004 -3662
rect 530004 675654 530604 708882
rect 530004 675418 530186 675654
rect 530422 675418 530604 675654
rect 530004 675334 530604 675418
rect 530004 675098 530186 675334
rect 530422 675098 530604 675334
rect 530004 639654 530604 675098
rect 530004 639418 530186 639654
rect 530422 639418 530604 639654
rect 530004 639334 530604 639418
rect 530004 639098 530186 639334
rect 530422 639098 530604 639334
rect 530004 603654 530604 639098
rect 530004 603418 530186 603654
rect 530422 603418 530604 603654
rect 530004 603334 530604 603418
rect 530004 603098 530186 603334
rect 530422 603098 530604 603334
rect 530004 567654 530604 603098
rect 530004 567418 530186 567654
rect 530422 567418 530604 567654
rect 530004 567334 530604 567418
rect 530004 567098 530186 567334
rect 530422 567098 530604 567334
rect 530004 531654 530604 567098
rect 530004 531418 530186 531654
rect 530422 531418 530604 531654
rect 530004 531334 530604 531418
rect 530004 531098 530186 531334
rect 530422 531098 530604 531334
rect 530004 495654 530604 531098
rect 530004 495418 530186 495654
rect 530422 495418 530604 495654
rect 530004 495334 530604 495418
rect 530004 495098 530186 495334
rect 530422 495098 530604 495334
rect 530004 459654 530604 495098
rect 530004 459418 530186 459654
rect 530422 459418 530604 459654
rect 530004 459334 530604 459418
rect 530004 459098 530186 459334
rect 530422 459098 530604 459334
rect 530004 423654 530604 459098
rect 530004 423418 530186 423654
rect 530422 423418 530604 423654
rect 530004 423334 530604 423418
rect 530004 423098 530186 423334
rect 530422 423098 530604 423334
rect 530004 387654 530604 423098
rect 530004 387418 530186 387654
rect 530422 387418 530604 387654
rect 530004 387334 530604 387418
rect 530004 387098 530186 387334
rect 530422 387098 530604 387334
rect 530004 351654 530604 387098
rect 530004 351418 530186 351654
rect 530422 351418 530604 351654
rect 530004 351334 530604 351418
rect 530004 351098 530186 351334
rect 530422 351098 530604 351334
rect 530004 315654 530604 351098
rect 530004 315418 530186 315654
rect 530422 315418 530604 315654
rect 530004 315334 530604 315418
rect 530004 315098 530186 315334
rect 530422 315098 530604 315334
rect 530004 279654 530604 315098
rect 530004 279418 530186 279654
rect 530422 279418 530604 279654
rect 530004 279334 530604 279418
rect 530004 279098 530186 279334
rect 530422 279098 530604 279334
rect 530004 243654 530604 279098
rect 530004 243418 530186 243654
rect 530422 243418 530604 243654
rect 530004 243334 530604 243418
rect 530004 243098 530186 243334
rect 530422 243098 530604 243334
rect 530004 207654 530604 243098
rect 530004 207418 530186 207654
rect 530422 207418 530604 207654
rect 530004 207334 530604 207418
rect 530004 207098 530186 207334
rect 530422 207098 530604 207334
rect 530004 171654 530604 207098
rect 530004 171418 530186 171654
rect 530422 171418 530604 171654
rect 530004 171334 530604 171418
rect 530004 171098 530186 171334
rect 530422 171098 530604 171334
rect 530004 135654 530604 171098
rect 530004 135418 530186 135654
rect 530422 135418 530604 135654
rect 530004 135334 530604 135418
rect 530004 135098 530186 135334
rect 530422 135098 530604 135334
rect 530004 99654 530604 135098
rect 530004 99418 530186 99654
rect 530422 99418 530604 99654
rect 530004 99334 530604 99418
rect 530004 99098 530186 99334
rect 530422 99098 530604 99334
rect 530004 63654 530604 99098
rect 530004 63418 530186 63654
rect 530422 63418 530604 63654
rect 530004 63334 530604 63418
rect 530004 63098 530186 63334
rect 530422 63098 530604 63334
rect 530004 27654 530604 63098
rect 530004 27418 530186 27654
rect 530422 27418 530604 27654
rect 530004 27334 530604 27418
rect 530004 27098 530186 27334
rect 530422 27098 530604 27334
rect 530004 -4946 530604 27098
rect 530004 -5182 530186 -4946
rect 530422 -5182 530604 -4946
rect 530004 -5266 530604 -5182
rect 530004 -5502 530186 -5266
rect 530422 -5502 530604 -5266
rect 530004 -5524 530604 -5502
rect 533604 679254 534204 710722
rect 551604 710358 552204 711300
rect 551604 710122 551786 710358
rect 552022 710122 552204 710358
rect 551604 710038 552204 710122
rect 551604 709802 551786 710038
rect 552022 709802 552204 710038
rect 548004 708518 548604 709460
rect 548004 708282 548186 708518
rect 548422 708282 548604 708518
rect 548004 708198 548604 708282
rect 548004 707962 548186 708198
rect 548422 707962 548604 708198
rect 544404 706678 545004 707620
rect 544404 706442 544586 706678
rect 544822 706442 545004 706678
rect 544404 706358 545004 706442
rect 544404 706122 544586 706358
rect 544822 706122 545004 706358
rect 533604 679018 533786 679254
rect 534022 679018 534204 679254
rect 533604 678934 534204 679018
rect 533604 678698 533786 678934
rect 534022 678698 534204 678934
rect 533604 643254 534204 678698
rect 533604 643018 533786 643254
rect 534022 643018 534204 643254
rect 533604 642934 534204 643018
rect 533604 642698 533786 642934
rect 534022 642698 534204 642934
rect 533604 607254 534204 642698
rect 533604 607018 533786 607254
rect 534022 607018 534204 607254
rect 533604 606934 534204 607018
rect 533604 606698 533786 606934
rect 534022 606698 534204 606934
rect 533604 571254 534204 606698
rect 533604 571018 533786 571254
rect 534022 571018 534204 571254
rect 533604 570934 534204 571018
rect 533604 570698 533786 570934
rect 534022 570698 534204 570934
rect 533604 535254 534204 570698
rect 533604 535018 533786 535254
rect 534022 535018 534204 535254
rect 533604 534934 534204 535018
rect 533604 534698 533786 534934
rect 534022 534698 534204 534934
rect 533604 499254 534204 534698
rect 533604 499018 533786 499254
rect 534022 499018 534204 499254
rect 533604 498934 534204 499018
rect 533604 498698 533786 498934
rect 534022 498698 534204 498934
rect 533604 463254 534204 498698
rect 533604 463018 533786 463254
rect 534022 463018 534204 463254
rect 533604 462934 534204 463018
rect 533604 462698 533786 462934
rect 534022 462698 534204 462934
rect 533604 427254 534204 462698
rect 533604 427018 533786 427254
rect 534022 427018 534204 427254
rect 533604 426934 534204 427018
rect 533604 426698 533786 426934
rect 534022 426698 534204 426934
rect 533604 391254 534204 426698
rect 533604 391018 533786 391254
rect 534022 391018 534204 391254
rect 533604 390934 534204 391018
rect 533604 390698 533786 390934
rect 534022 390698 534204 390934
rect 533604 355254 534204 390698
rect 533604 355018 533786 355254
rect 534022 355018 534204 355254
rect 533604 354934 534204 355018
rect 533604 354698 533786 354934
rect 534022 354698 534204 354934
rect 533604 319254 534204 354698
rect 533604 319018 533786 319254
rect 534022 319018 534204 319254
rect 533604 318934 534204 319018
rect 533604 318698 533786 318934
rect 534022 318698 534204 318934
rect 533604 283254 534204 318698
rect 533604 283018 533786 283254
rect 534022 283018 534204 283254
rect 533604 282934 534204 283018
rect 533604 282698 533786 282934
rect 534022 282698 534204 282934
rect 533604 247254 534204 282698
rect 533604 247018 533786 247254
rect 534022 247018 534204 247254
rect 533604 246934 534204 247018
rect 533604 246698 533786 246934
rect 534022 246698 534204 246934
rect 533604 211254 534204 246698
rect 533604 211018 533786 211254
rect 534022 211018 534204 211254
rect 533604 210934 534204 211018
rect 533604 210698 533786 210934
rect 534022 210698 534204 210934
rect 533604 175254 534204 210698
rect 533604 175018 533786 175254
rect 534022 175018 534204 175254
rect 533604 174934 534204 175018
rect 533604 174698 533786 174934
rect 534022 174698 534204 174934
rect 533604 139254 534204 174698
rect 533604 139018 533786 139254
rect 534022 139018 534204 139254
rect 533604 138934 534204 139018
rect 533604 138698 533786 138934
rect 534022 138698 534204 138934
rect 533604 103254 534204 138698
rect 533604 103018 533786 103254
rect 534022 103018 534204 103254
rect 533604 102934 534204 103018
rect 533604 102698 533786 102934
rect 534022 102698 534204 102934
rect 533604 67254 534204 102698
rect 533604 67018 533786 67254
rect 534022 67018 534204 67254
rect 533604 66934 534204 67018
rect 533604 66698 533786 66934
rect 534022 66698 534204 66934
rect 533604 31254 534204 66698
rect 533604 31018 533786 31254
rect 534022 31018 534204 31254
rect 533604 30934 534204 31018
rect 533604 30698 533786 30934
rect 534022 30698 534204 30934
rect 515604 -6102 515786 -5866
rect 516022 -6102 516204 -5866
rect 515604 -6186 516204 -6102
rect 515604 -6422 515786 -6186
rect 516022 -6422 516204 -6186
rect 515604 -7364 516204 -6422
rect 533604 -6786 534204 30698
rect 540804 704838 541404 705780
rect 540804 704602 540986 704838
rect 541222 704602 541404 704838
rect 540804 704518 541404 704602
rect 540804 704282 540986 704518
rect 541222 704282 541404 704518
rect 540804 686454 541404 704282
rect 540804 686218 540986 686454
rect 541222 686218 541404 686454
rect 540804 686134 541404 686218
rect 540804 685898 540986 686134
rect 541222 685898 541404 686134
rect 540804 650454 541404 685898
rect 540804 650218 540986 650454
rect 541222 650218 541404 650454
rect 540804 650134 541404 650218
rect 540804 649898 540986 650134
rect 541222 649898 541404 650134
rect 540804 614454 541404 649898
rect 540804 614218 540986 614454
rect 541222 614218 541404 614454
rect 540804 614134 541404 614218
rect 540804 613898 540986 614134
rect 541222 613898 541404 614134
rect 540804 578454 541404 613898
rect 540804 578218 540986 578454
rect 541222 578218 541404 578454
rect 540804 578134 541404 578218
rect 540804 577898 540986 578134
rect 541222 577898 541404 578134
rect 540804 542454 541404 577898
rect 540804 542218 540986 542454
rect 541222 542218 541404 542454
rect 540804 542134 541404 542218
rect 540804 541898 540986 542134
rect 541222 541898 541404 542134
rect 540804 506454 541404 541898
rect 540804 506218 540986 506454
rect 541222 506218 541404 506454
rect 540804 506134 541404 506218
rect 540804 505898 540986 506134
rect 541222 505898 541404 506134
rect 540804 470454 541404 505898
rect 540804 470218 540986 470454
rect 541222 470218 541404 470454
rect 540804 470134 541404 470218
rect 540804 469898 540986 470134
rect 541222 469898 541404 470134
rect 540804 434454 541404 469898
rect 540804 434218 540986 434454
rect 541222 434218 541404 434454
rect 540804 434134 541404 434218
rect 540804 433898 540986 434134
rect 541222 433898 541404 434134
rect 540804 398454 541404 433898
rect 540804 398218 540986 398454
rect 541222 398218 541404 398454
rect 540804 398134 541404 398218
rect 540804 397898 540986 398134
rect 541222 397898 541404 398134
rect 540804 362454 541404 397898
rect 540804 362218 540986 362454
rect 541222 362218 541404 362454
rect 540804 362134 541404 362218
rect 540804 361898 540986 362134
rect 541222 361898 541404 362134
rect 540804 326454 541404 361898
rect 540804 326218 540986 326454
rect 541222 326218 541404 326454
rect 540804 326134 541404 326218
rect 540804 325898 540986 326134
rect 541222 325898 541404 326134
rect 540804 290454 541404 325898
rect 540804 290218 540986 290454
rect 541222 290218 541404 290454
rect 540804 290134 541404 290218
rect 540804 289898 540986 290134
rect 541222 289898 541404 290134
rect 540804 254454 541404 289898
rect 540804 254218 540986 254454
rect 541222 254218 541404 254454
rect 540804 254134 541404 254218
rect 540804 253898 540986 254134
rect 541222 253898 541404 254134
rect 540804 218454 541404 253898
rect 540804 218218 540986 218454
rect 541222 218218 541404 218454
rect 540804 218134 541404 218218
rect 540804 217898 540986 218134
rect 541222 217898 541404 218134
rect 540804 182454 541404 217898
rect 540804 182218 540986 182454
rect 541222 182218 541404 182454
rect 540804 182134 541404 182218
rect 540804 181898 540986 182134
rect 541222 181898 541404 182134
rect 540804 146454 541404 181898
rect 540804 146218 540986 146454
rect 541222 146218 541404 146454
rect 540804 146134 541404 146218
rect 540804 145898 540986 146134
rect 541222 145898 541404 146134
rect 540804 110454 541404 145898
rect 540804 110218 540986 110454
rect 541222 110218 541404 110454
rect 540804 110134 541404 110218
rect 540804 109898 540986 110134
rect 541222 109898 541404 110134
rect 540804 74454 541404 109898
rect 540804 74218 540986 74454
rect 541222 74218 541404 74454
rect 540804 74134 541404 74218
rect 540804 73898 540986 74134
rect 541222 73898 541404 74134
rect 540804 38454 541404 73898
rect 540804 38218 540986 38454
rect 541222 38218 541404 38454
rect 540804 38134 541404 38218
rect 540804 37898 540986 38134
rect 541222 37898 541404 38134
rect 540804 2454 541404 37898
rect 540804 2218 540986 2454
rect 541222 2218 541404 2454
rect 540804 2134 541404 2218
rect 540804 1898 540986 2134
rect 541222 1898 541404 2134
rect 540804 -346 541404 1898
rect 540804 -582 540986 -346
rect 541222 -582 541404 -346
rect 540804 -666 541404 -582
rect 540804 -902 540986 -666
rect 541222 -902 541404 -666
rect 540804 -1844 541404 -902
rect 544404 690054 545004 706122
rect 544404 689818 544586 690054
rect 544822 689818 545004 690054
rect 544404 689734 545004 689818
rect 544404 689498 544586 689734
rect 544822 689498 545004 689734
rect 544404 654054 545004 689498
rect 544404 653818 544586 654054
rect 544822 653818 545004 654054
rect 544404 653734 545004 653818
rect 544404 653498 544586 653734
rect 544822 653498 545004 653734
rect 544404 618054 545004 653498
rect 544404 617818 544586 618054
rect 544822 617818 545004 618054
rect 544404 617734 545004 617818
rect 544404 617498 544586 617734
rect 544822 617498 545004 617734
rect 544404 582054 545004 617498
rect 544404 581818 544586 582054
rect 544822 581818 545004 582054
rect 544404 581734 545004 581818
rect 544404 581498 544586 581734
rect 544822 581498 545004 581734
rect 544404 546054 545004 581498
rect 544404 545818 544586 546054
rect 544822 545818 545004 546054
rect 544404 545734 545004 545818
rect 544404 545498 544586 545734
rect 544822 545498 545004 545734
rect 544404 510054 545004 545498
rect 544404 509818 544586 510054
rect 544822 509818 545004 510054
rect 544404 509734 545004 509818
rect 544404 509498 544586 509734
rect 544822 509498 545004 509734
rect 544404 474054 545004 509498
rect 544404 473818 544586 474054
rect 544822 473818 545004 474054
rect 544404 473734 545004 473818
rect 544404 473498 544586 473734
rect 544822 473498 545004 473734
rect 544404 438054 545004 473498
rect 544404 437818 544586 438054
rect 544822 437818 545004 438054
rect 544404 437734 545004 437818
rect 544404 437498 544586 437734
rect 544822 437498 545004 437734
rect 544404 402054 545004 437498
rect 544404 401818 544586 402054
rect 544822 401818 545004 402054
rect 544404 401734 545004 401818
rect 544404 401498 544586 401734
rect 544822 401498 545004 401734
rect 544404 366054 545004 401498
rect 544404 365818 544586 366054
rect 544822 365818 545004 366054
rect 544404 365734 545004 365818
rect 544404 365498 544586 365734
rect 544822 365498 545004 365734
rect 544404 330054 545004 365498
rect 544404 329818 544586 330054
rect 544822 329818 545004 330054
rect 544404 329734 545004 329818
rect 544404 329498 544586 329734
rect 544822 329498 545004 329734
rect 544404 294054 545004 329498
rect 544404 293818 544586 294054
rect 544822 293818 545004 294054
rect 544404 293734 545004 293818
rect 544404 293498 544586 293734
rect 544822 293498 545004 293734
rect 544404 258054 545004 293498
rect 544404 257818 544586 258054
rect 544822 257818 545004 258054
rect 544404 257734 545004 257818
rect 544404 257498 544586 257734
rect 544822 257498 545004 257734
rect 544404 222054 545004 257498
rect 544404 221818 544586 222054
rect 544822 221818 545004 222054
rect 544404 221734 545004 221818
rect 544404 221498 544586 221734
rect 544822 221498 545004 221734
rect 544404 186054 545004 221498
rect 544404 185818 544586 186054
rect 544822 185818 545004 186054
rect 544404 185734 545004 185818
rect 544404 185498 544586 185734
rect 544822 185498 545004 185734
rect 544404 150054 545004 185498
rect 544404 149818 544586 150054
rect 544822 149818 545004 150054
rect 544404 149734 545004 149818
rect 544404 149498 544586 149734
rect 544822 149498 545004 149734
rect 544404 114054 545004 149498
rect 544404 113818 544586 114054
rect 544822 113818 545004 114054
rect 544404 113734 545004 113818
rect 544404 113498 544586 113734
rect 544822 113498 545004 113734
rect 544404 78054 545004 113498
rect 544404 77818 544586 78054
rect 544822 77818 545004 78054
rect 544404 77734 545004 77818
rect 544404 77498 544586 77734
rect 544822 77498 545004 77734
rect 544404 42054 545004 77498
rect 544404 41818 544586 42054
rect 544822 41818 545004 42054
rect 544404 41734 545004 41818
rect 544404 41498 544586 41734
rect 544822 41498 545004 41734
rect 544404 6054 545004 41498
rect 544404 5818 544586 6054
rect 544822 5818 545004 6054
rect 544404 5734 545004 5818
rect 544404 5498 544586 5734
rect 544822 5498 545004 5734
rect 544404 -2186 545004 5498
rect 544404 -2422 544586 -2186
rect 544822 -2422 545004 -2186
rect 544404 -2506 545004 -2422
rect 544404 -2742 544586 -2506
rect 544822 -2742 545004 -2506
rect 544404 -3684 545004 -2742
rect 548004 693654 548604 707962
rect 548004 693418 548186 693654
rect 548422 693418 548604 693654
rect 548004 693334 548604 693418
rect 548004 693098 548186 693334
rect 548422 693098 548604 693334
rect 548004 657654 548604 693098
rect 548004 657418 548186 657654
rect 548422 657418 548604 657654
rect 548004 657334 548604 657418
rect 548004 657098 548186 657334
rect 548422 657098 548604 657334
rect 548004 621654 548604 657098
rect 548004 621418 548186 621654
rect 548422 621418 548604 621654
rect 548004 621334 548604 621418
rect 548004 621098 548186 621334
rect 548422 621098 548604 621334
rect 548004 585654 548604 621098
rect 548004 585418 548186 585654
rect 548422 585418 548604 585654
rect 548004 585334 548604 585418
rect 548004 585098 548186 585334
rect 548422 585098 548604 585334
rect 548004 549654 548604 585098
rect 548004 549418 548186 549654
rect 548422 549418 548604 549654
rect 548004 549334 548604 549418
rect 548004 549098 548186 549334
rect 548422 549098 548604 549334
rect 548004 513654 548604 549098
rect 548004 513418 548186 513654
rect 548422 513418 548604 513654
rect 548004 513334 548604 513418
rect 548004 513098 548186 513334
rect 548422 513098 548604 513334
rect 548004 477654 548604 513098
rect 548004 477418 548186 477654
rect 548422 477418 548604 477654
rect 548004 477334 548604 477418
rect 548004 477098 548186 477334
rect 548422 477098 548604 477334
rect 548004 441654 548604 477098
rect 548004 441418 548186 441654
rect 548422 441418 548604 441654
rect 548004 441334 548604 441418
rect 548004 441098 548186 441334
rect 548422 441098 548604 441334
rect 548004 405654 548604 441098
rect 548004 405418 548186 405654
rect 548422 405418 548604 405654
rect 548004 405334 548604 405418
rect 548004 405098 548186 405334
rect 548422 405098 548604 405334
rect 548004 369654 548604 405098
rect 548004 369418 548186 369654
rect 548422 369418 548604 369654
rect 548004 369334 548604 369418
rect 548004 369098 548186 369334
rect 548422 369098 548604 369334
rect 548004 333654 548604 369098
rect 548004 333418 548186 333654
rect 548422 333418 548604 333654
rect 548004 333334 548604 333418
rect 548004 333098 548186 333334
rect 548422 333098 548604 333334
rect 548004 297654 548604 333098
rect 548004 297418 548186 297654
rect 548422 297418 548604 297654
rect 548004 297334 548604 297418
rect 548004 297098 548186 297334
rect 548422 297098 548604 297334
rect 548004 261654 548604 297098
rect 548004 261418 548186 261654
rect 548422 261418 548604 261654
rect 548004 261334 548604 261418
rect 548004 261098 548186 261334
rect 548422 261098 548604 261334
rect 548004 225654 548604 261098
rect 548004 225418 548186 225654
rect 548422 225418 548604 225654
rect 548004 225334 548604 225418
rect 548004 225098 548186 225334
rect 548422 225098 548604 225334
rect 548004 189654 548604 225098
rect 548004 189418 548186 189654
rect 548422 189418 548604 189654
rect 548004 189334 548604 189418
rect 548004 189098 548186 189334
rect 548422 189098 548604 189334
rect 548004 153654 548604 189098
rect 548004 153418 548186 153654
rect 548422 153418 548604 153654
rect 548004 153334 548604 153418
rect 548004 153098 548186 153334
rect 548422 153098 548604 153334
rect 548004 117654 548604 153098
rect 548004 117418 548186 117654
rect 548422 117418 548604 117654
rect 548004 117334 548604 117418
rect 548004 117098 548186 117334
rect 548422 117098 548604 117334
rect 548004 81654 548604 117098
rect 548004 81418 548186 81654
rect 548422 81418 548604 81654
rect 548004 81334 548604 81418
rect 548004 81098 548186 81334
rect 548422 81098 548604 81334
rect 548004 45654 548604 81098
rect 548004 45418 548186 45654
rect 548422 45418 548604 45654
rect 548004 45334 548604 45418
rect 548004 45098 548186 45334
rect 548422 45098 548604 45334
rect 548004 9654 548604 45098
rect 548004 9418 548186 9654
rect 548422 9418 548604 9654
rect 548004 9334 548604 9418
rect 548004 9098 548186 9334
rect 548422 9098 548604 9334
rect 548004 -4026 548604 9098
rect 548004 -4262 548186 -4026
rect 548422 -4262 548604 -4026
rect 548004 -4346 548604 -4262
rect 548004 -4582 548186 -4346
rect 548422 -4582 548604 -4346
rect 548004 -5524 548604 -4582
rect 551604 697254 552204 709802
rect 569604 711278 570204 711300
rect 569604 711042 569786 711278
rect 570022 711042 570204 711278
rect 569604 710958 570204 711042
rect 569604 710722 569786 710958
rect 570022 710722 570204 710958
rect 566004 709438 566604 709460
rect 566004 709202 566186 709438
rect 566422 709202 566604 709438
rect 566004 709118 566604 709202
rect 566004 708882 566186 709118
rect 566422 708882 566604 709118
rect 562404 707598 563004 707620
rect 562404 707362 562586 707598
rect 562822 707362 563004 707598
rect 562404 707278 563004 707362
rect 562404 707042 562586 707278
rect 562822 707042 563004 707278
rect 551604 697018 551786 697254
rect 552022 697018 552204 697254
rect 551604 696934 552204 697018
rect 551604 696698 551786 696934
rect 552022 696698 552204 696934
rect 551604 661254 552204 696698
rect 551604 661018 551786 661254
rect 552022 661018 552204 661254
rect 551604 660934 552204 661018
rect 551604 660698 551786 660934
rect 552022 660698 552204 660934
rect 551604 625254 552204 660698
rect 551604 625018 551786 625254
rect 552022 625018 552204 625254
rect 551604 624934 552204 625018
rect 551604 624698 551786 624934
rect 552022 624698 552204 624934
rect 551604 589254 552204 624698
rect 551604 589018 551786 589254
rect 552022 589018 552204 589254
rect 551604 588934 552204 589018
rect 551604 588698 551786 588934
rect 552022 588698 552204 588934
rect 551604 553254 552204 588698
rect 551604 553018 551786 553254
rect 552022 553018 552204 553254
rect 551604 552934 552204 553018
rect 551604 552698 551786 552934
rect 552022 552698 552204 552934
rect 551604 517254 552204 552698
rect 551604 517018 551786 517254
rect 552022 517018 552204 517254
rect 551604 516934 552204 517018
rect 551604 516698 551786 516934
rect 552022 516698 552204 516934
rect 551604 481254 552204 516698
rect 551604 481018 551786 481254
rect 552022 481018 552204 481254
rect 551604 480934 552204 481018
rect 551604 480698 551786 480934
rect 552022 480698 552204 480934
rect 551604 445254 552204 480698
rect 551604 445018 551786 445254
rect 552022 445018 552204 445254
rect 551604 444934 552204 445018
rect 551604 444698 551786 444934
rect 552022 444698 552204 444934
rect 551604 409254 552204 444698
rect 551604 409018 551786 409254
rect 552022 409018 552204 409254
rect 551604 408934 552204 409018
rect 551604 408698 551786 408934
rect 552022 408698 552204 408934
rect 551604 373254 552204 408698
rect 551604 373018 551786 373254
rect 552022 373018 552204 373254
rect 551604 372934 552204 373018
rect 551604 372698 551786 372934
rect 552022 372698 552204 372934
rect 551604 337254 552204 372698
rect 551604 337018 551786 337254
rect 552022 337018 552204 337254
rect 551604 336934 552204 337018
rect 551604 336698 551786 336934
rect 552022 336698 552204 336934
rect 551604 301254 552204 336698
rect 551604 301018 551786 301254
rect 552022 301018 552204 301254
rect 551604 300934 552204 301018
rect 551604 300698 551786 300934
rect 552022 300698 552204 300934
rect 551604 265254 552204 300698
rect 551604 265018 551786 265254
rect 552022 265018 552204 265254
rect 551604 264934 552204 265018
rect 551604 264698 551786 264934
rect 552022 264698 552204 264934
rect 551604 229254 552204 264698
rect 551604 229018 551786 229254
rect 552022 229018 552204 229254
rect 551604 228934 552204 229018
rect 551604 228698 551786 228934
rect 552022 228698 552204 228934
rect 551604 193254 552204 228698
rect 551604 193018 551786 193254
rect 552022 193018 552204 193254
rect 551604 192934 552204 193018
rect 551604 192698 551786 192934
rect 552022 192698 552204 192934
rect 551604 157254 552204 192698
rect 551604 157018 551786 157254
rect 552022 157018 552204 157254
rect 551604 156934 552204 157018
rect 551604 156698 551786 156934
rect 552022 156698 552204 156934
rect 551604 121254 552204 156698
rect 551604 121018 551786 121254
rect 552022 121018 552204 121254
rect 551604 120934 552204 121018
rect 551604 120698 551786 120934
rect 552022 120698 552204 120934
rect 551604 85254 552204 120698
rect 551604 85018 551786 85254
rect 552022 85018 552204 85254
rect 551604 84934 552204 85018
rect 551604 84698 551786 84934
rect 552022 84698 552204 84934
rect 551604 49254 552204 84698
rect 551604 49018 551786 49254
rect 552022 49018 552204 49254
rect 551604 48934 552204 49018
rect 551604 48698 551786 48934
rect 552022 48698 552204 48934
rect 551604 13254 552204 48698
rect 551604 13018 551786 13254
rect 552022 13018 552204 13254
rect 551604 12934 552204 13018
rect 551604 12698 551786 12934
rect 552022 12698 552204 12934
rect 533604 -7022 533786 -6786
rect 534022 -7022 534204 -6786
rect 533604 -7106 534204 -7022
rect 533604 -7342 533786 -7106
rect 534022 -7342 534204 -7106
rect 533604 -7364 534204 -7342
rect 551604 -5866 552204 12698
rect 558804 705758 559404 705780
rect 558804 705522 558986 705758
rect 559222 705522 559404 705758
rect 558804 705438 559404 705522
rect 558804 705202 558986 705438
rect 559222 705202 559404 705438
rect 558804 668454 559404 705202
rect 558804 668218 558986 668454
rect 559222 668218 559404 668454
rect 558804 668134 559404 668218
rect 558804 667898 558986 668134
rect 559222 667898 559404 668134
rect 558804 632454 559404 667898
rect 558804 632218 558986 632454
rect 559222 632218 559404 632454
rect 558804 632134 559404 632218
rect 558804 631898 558986 632134
rect 559222 631898 559404 632134
rect 558804 596454 559404 631898
rect 558804 596218 558986 596454
rect 559222 596218 559404 596454
rect 558804 596134 559404 596218
rect 558804 595898 558986 596134
rect 559222 595898 559404 596134
rect 558804 560454 559404 595898
rect 558804 560218 558986 560454
rect 559222 560218 559404 560454
rect 558804 560134 559404 560218
rect 558804 559898 558986 560134
rect 559222 559898 559404 560134
rect 558804 524454 559404 559898
rect 558804 524218 558986 524454
rect 559222 524218 559404 524454
rect 558804 524134 559404 524218
rect 558804 523898 558986 524134
rect 559222 523898 559404 524134
rect 558804 488454 559404 523898
rect 558804 488218 558986 488454
rect 559222 488218 559404 488454
rect 558804 488134 559404 488218
rect 558804 487898 558986 488134
rect 559222 487898 559404 488134
rect 558804 452454 559404 487898
rect 558804 452218 558986 452454
rect 559222 452218 559404 452454
rect 558804 452134 559404 452218
rect 558804 451898 558986 452134
rect 559222 451898 559404 452134
rect 558804 416454 559404 451898
rect 558804 416218 558986 416454
rect 559222 416218 559404 416454
rect 558804 416134 559404 416218
rect 558804 415898 558986 416134
rect 559222 415898 559404 416134
rect 558804 380454 559404 415898
rect 558804 380218 558986 380454
rect 559222 380218 559404 380454
rect 558804 380134 559404 380218
rect 558804 379898 558986 380134
rect 559222 379898 559404 380134
rect 558804 344454 559404 379898
rect 558804 344218 558986 344454
rect 559222 344218 559404 344454
rect 558804 344134 559404 344218
rect 558804 343898 558986 344134
rect 559222 343898 559404 344134
rect 558804 308454 559404 343898
rect 558804 308218 558986 308454
rect 559222 308218 559404 308454
rect 558804 308134 559404 308218
rect 558804 307898 558986 308134
rect 559222 307898 559404 308134
rect 558804 272454 559404 307898
rect 558804 272218 558986 272454
rect 559222 272218 559404 272454
rect 558804 272134 559404 272218
rect 558804 271898 558986 272134
rect 559222 271898 559404 272134
rect 558804 236454 559404 271898
rect 558804 236218 558986 236454
rect 559222 236218 559404 236454
rect 558804 236134 559404 236218
rect 558804 235898 558986 236134
rect 559222 235898 559404 236134
rect 558804 200454 559404 235898
rect 558804 200218 558986 200454
rect 559222 200218 559404 200454
rect 558804 200134 559404 200218
rect 558804 199898 558986 200134
rect 559222 199898 559404 200134
rect 558804 164454 559404 199898
rect 558804 164218 558986 164454
rect 559222 164218 559404 164454
rect 558804 164134 559404 164218
rect 558804 163898 558986 164134
rect 559222 163898 559404 164134
rect 558804 128454 559404 163898
rect 558804 128218 558986 128454
rect 559222 128218 559404 128454
rect 558804 128134 559404 128218
rect 558804 127898 558986 128134
rect 559222 127898 559404 128134
rect 558804 92454 559404 127898
rect 558804 92218 558986 92454
rect 559222 92218 559404 92454
rect 558804 92134 559404 92218
rect 558804 91898 558986 92134
rect 559222 91898 559404 92134
rect 558804 56454 559404 91898
rect 558804 56218 558986 56454
rect 559222 56218 559404 56454
rect 558804 56134 559404 56218
rect 558804 55898 558986 56134
rect 559222 55898 559404 56134
rect 558804 20454 559404 55898
rect 558804 20218 558986 20454
rect 559222 20218 559404 20454
rect 558804 20134 559404 20218
rect 558804 19898 558986 20134
rect 559222 19898 559404 20134
rect 558804 -1266 559404 19898
rect 558804 -1502 558986 -1266
rect 559222 -1502 559404 -1266
rect 558804 -1586 559404 -1502
rect 558804 -1822 558986 -1586
rect 559222 -1822 559404 -1586
rect 558804 -1844 559404 -1822
rect 562404 672054 563004 707042
rect 562404 671818 562586 672054
rect 562822 671818 563004 672054
rect 562404 671734 563004 671818
rect 562404 671498 562586 671734
rect 562822 671498 563004 671734
rect 562404 636054 563004 671498
rect 562404 635818 562586 636054
rect 562822 635818 563004 636054
rect 562404 635734 563004 635818
rect 562404 635498 562586 635734
rect 562822 635498 563004 635734
rect 562404 600054 563004 635498
rect 562404 599818 562586 600054
rect 562822 599818 563004 600054
rect 562404 599734 563004 599818
rect 562404 599498 562586 599734
rect 562822 599498 563004 599734
rect 562404 564054 563004 599498
rect 562404 563818 562586 564054
rect 562822 563818 563004 564054
rect 562404 563734 563004 563818
rect 562404 563498 562586 563734
rect 562822 563498 563004 563734
rect 562404 528054 563004 563498
rect 562404 527818 562586 528054
rect 562822 527818 563004 528054
rect 562404 527734 563004 527818
rect 562404 527498 562586 527734
rect 562822 527498 563004 527734
rect 562404 492054 563004 527498
rect 562404 491818 562586 492054
rect 562822 491818 563004 492054
rect 562404 491734 563004 491818
rect 562404 491498 562586 491734
rect 562822 491498 563004 491734
rect 562404 456054 563004 491498
rect 562404 455818 562586 456054
rect 562822 455818 563004 456054
rect 562404 455734 563004 455818
rect 562404 455498 562586 455734
rect 562822 455498 563004 455734
rect 562404 420054 563004 455498
rect 562404 419818 562586 420054
rect 562822 419818 563004 420054
rect 562404 419734 563004 419818
rect 562404 419498 562586 419734
rect 562822 419498 563004 419734
rect 562404 384054 563004 419498
rect 562404 383818 562586 384054
rect 562822 383818 563004 384054
rect 562404 383734 563004 383818
rect 562404 383498 562586 383734
rect 562822 383498 563004 383734
rect 562404 348054 563004 383498
rect 562404 347818 562586 348054
rect 562822 347818 563004 348054
rect 562404 347734 563004 347818
rect 562404 347498 562586 347734
rect 562822 347498 563004 347734
rect 562404 312054 563004 347498
rect 562404 311818 562586 312054
rect 562822 311818 563004 312054
rect 562404 311734 563004 311818
rect 562404 311498 562586 311734
rect 562822 311498 563004 311734
rect 562404 276054 563004 311498
rect 562404 275818 562586 276054
rect 562822 275818 563004 276054
rect 562404 275734 563004 275818
rect 562404 275498 562586 275734
rect 562822 275498 563004 275734
rect 562404 240054 563004 275498
rect 562404 239818 562586 240054
rect 562822 239818 563004 240054
rect 562404 239734 563004 239818
rect 562404 239498 562586 239734
rect 562822 239498 563004 239734
rect 562404 204054 563004 239498
rect 562404 203818 562586 204054
rect 562822 203818 563004 204054
rect 562404 203734 563004 203818
rect 562404 203498 562586 203734
rect 562822 203498 563004 203734
rect 562404 168054 563004 203498
rect 562404 167818 562586 168054
rect 562822 167818 563004 168054
rect 562404 167734 563004 167818
rect 562404 167498 562586 167734
rect 562822 167498 563004 167734
rect 562404 132054 563004 167498
rect 562404 131818 562586 132054
rect 562822 131818 563004 132054
rect 562404 131734 563004 131818
rect 562404 131498 562586 131734
rect 562822 131498 563004 131734
rect 562404 96054 563004 131498
rect 562404 95818 562586 96054
rect 562822 95818 563004 96054
rect 562404 95734 563004 95818
rect 562404 95498 562586 95734
rect 562822 95498 563004 95734
rect 562404 60054 563004 95498
rect 562404 59818 562586 60054
rect 562822 59818 563004 60054
rect 562404 59734 563004 59818
rect 562404 59498 562586 59734
rect 562822 59498 563004 59734
rect 562404 24054 563004 59498
rect 562404 23818 562586 24054
rect 562822 23818 563004 24054
rect 562404 23734 563004 23818
rect 562404 23498 562586 23734
rect 562822 23498 563004 23734
rect 562404 -3106 563004 23498
rect 562404 -3342 562586 -3106
rect 562822 -3342 563004 -3106
rect 562404 -3426 563004 -3342
rect 562404 -3662 562586 -3426
rect 562822 -3662 563004 -3426
rect 562404 -3684 563004 -3662
rect 566004 675654 566604 708882
rect 566004 675418 566186 675654
rect 566422 675418 566604 675654
rect 566004 675334 566604 675418
rect 566004 675098 566186 675334
rect 566422 675098 566604 675334
rect 566004 639654 566604 675098
rect 566004 639418 566186 639654
rect 566422 639418 566604 639654
rect 566004 639334 566604 639418
rect 566004 639098 566186 639334
rect 566422 639098 566604 639334
rect 566004 603654 566604 639098
rect 566004 603418 566186 603654
rect 566422 603418 566604 603654
rect 566004 603334 566604 603418
rect 566004 603098 566186 603334
rect 566422 603098 566604 603334
rect 566004 567654 566604 603098
rect 566004 567418 566186 567654
rect 566422 567418 566604 567654
rect 566004 567334 566604 567418
rect 566004 567098 566186 567334
rect 566422 567098 566604 567334
rect 566004 531654 566604 567098
rect 566004 531418 566186 531654
rect 566422 531418 566604 531654
rect 566004 531334 566604 531418
rect 566004 531098 566186 531334
rect 566422 531098 566604 531334
rect 566004 495654 566604 531098
rect 566004 495418 566186 495654
rect 566422 495418 566604 495654
rect 566004 495334 566604 495418
rect 566004 495098 566186 495334
rect 566422 495098 566604 495334
rect 566004 459654 566604 495098
rect 566004 459418 566186 459654
rect 566422 459418 566604 459654
rect 566004 459334 566604 459418
rect 566004 459098 566186 459334
rect 566422 459098 566604 459334
rect 566004 423654 566604 459098
rect 566004 423418 566186 423654
rect 566422 423418 566604 423654
rect 566004 423334 566604 423418
rect 566004 423098 566186 423334
rect 566422 423098 566604 423334
rect 566004 387654 566604 423098
rect 566004 387418 566186 387654
rect 566422 387418 566604 387654
rect 566004 387334 566604 387418
rect 566004 387098 566186 387334
rect 566422 387098 566604 387334
rect 566004 351654 566604 387098
rect 566004 351418 566186 351654
rect 566422 351418 566604 351654
rect 566004 351334 566604 351418
rect 566004 351098 566186 351334
rect 566422 351098 566604 351334
rect 566004 315654 566604 351098
rect 566004 315418 566186 315654
rect 566422 315418 566604 315654
rect 566004 315334 566604 315418
rect 566004 315098 566186 315334
rect 566422 315098 566604 315334
rect 566004 279654 566604 315098
rect 566004 279418 566186 279654
rect 566422 279418 566604 279654
rect 566004 279334 566604 279418
rect 566004 279098 566186 279334
rect 566422 279098 566604 279334
rect 566004 243654 566604 279098
rect 566004 243418 566186 243654
rect 566422 243418 566604 243654
rect 566004 243334 566604 243418
rect 566004 243098 566186 243334
rect 566422 243098 566604 243334
rect 566004 207654 566604 243098
rect 566004 207418 566186 207654
rect 566422 207418 566604 207654
rect 566004 207334 566604 207418
rect 566004 207098 566186 207334
rect 566422 207098 566604 207334
rect 566004 171654 566604 207098
rect 566004 171418 566186 171654
rect 566422 171418 566604 171654
rect 566004 171334 566604 171418
rect 566004 171098 566186 171334
rect 566422 171098 566604 171334
rect 566004 135654 566604 171098
rect 566004 135418 566186 135654
rect 566422 135418 566604 135654
rect 566004 135334 566604 135418
rect 566004 135098 566186 135334
rect 566422 135098 566604 135334
rect 566004 99654 566604 135098
rect 566004 99418 566186 99654
rect 566422 99418 566604 99654
rect 566004 99334 566604 99418
rect 566004 99098 566186 99334
rect 566422 99098 566604 99334
rect 566004 63654 566604 99098
rect 566004 63418 566186 63654
rect 566422 63418 566604 63654
rect 566004 63334 566604 63418
rect 566004 63098 566186 63334
rect 566422 63098 566604 63334
rect 566004 27654 566604 63098
rect 566004 27418 566186 27654
rect 566422 27418 566604 27654
rect 566004 27334 566604 27418
rect 566004 27098 566186 27334
rect 566422 27098 566604 27334
rect 566004 -4946 566604 27098
rect 566004 -5182 566186 -4946
rect 566422 -5182 566604 -4946
rect 566004 -5266 566604 -5182
rect 566004 -5502 566186 -5266
rect 566422 -5502 566604 -5266
rect 566004 -5524 566604 -5502
rect 569604 679254 570204 710722
rect 591760 711278 592360 711300
rect 591760 711042 591942 711278
rect 592178 711042 592360 711278
rect 591760 710958 592360 711042
rect 591760 710722 591942 710958
rect 592178 710722 592360 710958
rect 590840 710358 591440 710380
rect 590840 710122 591022 710358
rect 591258 710122 591440 710358
rect 590840 710038 591440 710122
rect 590840 709802 591022 710038
rect 591258 709802 591440 710038
rect 589920 709438 590520 709460
rect 589920 709202 590102 709438
rect 590338 709202 590520 709438
rect 589920 709118 590520 709202
rect 589920 708882 590102 709118
rect 590338 708882 590520 709118
rect 589000 708518 589600 708540
rect 589000 708282 589182 708518
rect 589418 708282 589600 708518
rect 589000 708198 589600 708282
rect 589000 707962 589182 708198
rect 589418 707962 589600 708198
rect 580404 706678 581004 707620
rect 588080 707598 588680 707620
rect 588080 707362 588262 707598
rect 588498 707362 588680 707598
rect 588080 707278 588680 707362
rect 588080 707042 588262 707278
rect 588498 707042 588680 707278
rect 580404 706442 580586 706678
rect 580822 706442 581004 706678
rect 580404 706358 581004 706442
rect 580404 706122 580586 706358
rect 580822 706122 581004 706358
rect 569604 679018 569786 679254
rect 570022 679018 570204 679254
rect 569604 678934 570204 679018
rect 569604 678698 569786 678934
rect 570022 678698 570204 678934
rect 569604 643254 570204 678698
rect 569604 643018 569786 643254
rect 570022 643018 570204 643254
rect 569604 642934 570204 643018
rect 569604 642698 569786 642934
rect 570022 642698 570204 642934
rect 569604 607254 570204 642698
rect 569604 607018 569786 607254
rect 570022 607018 570204 607254
rect 569604 606934 570204 607018
rect 569604 606698 569786 606934
rect 570022 606698 570204 606934
rect 569604 571254 570204 606698
rect 569604 571018 569786 571254
rect 570022 571018 570204 571254
rect 569604 570934 570204 571018
rect 569604 570698 569786 570934
rect 570022 570698 570204 570934
rect 569604 535254 570204 570698
rect 569604 535018 569786 535254
rect 570022 535018 570204 535254
rect 569604 534934 570204 535018
rect 569604 534698 569786 534934
rect 570022 534698 570204 534934
rect 569604 499254 570204 534698
rect 569604 499018 569786 499254
rect 570022 499018 570204 499254
rect 569604 498934 570204 499018
rect 569604 498698 569786 498934
rect 570022 498698 570204 498934
rect 569604 463254 570204 498698
rect 569604 463018 569786 463254
rect 570022 463018 570204 463254
rect 569604 462934 570204 463018
rect 569604 462698 569786 462934
rect 570022 462698 570204 462934
rect 569604 427254 570204 462698
rect 569604 427018 569786 427254
rect 570022 427018 570204 427254
rect 569604 426934 570204 427018
rect 569604 426698 569786 426934
rect 570022 426698 570204 426934
rect 569604 391254 570204 426698
rect 569604 391018 569786 391254
rect 570022 391018 570204 391254
rect 569604 390934 570204 391018
rect 569604 390698 569786 390934
rect 570022 390698 570204 390934
rect 569604 355254 570204 390698
rect 569604 355018 569786 355254
rect 570022 355018 570204 355254
rect 569604 354934 570204 355018
rect 569604 354698 569786 354934
rect 570022 354698 570204 354934
rect 569604 319254 570204 354698
rect 569604 319018 569786 319254
rect 570022 319018 570204 319254
rect 569604 318934 570204 319018
rect 569604 318698 569786 318934
rect 570022 318698 570204 318934
rect 569604 283254 570204 318698
rect 569604 283018 569786 283254
rect 570022 283018 570204 283254
rect 569604 282934 570204 283018
rect 569604 282698 569786 282934
rect 570022 282698 570204 282934
rect 569604 247254 570204 282698
rect 569604 247018 569786 247254
rect 570022 247018 570204 247254
rect 569604 246934 570204 247018
rect 569604 246698 569786 246934
rect 570022 246698 570204 246934
rect 569604 211254 570204 246698
rect 569604 211018 569786 211254
rect 570022 211018 570204 211254
rect 569604 210934 570204 211018
rect 569604 210698 569786 210934
rect 570022 210698 570204 210934
rect 569604 175254 570204 210698
rect 569604 175018 569786 175254
rect 570022 175018 570204 175254
rect 569604 174934 570204 175018
rect 569604 174698 569786 174934
rect 570022 174698 570204 174934
rect 569604 139254 570204 174698
rect 569604 139018 569786 139254
rect 570022 139018 570204 139254
rect 569604 138934 570204 139018
rect 569604 138698 569786 138934
rect 570022 138698 570204 138934
rect 569604 103254 570204 138698
rect 569604 103018 569786 103254
rect 570022 103018 570204 103254
rect 569604 102934 570204 103018
rect 569604 102698 569786 102934
rect 570022 102698 570204 102934
rect 569604 67254 570204 102698
rect 569604 67018 569786 67254
rect 570022 67018 570204 67254
rect 569604 66934 570204 67018
rect 569604 66698 569786 66934
rect 570022 66698 570204 66934
rect 569604 31254 570204 66698
rect 569604 31018 569786 31254
rect 570022 31018 570204 31254
rect 569604 30934 570204 31018
rect 569604 30698 569786 30934
rect 570022 30698 570204 30934
rect 551604 -6102 551786 -5866
rect 552022 -6102 552204 -5866
rect 551604 -6186 552204 -6102
rect 551604 -6422 551786 -6186
rect 552022 -6422 552204 -6186
rect 551604 -7364 552204 -6422
rect 569604 -6786 570204 30698
rect 576804 704838 577404 705780
rect 576804 704602 576986 704838
rect 577222 704602 577404 704838
rect 576804 704518 577404 704602
rect 576804 704282 576986 704518
rect 577222 704282 577404 704518
rect 576804 686454 577404 704282
rect 576804 686218 576986 686454
rect 577222 686218 577404 686454
rect 576804 686134 577404 686218
rect 576804 685898 576986 686134
rect 577222 685898 577404 686134
rect 576804 650454 577404 685898
rect 576804 650218 576986 650454
rect 577222 650218 577404 650454
rect 576804 650134 577404 650218
rect 576804 649898 576986 650134
rect 577222 649898 577404 650134
rect 576804 614454 577404 649898
rect 576804 614218 576986 614454
rect 577222 614218 577404 614454
rect 576804 614134 577404 614218
rect 576804 613898 576986 614134
rect 577222 613898 577404 614134
rect 576804 578454 577404 613898
rect 576804 578218 576986 578454
rect 577222 578218 577404 578454
rect 576804 578134 577404 578218
rect 576804 577898 576986 578134
rect 577222 577898 577404 578134
rect 576804 542454 577404 577898
rect 576804 542218 576986 542454
rect 577222 542218 577404 542454
rect 576804 542134 577404 542218
rect 576804 541898 576986 542134
rect 577222 541898 577404 542134
rect 576804 506454 577404 541898
rect 576804 506218 576986 506454
rect 577222 506218 577404 506454
rect 576804 506134 577404 506218
rect 576804 505898 576986 506134
rect 577222 505898 577404 506134
rect 576804 470454 577404 505898
rect 576804 470218 576986 470454
rect 577222 470218 577404 470454
rect 576804 470134 577404 470218
rect 576804 469898 576986 470134
rect 577222 469898 577404 470134
rect 576804 434454 577404 469898
rect 576804 434218 576986 434454
rect 577222 434218 577404 434454
rect 576804 434134 577404 434218
rect 576804 433898 576986 434134
rect 577222 433898 577404 434134
rect 576804 398454 577404 433898
rect 576804 398218 576986 398454
rect 577222 398218 577404 398454
rect 576804 398134 577404 398218
rect 576804 397898 576986 398134
rect 577222 397898 577404 398134
rect 576804 362454 577404 397898
rect 576804 362218 576986 362454
rect 577222 362218 577404 362454
rect 576804 362134 577404 362218
rect 576804 361898 576986 362134
rect 577222 361898 577404 362134
rect 576804 326454 577404 361898
rect 576804 326218 576986 326454
rect 577222 326218 577404 326454
rect 576804 326134 577404 326218
rect 576804 325898 576986 326134
rect 577222 325898 577404 326134
rect 576804 290454 577404 325898
rect 576804 290218 576986 290454
rect 577222 290218 577404 290454
rect 576804 290134 577404 290218
rect 576804 289898 576986 290134
rect 577222 289898 577404 290134
rect 576804 254454 577404 289898
rect 576804 254218 576986 254454
rect 577222 254218 577404 254454
rect 576804 254134 577404 254218
rect 576804 253898 576986 254134
rect 577222 253898 577404 254134
rect 576804 218454 577404 253898
rect 576804 218218 576986 218454
rect 577222 218218 577404 218454
rect 576804 218134 577404 218218
rect 576804 217898 576986 218134
rect 577222 217898 577404 218134
rect 576804 182454 577404 217898
rect 576804 182218 576986 182454
rect 577222 182218 577404 182454
rect 576804 182134 577404 182218
rect 576804 181898 576986 182134
rect 577222 181898 577404 182134
rect 576804 146454 577404 181898
rect 576804 146218 576986 146454
rect 577222 146218 577404 146454
rect 576804 146134 577404 146218
rect 576804 145898 576986 146134
rect 577222 145898 577404 146134
rect 576804 110454 577404 145898
rect 576804 110218 576986 110454
rect 577222 110218 577404 110454
rect 576804 110134 577404 110218
rect 576804 109898 576986 110134
rect 577222 109898 577404 110134
rect 576804 74454 577404 109898
rect 576804 74218 576986 74454
rect 577222 74218 577404 74454
rect 576804 74134 577404 74218
rect 576804 73898 576986 74134
rect 577222 73898 577404 74134
rect 576804 38454 577404 73898
rect 576804 38218 576986 38454
rect 577222 38218 577404 38454
rect 576804 38134 577404 38218
rect 576804 37898 576986 38134
rect 577222 37898 577404 38134
rect 576804 2454 577404 37898
rect 576804 2218 576986 2454
rect 577222 2218 577404 2454
rect 576804 2134 577404 2218
rect 576804 1898 576986 2134
rect 577222 1898 577404 2134
rect 576804 -346 577404 1898
rect 576804 -582 576986 -346
rect 577222 -582 577404 -346
rect 576804 -666 577404 -582
rect 576804 -902 576986 -666
rect 577222 -902 577404 -666
rect 576804 -1844 577404 -902
rect 580404 690054 581004 706122
rect 587160 706678 587760 706700
rect 587160 706442 587342 706678
rect 587578 706442 587760 706678
rect 587160 706358 587760 706442
rect 587160 706122 587342 706358
rect 587578 706122 587760 706358
rect 586240 705758 586840 705780
rect 586240 705522 586422 705758
rect 586658 705522 586840 705758
rect 586240 705438 586840 705522
rect 586240 705202 586422 705438
rect 586658 705202 586840 705438
rect 580404 689818 580586 690054
rect 580822 689818 581004 690054
rect 580404 689734 581004 689818
rect 580404 689498 580586 689734
rect 580822 689498 581004 689734
rect 580404 654054 581004 689498
rect 580404 653818 580586 654054
rect 580822 653818 581004 654054
rect 580404 653734 581004 653818
rect 580404 653498 580586 653734
rect 580822 653498 581004 653734
rect 580404 618054 581004 653498
rect 580404 617818 580586 618054
rect 580822 617818 581004 618054
rect 580404 617734 581004 617818
rect 580404 617498 580586 617734
rect 580822 617498 581004 617734
rect 580404 582054 581004 617498
rect 580404 581818 580586 582054
rect 580822 581818 581004 582054
rect 580404 581734 581004 581818
rect 580404 581498 580586 581734
rect 580822 581498 581004 581734
rect 580404 546054 581004 581498
rect 580404 545818 580586 546054
rect 580822 545818 581004 546054
rect 580404 545734 581004 545818
rect 580404 545498 580586 545734
rect 580822 545498 581004 545734
rect 580404 510054 581004 545498
rect 580404 509818 580586 510054
rect 580822 509818 581004 510054
rect 580404 509734 581004 509818
rect 580404 509498 580586 509734
rect 580822 509498 581004 509734
rect 580404 474054 581004 509498
rect 580404 473818 580586 474054
rect 580822 473818 581004 474054
rect 580404 473734 581004 473818
rect 580404 473498 580586 473734
rect 580822 473498 581004 473734
rect 580404 438054 581004 473498
rect 580404 437818 580586 438054
rect 580822 437818 581004 438054
rect 580404 437734 581004 437818
rect 580404 437498 580586 437734
rect 580822 437498 581004 437734
rect 580404 402054 581004 437498
rect 580404 401818 580586 402054
rect 580822 401818 581004 402054
rect 580404 401734 581004 401818
rect 580404 401498 580586 401734
rect 580822 401498 581004 401734
rect 580404 366054 581004 401498
rect 580404 365818 580586 366054
rect 580822 365818 581004 366054
rect 580404 365734 581004 365818
rect 580404 365498 580586 365734
rect 580822 365498 581004 365734
rect 580404 330054 581004 365498
rect 580404 329818 580586 330054
rect 580822 329818 581004 330054
rect 580404 329734 581004 329818
rect 580404 329498 580586 329734
rect 580822 329498 581004 329734
rect 580404 294054 581004 329498
rect 580404 293818 580586 294054
rect 580822 293818 581004 294054
rect 580404 293734 581004 293818
rect 580404 293498 580586 293734
rect 580822 293498 581004 293734
rect 580404 258054 581004 293498
rect 580404 257818 580586 258054
rect 580822 257818 581004 258054
rect 580404 257734 581004 257818
rect 580404 257498 580586 257734
rect 580822 257498 581004 257734
rect 580404 222054 581004 257498
rect 580404 221818 580586 222054
rect 580822 221818 581004 222054
rect 580404 221734 581004 221818
rect 580404 221498 580586 221734
rect 580822 221498 581004 221734
rect 580404 186054 581004 221498
rect 580404 185818 580586 186054
rect 580822 185818 581004 186054
rect 580404 185734 581004 185818
rect 580404 185498 580586 185734
rect 580822 185498 581004 185734
rect 580404 150054 581004 185498
rect 580404 149818 580586 150054
rect 580822 149818 581004 150054
rect 580404 149734 581004 149818
rect 580404 149498 580586 149734
rect 580822 149498 581004 149734
rect 580404 114054 581004 149498
rect 580404 113818 580586 114054
rect 580822 113818 581004 114054
rect 580404 113734 581004 113818
rect 580404 113498 580586 113734
rect 580822 113498 581004 113734
rect 580404 78054 581004 113498
rect 580404 77818 580586 78054
rect 580822 77818 581004 78054
rect 580404 77734 581004 77818
rect 580404 77498 580586 77734
rect 580822 77498 581004 77734
rect 580404 42054 581004 77498
rect 580404 41818 580586 42054
rect 580822 41818 581004 42054
rect 580404 41734 581004 41818
rect 580404 41498 580586 41734
rect 580822 41498 581004 41734
rect 580404 6054 581004 41498
rect 580404 5818 580586 6054
rect 580822 5818 581004 6054
rect 580404 5734 581004 5818
rect 580404 5498 580586 5734
rect 580822 5498 581004 5734
rect 580404 -2186 581004 5498
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 686454 585920 704282
rect 585320 686218 585502 686454
rect 585738 686218 585920 686454
rect 585320 686134 585920 686218
rect 585320 685898 585502 686134
rect 585738 685898 585920 686134
rect 585320 650454 585920 685898
rect 585320 650218 585502 650454
rect 585738 650218 585920 650454
rect 585320 650134 585920 650218
rect 585320 649898 585502 650134
rect 585738 649898 585920 650134
rect 585320 614454 585920 649898
rect 585320 614218 585502 614454
rect 585738 614218 585920 614454
rect 585320 614134 585920 614218
rect 585320 613898 585502 614134
rect 585738 613898 585920 614134
rect 585320 578454 585920 613898
rect 585320 578218 585502 578454
rect 585738 578218 585920 578454
rect 585320 578134 585920 578218
rect 585320 577898 585502 578134
rect 585738 577898 585920 578134
rect 585320 542454 585920 577898
rect 585320 542218 585502 542454
rect 585738 542218 585920 542454
rect 585320 542134 585920 542218
rect 585320 541898 585502 542134
rect 585738 541898 585920 542134
rect 585320 506454 585920 541898
rect 585320 506218 585502 506454
rect 585738 506218 585920 506454
rect 585320 506134 585920 506218
rect 585320 505898 585502 506134
rect 585738 505898 585920 506134
rect 585320 470454 585920 505898
rect 585320 470218 585502 470454
rect 585738 470218 585920 470454
rect 585320 470134 585920 470218
rect 585320 469898 585502 470134
rect 585738 469898 585920 470134
rect 585320 434454 585920 469898
rect 585320 434218 585502 434454
rect 585738 434218 585920 434454
rect 585320 434134 585920 434218
rect 585320 433898 585502 434134
rect 585738 433898 585920 434134
rect 585320 398454 585920 433898
rect 585320 398218 585502 398454
rect 585738 398218 585920 398454
rect 585320 398134 585920 398218
rect 585320 397898 585502 398134
rect 585738 397898 585920 398134
rect 585320 362454 585920 397898
rect 585320 362218 585502 362454
rect 585738 362218 585920 362454
rect 585320 362134 585920 362218
rect 585320 361898 585502 362134
rect 585738 361898 585920 362134
rect 585320 326454 585920 361898
rect 585320 326218 585502 326454
rect 585738 326218 585920 326454
rect 585320 326134 585920 326218
rect 585320 325898 585502 326134
rect 585738 325898 585920 326134
rect 585320 290454 585920 325898
rect 585320 290218 585502 290454
rect 585738 290218 585920 290454
rect 585320 290134 585920 290218
rect 585320 289898 585502 290134
rect 585738 289898 585920 290134
rect 585320 254454 585920 289898
rect 585320 254218 585502 254454
rect 585738 254218 585920 254454
rect 585320 254134 585920 254218
rect 585320 253898 585502 254134
rect 585738 253898 585920 254134
rect 585320 218454 585920 253898
rect 585320 218218 585502 218454
rect 585738 218218 585920 218454
rect 585320 218134 585920 218218
rect 585320 217898 585502 218134
rect 585738 217898 585920 218134
rect 585320 182454 585920 217898
rect 585320 182218 585502 182454
rect 585738 182218 585920 182454
rect 585320 182134 585920 182218
rect 585320 181898 585502 182134
rect 585738 181898 585920 182134
rect 585320 146454 585920 181898
rect 585320 146218 585502 146454
rect 585738 146218 585920 146454
rect 585320 146134 585920 146218
rect 585320 145898 585502 146134
rect 585738 145898 585920 146134
rect 585320 110454 585920 145898
rect 585320 110218 585502 110454
rect 585738 110218 585920 110454
rect 585320 110134 585920 110218
rect 585320 109898 585502 110134
rect 585738 109898 585920 110134
rect 585320 74454 585920 109898
rect 585320 74218 585502 74454
rect 585738 74218 585920 74454
rect 585320 74134 585920 74218
rect 585320 73898 585502 74134
rect 585738 73898 585920 74134
rect 585320 38454 585920 73898
rect 585320 38218 585502 38454
rect 585738 38218 585920 38454
rect 585320 38134 585920 38218
rect 585320 37898 585502 38134
rect 585738 37898 585920 38134
rect 585320 2454 585920 37898
rect 585320 2218 585502 2454
rect 585738 2218 585920 2454
rect 585320 2134 585920 2218
rect 585320 1898 585502 2134
rect 585738 1898 585920 2134
rect 585320 -346 585920 1898
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586240 668454 586840 705202
rect 586240 668218 586422 668454
rect 586658 668218 586840 668454
rect 586240 668134 586840 668218
rect 586240 667898 586422 668134
rect 586658 667898 586840 668134
rect 586240 632454 586840 667898
rect 586240 632218 586422 632454
rect 586658 632218 586840 632454
rect 586240 632134 586840 632218
rect 586240 631898 586422 632134
rect 586658 631898 586840 632134
rect 586240 596454 586840 631898
rect 586240 596218 586422 596454
rect 586658 596218 586840 596454
rect 586240 596134 586840 596218
rect 586240 595898 586422 596134
rect 586658 595898 586840 596134
rect 586240 560454 586840 595898
rect 586240 560218 586422 560454
rect 586658 560218 586840 560454
rect 586240 560134 586840 560218
rect 586240 559898 586422 560134
rect 586658 559898 586840 560134
rect 586240 524454 586840 559898
rect 586240 524218 586422 524454
rect 586658 524218 586840 524454
rect 586240 524134 586840 524218
rect 586240 523898 586422 524134
rect 586658 523898 586840 524134
rect 586240 488454 586840 523898
rect 586240 488218 586422 488454
rect 586658 488218 586840 488454
rect 586240 488134 586840 488218
rect 586240 487898 586422 488134
rect 586658 487898 586840 488134
rect 586240 452454 586840 487898
rect 586240 452218 586422 452454
rect 586658 452218 586840 452454
rect 586240 452134 586840 452218
rect 586240 451898 586422 452134
rect 586658 451898 586840 452134
rect 586240 416454 586840 451898
rect 586240 416218 586422 416454
rect 586658 416218 586840 416454
rect 586240 416134 586840 416218
rect 586240 415898 586422 416134
rect 586658 415898 586840 416134
rect 586240 380454 586840 415898
rect 586240 380218 586422 380454
rect 586658 380218 586840 380454
rect 586240 380134 586840 380218
rect 586240 379898 586422 380134
rect 586658 379898 586840 380134
rect 586240 344454 586840 379898
rect 586240 344218 586422 344454
rect 586658 344218 586840 344454
rect 586240 344134 586840 344218
rect 586240 343898 586422 344134
rect 586658 343898 586840 344134
rect 586240 308454 586840 343898
rect 586240 308218 586422 308454
rect 586658 308218 586840 308454
rect 586240 308134 586840 308218
rect 586240 307898 586422 308134
rect 586658 307898 586840 308134
rect 586240 272454 586840 307898
rect 586240 272218 586422 272454
rect 586658 272218 586840 272454
rect 586240 272134 586840 272218
rect 586240 271898 586422 272134
rect 586658 271898 586840 272134
rect 586240 236454 586840 271898
rect 586240 236218 586422 236454
rect 586658 236218 586840 236454
rect 586240 236134 586840 236218
rect 586240 235898 586422 236134
rect 586658 235898 586840 236134
rect 586240 200454 586840 235898
rect 586240 200218 586422 200454
rect 586658 200218 586840 200454
rect 586240 200134 586840 200218
rect 586240 199898 586422 200134
rect 586658 199898 586840 200134
rect 586240 164454 586840 199898
rect 586240 164218 586422 164454
rect 586658 164218 586840 164454
rect 586240 164134 586840 164218
rect 586240 163898 586422 164134
rect 586658 163898 586840 164134
rect 586240 128454 586840 163898
rect 586240 128218 586422 128454
rect 586658 128218 586840 128454
rect 586240 128134 586840 128218
rect 586240 127898 586422 128134
rect 586658 127898 586840 128134
rect 586240 92454 586840 127898
rect 586240 92218 586422 92454
rect 586658 92218 586840 92454
rect 586240 92134 586840 92218
rect 586240 91898 586422 92134
rect 586658 91898 586840 92134
rect 586240 56454 586840 91898
rect 586240 56218 586422 56454
rect 586658 56218 586840 56454
rect 586240 56134 586840 56218
rect 586240 55898 586422 56134
rect 586658 55898 586840 56134
rect 586240 20454 586840 55898
rect 586240 20218 586422 20454
rect 586658 20218 586840 20454
rect 586240 20134 586840 20218
rect 586240 19898 586422 20134
rect 586658 19898 586840 20134
rect 586240 -1266 586840 19898
rect 586240 -1502 586422 -1266
rect 586658 -1502 586840 -1266
rect 586240 -1586 586840 -1502
rect 586240 -1822 586422 -1586
rect 586658 -1822 586840 -1586
rect 586240 -1844 586840 -1822
rect 587160 690054 587760 706122
rect 587160 689818 587342 690054
rect 587578 689818 587760 690054
rect 587160 689734 587760 689818
rect 587160 689498 587342 689734
rect 587578 689498 587760 689734
rect 587160 654054 587760 689498
rect 587160 653818 587342 654054
rect 587578 653818 587760 654054
rect 587160 653734 587760 653818
rect 587160 653498 587342 653734
rect 587578 653498 587760 653734
rect 587160 618054 587760 653498
rect 587160 617818 587342 618054
rect 587578 617818 587760 618054
rect 587160 617734 587760 617818
rect 587160 617498 587342 617734
rect 587578 617498 587760 617734
rect 587160 582054 587760 617498
rect 587160 581818 587342 582054
rect 587578 581818 587760 582054
rect 587160 581734 587760 581818
rect 587160 581498 587342 581734
rect 587578 581498 587760 581734
rect 587160 546054 587760 581498
rect 587160 545818 587342 546054
rect 587578 545818 587760 546054
rect 587160 545734 587760 545818
rect 587160 545498 587342 545734
rect 587578 545498 587760 545734
rect 587160 510054 587760 545498
rect 587160 509818 587342 510054
rect 587578 509818 587760 510054
rect 587160 509734 587760 509818
rect 587160 509498 587342 509734
rect 587578 509498 587760 509734
rect 587160 474054 587760 509498
rect 587160 473818 587342 474054
rect 587578 473818 587760 474054
rect 587160 473734 587760 473818
rect 587160 473498 587342 473734
rect 587578 473498 587760 473734
rect 587160 438054 587760 473498
rect 587160 437818 587342 438054
rect 587578 437818 587760 438054
rect 587160 437734 587760 437818
rect 587160 437498 587342 437734
rect 587578 437498 587760 437734
rect 587160 402054 587760 437498
rect 587160 401818 587342 402054
rect 587578 401818 587760 402054
rect 587160 401734 587760 401818
rect 587160 401498 587342 401734
rect 587578 401498 587760 401734
rect 587160 366054 587760 401498
rect 587160 365818 587342 366054
rect 587578 365818 587760 366054
rect 587160 365734 587760 365818
rect 587160 365498 587342 365734
rect 587578 365498 587760 365734
rect 587160 330054 587760 365498
rect 587160 329818 587342 330054
rect 587578 329818 587760 330054
rect 587160 329734 587760 329818
rect 587160 329498 587342 329734
rect 587578 329498 587760 329734
rect 587160 294054 587760 329498
rect 587160 293818 587342 294054
rect 587578 293818 587760 294054
rect 587160 293734 587760 293818
rect 587160 293498 587342 293734
rect 587578 293498 587760 293734
rect 587160 258054 587760 293498
rect 587160 257818 587342 258054
rect 587578 257818 587760 258054
rect 587160 257734 587760 257818
rect 587160 257498 587342 257734
rect 587578 257498 587760 257734
rect 587160 222054 587760 257498
rect 587160 221818 587342 222054
rect 587578 221818 587760 222054
rect 587160 221734 587760 221818
rect 587160 221498 587342 221734
rect 587578 221498 587760 221734
rect 587160 186054 587760 221498
rect 587160 185818 587342 186054
rect 587578 185818 587760 186054
rect 587160 185734 587760 185818
rect 587160 185498 587342 185734
rect 587578 185498 587760 185734
rect 587160 150054 587760 185498
rect 587160 149818 587342 150054
rect 587578 149818 587760 150054
rect 587160 149734 587760 149818
rect 587160 149498 587342 149734
rect 587578 149498 587760 149734
rect 587160 114054 587760 149498
rect 587160 113818 587342 114054
rect 587578 113818 587760 114054
rect 587160 113734 587760 113818
rect 587160 113498 587342 113734
rect 587578 113498 587760 113734
rect 587160 78054 587760 113498
rect 587160 77818 587342 78054
rect 587578 77818 587760 78054
rect 587160 77734 587760 77818
rect 587160 77498 587342 77734
rect 587578 77498 587760 77734
rect 587160 42054 587760 77498
rect 587160 41818 587342 42054
rect 587578 41818 587760 42054
rect 587160 41734 587760 41818
rect 587160 41498 587342 41734
rect 587578 41498 587760 41734
rect 587160 6054 587760 41498
rect 587160 5818 587342 6054
rect 587578 5818 587760 6054
rect 587160 5734 587760 5818
rect 587160 5498 587342 5734
rect 587578 5498 587760 5734
rect 580404 -2422 580586 -2186
rect 580822 -2422 581004 -2186
rect 580404 -2506 581004 -2422
rect 580404 -2742 580586 -2506
rect 580822 -2742 581004 -2506
rect 580404 -3684 581004 -2742
rect 587160 -2186 587760 5498
rect 587160 -2422 587342 -2186
rect 587578 -2422 587760 -2186
rect 587160 -2506 587760 -2422
rect 587160 -2742 587342 -2506
rect 587578 -2742 587760 -2506
rect 587160 -2764 587760 -2742
rect 588080 672054 588680 707042
rect 588080 671818 588262 672054
rect 588498 671818 588680 672054
rect 588080 671734 588680 671818
rect 588080 671498 588262 671734
rect 588498 671498 588680 671734
rect 588080 636054 588680 671498
rect 588080 635818 588262 636054
rect 588498 635818 588680 636054
rect 588080 635734 588680 635818
rect 588080 635498 588262 635734
rect 588498 635498 588680 635734
rect 588080 600054 588680 635498
rect 588080 599818 588262 600054
rect 588498 599818 588680 600054
rect 588080 599734 588680 599818
rect 588080 599498 588262 599734
rect 588498 599498 588680 599734
rect 588080 564054 588680 599498
rect 588080 563818 588262 564054
rect 588498 563818 588680 564054
rect 588080 563734 588680 563818
rect 588080 563498 588262 563734
rect 588498 563498 588680 563734
rect 588080 528054 588680 563498
rect 588080 527818 588262 528054
rect 588498 527818 588680 528054
rect 588080 527734 588680 527818
rect 588080 527498 588262 527734
rect 588498 527498 588680 527734
rect 588080 492054 588680 527498
rect 588080 491818 588262 492054
rect 588498 491818 588680 492054
rect 588080 491734 588680 491818
rect 588080 491498 588262 491734
rect 588498 491498 588680 491734
rect 588080 456054 588680 491498
rect 588080 455818 588262 456054
rect 588498 455818 588680 456054
rect 588080 455734 588680 455818
rect 588080 455498 588262 455734
rect 588498 455498 588680 455734
rect 588080 420054 588680 455498
rect 588080 419818 588262 420054
rect 588498 419818 588680 420054
rect 588080 419734 588680 419818
rect 588080 419498 588262 419734
rect 588498 419498 588680 419734
rect 588080 384054 588680 419498
rect 588080 383818 588262 384054
rect 588498 383818 588680 384054
rect 588080 383734 588680 383818
rect 588080 383498 588262 383734
rect 588498 383498 588680 383734
rect 588080 348054 588680 383498
rect 588080 347818 588262 348054
rect 588498 347818 588680 348054
rect 588080 347734 588680 347818
rect 588080 347498 588262 347734
rect 588498 347498 588680 347734
rect 588080 312054 588680 347498
rect 588080 311818 588262 312054
rect 588498 311818 588680 312054
rect 588080 311734 588680 311818
rect 588080 311498 588262 311734
rect 588498 311498 588680 311734
rect 588080 276054 588680 311498
rect 588080 275818 588262 276054
rect 588498 275818 588680 276054
rect 588080 275734 588680 275818
rect 588080 275498 588262 275734
rect 588498 275498 588680 275734
rect 588080 240054 588680 275498
rect 588080 239818 588262 240054
rect 588498 239818 588680 240054
rect 588080 239734 588680 239818
rect 588080 239498 588262 239734
rect 588498 239498 588680 239734
rect 588080 204054 588680 239498
rect 588080 203818 588262 204054
rect 588498 203818 588680 204054
rect 588080 203734 588680 203818
rect 588080 203498 588262 203734
rect 588498 203498 588680 203734
rect 588080 168054 588680 203498
rect 588080 167818 588262 168054
rect 588498 167818 588680 168054
rect 588080 167734 588680 167818
rect 588080 167498 588262 167734
rect 588498 167498 588680 167734
rect 588080 132054 588680 167498
rect 588080 131818 588262 132054
rect 588498 131818 588680 132054
rect 588080 131734 588680 131818
rect 588080 131498 588262 131734
rect 588498 131498 588680 131734
rect 588080 96054 588680 131498
rect 588080 95818 588262 96054
rect 588498 95818 588680 96054
rect 588080 95734 588680 95818
rect 588080 95498 588262 95734
rect 588498 95498 588680 95734
rect 588080 60054 588680 95498
rect 588080 59818 588262 60054
rect 588498 59818 588680 60054
rect 588080 59734 588680 59818
rect 588080 59498 588262 59734
rect 588498 59498 588680 59734
rect 588080 24054 588680 59498
rect 588080 23818 588262 24054
rect 588498 23818 588680 24054
rect 588080 23734 588680 23818
rect 588080 23498 588262 23734
rect 588498 23498 588680 23734
rect 588080 -3106 588680 23498
rect 588080 -3342 588262 -3106
rect 588498 -3342 588680 -3106
rect 588080 -3426 588680 -3342
rect 588080 -3662 588262 -3426
rect 588498 -3662 588680 -3426
rect 588080 -3684 588680 -3662
rect 589000 693654 589600 707962
rect 589000 693418 589182 693654
rect 589418 693418 589600 693654
rect 589000 693334 589600 693418
rect 589000 693098 589182 693334
rect 589418 693098 589600 693334
rect 589000 657654 589600 693098
rect 589000 657418 589182 657654
rect 589418 657418 589600 657654
rect 589000 657334 589600 657418
rect 589000 657098 589182 657334
rect 589418 657098 589600 657334
rect 589000 621654 589600 657098
rect 589000 621418 589182 621654
rect 589418 621418 589600 621654
rect 589000 621334 589600 621418
rect 589000 621098 589182 621334
rect 589418 621098 589600 621334
rect 589000 585654 589600 621098
rect 589000 585418 589182 585654
rect 589418 585418 589600 585654
rect 589000 585334 589600 585418
rect 589000 585098 589182 585334
rect 589418 585098 589600 585334
rect 589000 549654 589600 585098
rect 589000 549418 589182 549654
rect 589418 549418 589600 549654
rect 589000 549334 589600 549418
rect 589000 549098 589182 549334
rect 589418 549098 589600 549334
rect 589000 513654 589600 549098
rect 589000 513418 589182 513654
rect 589418 513418 589600 513654
rect 589000 513334 589600 513418
rect 589000 513098 589182 513334
rect 589418 513098 589600 513334
rect 589000 477654 589600 513098
rect 589000 477418 589182 477654
rect 589418 477418 589600 477654
rect 589000 477334 589600 477418
rect 589000 477098 589182 477334
rect 589418 477098 589600 477334
rect 589000 441654 589600 477098
rect 589000 441418 589182 441654
rect 589418 441418 589600 441654
rect 589000 441334 589600 441418
rect 589000 441098 589182 441334
rect 589418 441098 589600 441334
rect 589000 405654 589600 441098
rect 589000 405418 589182 405654
rect 589418 405418 589600 405654
rect 589000 405334 589600 405418
rect 589000 405098 589182 405334
rect 589418 405098 589600 405334
rect 589000 369654 589600 405098
rect 589000 369418 589182 369654
rect 589418 369418 589600 369654
rect 589000 369334 589600 369418
rect 589000 369098 589182 369334
rect 589418 369098 589600 369334
rect 589000 333654 589600 369098
rect 589000 333418 589182 333654
rect 589418 333418 589600 333654
rect 589000 333334 589600 333418
rect 589000 333098 589182 333334
rect 589418 333098 589600 333334
rect 589000 297654 589600 333098
rect 589000 297418 589182 297654
rect 589418 297418 589600 297654
rect 589000 297334 589600 297418
rect 589000 297098 589182 297334
rect 589418 297098 589600 297334
rect 589000 261654 589600 297098
rect 589000 261418 589182 261654
rect 589418 261418 589600 261654
rect 589000 261334 589600 261418
rect 589000 261098 589182 261334
rect 589418 261098 589600 261334
rect 589000 225654 589600 261098
rect 589000 225418 589182 225654
rect 589418 225418 589600 225654
rect 589000 225334 589600 225418
rect 589000 225098 589182 225334
rect 589418 225098 589600 225334
rect 589000 189654 589600 225098
rect 589000 189418 589182 189654
rect 589418 189418 589600 189654
rect 589000 189334 589600 189418
rect 589000 189098 589182 189334
rect 589418 189098 589600 189334
rect 589000 153654 589600 189098
rect 589000 153418 589182 153654
rect 589418 153418 589600 153654
rect 589000 153334 589600 153418
rect 589000 153098 589182 153334
rect 589418 153098 589600 153334
rect 589000 117654 589600 153098
rect 589000 117418 589182 117654
rect 589418 117418 589600 117654
rect 589000 117334 589600 117418
rect 589000 117098 589182 117334
rect 589418 117098 589600 117334
rect 589000 81654 589600 117098
rect 589000 81418 589182 81654
rect 589418 81418 589600 81654
rect 589000 81334 589600 81418
rect 589000 81098 589182 81334
rect 589418 81098 589600 81334
rect 589000 45654 589600 81098
rect 589000 45418 589182 45654
rect 589418 45418 589600 45654
rect 589000 45334 589600 45418
rect 589000 45098 589182 45334
rect 589418 45098 589600 45334
rect 589000 9654 589600 45098
rect 589000 9418 589182 9654
rect 589418 9418 589600 9654
rect 589000 9334 589600 9418
rect 589000 9098 589182 9334
rect 589418 9098 589600 9334
rect 589000 -4026 589600 9098
rect 589000 -4262 589182 -4026
rect 589418 -4262 589600 -4026
rect 589000 -4346 589600 -4262
rect 589000 -4582 589182 -4346
rect 589418 -4582 589600 -4346
rect 589000 -4604 589600 -4582
rect 589920 675654 590520 708882
rect 589920 675418 590102 675654
rect 590338 675418 590520 675654
rect 589920 675334 590520 675418
rect 589920 675098 590102 675334
rect 590338 675098 590520 675334
rect 589920 639654 590520 675098
rect 589920 639418 590102 639654
rect 590338 639418 590520 639654
rect 589920 639334 590520 639418
rect 589920 639098 590102 639334
rect 590338 639098 590520 639334
rect 589920 603654 590520 639098
rect 589920 603418 590102 603654
rect 590338 603418 590520 603654
rect 589920 603334 590520 603418
rect 589920 603098 590102 603334
rect 590338 603098 590520 603334
rect 589920 567654 590520 603098
rect 589920 567418 590102 567654
rect 590338 567418 590520 567654
rect 589920 567334 590520 567418
rect 589920 567098 590102 567334
rect 590338 567098 590520 567334
rect 589920 531654 590520 567098
rect 589920 531418 590102 531654
rect 590338 531418 590520 531654
rect 589920 531334 590520 531418
rect 589920 531098 590102 531334
rect 590338 531098 590520 531334
rect 589920 495654 590520 531098
rect 589920 495418 590102 495654
rect 590338 495418 590520 495654
rect 589920 495334 590520 495418
rect 589920 495098 590102 495334
rect 590338 495098 590520 495334
rect 589920 459654 590520 495098
rect 589920 459418 590102 459654
rect 590338 459418 590520 459654
rect 589920 459334 590520 459418
rect 589920 459098 590102 459334
rect 590338 459098 590520 459334
rect 589920 423654 590520 459098
rect 589920 423418 590102 423654
rect 590338 423418 590520 423654
rect 589920 423334 590520 423418
rect 589920 423098 590102 423334
rect 590338 423098 590520 423334
rect 589920 387654 590520 423098
rect 589920 387418 590102 387654
rect 590338 387418 590520 387654
rect 589920 387334 590520 387418
rect 589920 387098 590102 387334
rect 590338 387098 590520 387334
rect 589920 351654 590520 387098
rect 589920 351418 590102 351654
rect 590338 351418 590520 351654
rect 589920 351334 590520 351418
rect 589920 351098 590102 351334
rect 590338 351098 590520 351334
rect 589920 315654 590520 351098
rect 589920 315418 590102 315654
rect 590338 315418 590520 315654
rect 589920 315334 590520 315418
rect 589920 315098 590102 315334
rect 590338 315098 590520 315334
rect 589920 279654 590520 315098
rect 589920 279418 590102 279654
rect 590338 279418 590520 279654
rect 589920 279334 590520 279418
rect 589920 279098 590102 279334
rect 590338 279098 590520 279334
rect 589920 243654 590520 279098
rect 589920 243418 590102 243654
rect 590338 243418 590520 243654
rect 589920 243334 590520 243418
rect 589920 243098 590102 243334
rect 590338 243098 590520 243334
rect 589920 207654 590520 243098
rect 589920 207418 590102 207654
rect 590338 207418 590520 207654
rect 589920 207334 590520 207418
rect 589920 207098 590102 207334
rect 590338 207098 590520 207334
rect 589920 171654 590520 207098
rect 589920 171418 590102 171654
rect 590338 171418 590520 171654
rect 589920 171334 590520 171418
rect 589920 171098 590102 171334
rect 590338 171098 590520 171334
rect 589920 135654 590520 171098
rect 589920 135418 590102 135654
rect 590338 135418 590520 135654
rect 589920 135334 590520 135418
rect 589920 135098 590102 135334
rect 590338 135098 590520 135334
rect 589920 99654 590520 135098
rect 589920 99418 590102 99654
rect 590338 99418 590520 99654
rect 589920 99334 590520 99418
rect 589920 99098 590102 99334
rect 590338 99098 590520 99334
rect 589920 63654 590520 99098
rect 589920 63418 590102 63654
rect 590338 63418 590520 63654
rect 589920 63334 590520 63418
rect 589920 63098 590102 63334
rect 590338 63098 590520 63334
rect 589920 27654 590520 63098
rect 589920 27418 590102 27654
rect 590338 27418 590520 27654
rect 589920 27334 590520 27418
rect 589920 27098 590102 27334
rect 590338 27098 590520 27334
rect 589920 -4946 590520 27098
rect 589920 -5182 590102 -4946
rect 590338 -5182 590520 -4946
rect 589920 -5266 590520 -5182
rect 589920 -5502 590102 -5266
rect 590338 -5502 590520 -5266
rect 589920 -5524 590520 -5502
rect 590840 697254 591440 709802
rect 590840 697018 591022 697254
rect 591258 697018 591440 697254
rect 590840 696934 591440 697018
rect 590840 696698 591022 696934
rect 591258 696698 591440 696934
rect 590840 661254 591440 696698
rect 590840 661018 591022 661254
rect 591258 661018 591440 661254
rect 590840 660934 591440 661018
rect 590840 660698 591022 660934
rect 591258 660698 591440 660934
rect 590840 625254 591440 660698
rect 590840 625018 591022 625254
rect 591258 625018 591440 625254
rect 590840 624934 591440 625018
rect 590840 624698 591022 624934
rect 591258 624698 591440 624934
rect 590840 589254 591440 624698
rect 590840 589018 591022 589254
rect 591258 589018 591440 589254
rect 590840 588934 591440 589018
rect 590840 588698 591022 588934
rect 591258 588698 591440 588934
rect 590840 553254 591440 588698
rect 590840 553018 591022 553254
rect 591258 553018 591440 553254
rect 590840 552934 591440 553018
rect 590840 552698 591022 552934
rect 591258 552698 591440 552934
rect 590840 517254 591440 552698
rect 590840 517018 591022 517254
rect 591258 517018 591440 517254
rect 590840 516934 591440 517018
rect 590840 516698 591022 516934
rect 591258 516698 591440 516934
rect 590840 481254 591440 516698
rect 590840 481018 591022 481254
rect 591258 481018 591440 481254
rect 590840 480934 591440 481018
rect 590840 480698 591022 480934
rect 591258 480698 591440 480934
rect 590840 445254 591440 480698
rect 590840 445018 591022 445254
rect 591258 445018 591440 445254
rect 590840 444934 591440 445018
rect 590840 444698 591022 444934
rect 591258 444698 591440 444934
rect 590840 409254 591440 444698
rect 590840 409018 591022 409254
rect 591258 409018 591440 409254
rect 590840 408934 591440 409018
rect 590840 408698 591022 408934
rect 591258 408698 591440 408934
rect 590840 373254 591440 408698
rect 590840 373018 591022 373254
rect 591258 373018 591440 373254
rect 590840 372934 591440 373018
rect 590840 372698 591022 372934
rect 591258 372698 591440 372934
rect 590840 337254 591440 372698
rect 590840 337018 591022 337254
rect 591258 337018 591440 337254
rect 590840 336934 591440 337018
rect 590840 336698 591022 336934
rect 591258 336698 591440 336934
rect 590840 301254 591440 336698
rect 590840 301018 591022 301254
rect 591258 301018 591440 301254
rect 590840 300934 591440 301018
rect 590840 300698 591022 300934
rect 591258 300698 591440 300934
rect 590840 265254 591440 300698
rect 590840 265018 591022 265254
rect 591258 265018 591440 265254
rect 590840 264934 591440 265018
rect 590840 264698 591022 264934
rect 591258 264698 591440 264934
rect 590840 229254 591440 264698
rect 590840 229018 591022 229254
rect 591258 229018 591440 229254
rect 590840 228934 591440 229018
rect 590840 228698 591022 228934
rect 591258 228698 591440 228934
rect 590840 193254 591440 228698
rect 590840 193018 591022 193254
rect 591258 193018 591440 193254
rect 590840 192934 591440 193018
rect 590840 192698 591022 192934
rect 591258 192698 591440 192934
rect 590840 157254 591440 192698
rect 590840 157018 591022 157254
rect 591258 157018 591440 157254
rect 590840 156934 591440 157018
rect 590840 156698 591022 156934
rect 591258 156698 591440 156934
rect 590840 121254 591440 156698
rect 590840 121018 591022 121254
rect 591258 121018 591440 121254
rect 590840 120934 591440 121018
rect 590840 120698 591022 120934
rect 591258 120698 591440 120934
rect 590840 85254 591440 120698
rect 590840 85018 591022 85254
rect 591258 85018 591440 85254
rect 590840 84934 591440 85018
rect 590840 84698 591022 84934
rect 591258 84698 591440 84934
rect 590840 49254 591440 84698
rect 590840 49018 591022 49254
rect 591258 49018 591440 49254
rect 590840 48934 591440 49018
rect 590840 48698 591022 48934
rect 591258 48698 591440 48934
rect 590840 13254 591440 48698
rect 590840 13018 591022 13254
rect 591258 13018 591440 13254
rect 590840 12934 591440 13018
rect 590840 12698 591022 12934
rect 591258 12698 591440 12934
rect 590840 -5866 591440 12698
rect 590840 -6102 591022 -5866
rect 591258 -6102 591440 -5866
rect 590840 -6186 591440 -6102
rect 590840 -6422 591022 -6186
rect 591258 -6422 591440 -6186
rect 590840 -6444 591440 -6422
rect 591760 679254 592360 710722
rect 591760 679018 591942 679254
rect 592178 679018 592360 679254
rect 591760 678934 592360 679018
rect 591760 678698 591942 678934
rect 592178 678698 592360 678934
rect 591760 643254 592360 678698
rect 591760 643018 591942 643254
rect 592178 643018 592360 643254
rect 591760 642934 592360 643018
rect 591760 642698 591942 642934
rect 592178 642698 592360 642934
rect 591760 607254 592360 642698
rect 591760 607018 591942 607254
rect 592178 607018 592360 607254
rect 591760 606934 592360 607018
rect 591760 606698 591942 606934
rect 592178 606698 592360 606934
rect 591760 571254 592360 606698
rect 591760 571018 591942 571254
rect 592178 571018 592360 571254
rect 591760 570934 592360 571018
rect 591760 570698 591942 570934
rect 592178 570698 592360 570934
rect 591760 535254 592360 570698
rect 591760 535018 591942 535254
rect 592178 535018 592360 535254
rect 591760 534934 592360 535018
rect 591760 534698 591942 534934
rect 592178 534698 592360 534934
rect 591760 499254 592360 534698
rect 591760 499018 591942 499254
rect 592178 499018 592360 499254
rect 591760 498934 592360 499018
rect 591760 498698 591942 498934
rect 592178 498698 592360 498934
rect 591760 463254 592360 498698
rect 591760 463018 591942 463254
rect 592178 463018 592360 463254
rect 591760 462934 592360 463018
rect 591760 462698 591942 462934
rect 592178 462698 592360 462934
rect 591760 427254 592360 462698
rect 591760 427018 591942 427254
rect 592178 427018 592360 427254
rect 591760 426934 592360 427018
rect 591760 426698 591942 426934
rect 592178 426698 592360 426934
rect 591760 391254 592360 426698
rect 591760 391018 591942 391254
rect 592178 391018 592360 391254
rect 591760 390934 592360 391018
rect 591760 390698 591942 390934
rect 592178 390698 592360 390934
rect 591760 355254 592360 390698
rect 591760 355018 591942 355254
rect 592178 355018 592360 355254
rect 591760 354934 592360 355018
rect 591760 354698 591942 354934
rect 592178 354698 592360 354934
rect 591760 319254 592360 354698
rect 591760 319018 591942 319254
rect 592178 319018 592360 319254
rect 591760 318934 592360 319018
rect 591760 318698 591942 318934
rect 592178 318698 592360 318934
rect 591760 283254 592360 318698
rect 591760 283018 591942 283254
rect 592178 283018 592360 283254
rect 591760 282934 592360 283018
rect 591760 282698 591942 282934
rect 592178 282698 592360 282934
rect 591760 247254 592360 282698
rect 591760 247018 591942 247254
rect 592178 247018 592360 247254
rect 591760 246934 592360 247018
rect 591760 246698 591942 246934
rect 592178 246698 592360 246934
rect 591760 211254 592360 246698
rect 591760 211018 591942 211254
rect 592178 211018 592360 211254
rect 591760 210934 592360 211018
rect 591760 210698 591942 210934
rect 592178 210698 592360 210934
rect 591760 175254 592360 210698
rect 591760 175018 591942 175254
rect 592178 175018 592360 175254
rect 591760 174934 592360 175018
rect 591760 174698 591942 174934
rect 592178 174698 592360 174934
rect 591760 139254 592360 174698
rect 591760 139018 591942 139254
rect 592178 139018 592360 139254
rect 591760 138934 592360 139018
rect 591760 138698 591942 138934
rect 592178 138698 592360 138934
rect 591760 103254 592360 138698
rect 591760 103018 591942 103254
rect 592178 103018 592360 103254
rect 591760 102934 592360 103018
rect 591760 102698 591942 102934
rect 592178 102698 592360 102934
rect 591760 67254 592360 102698
rect 591760 67018 591942 67254
rect 592178 67018 592360 67254
rect 591760 66934 592360 67018
rect 591760 66698 591942 66934
rect 592178 66698 592360 66934
rect 591760 31254 592360 66698
rect 591760 31018 591942 31254
rect 592178 31018 592360 31254
rect 591760 30934 592360 31018
rect 591760 30698 591942 30934
rect 592178 30698 592360 30934
rect 569604 -7022 569786 -6786
rect 570022 -7022 570204 -6786
rect 569604 -7106 570204 -7022
rect 569604 -7342 569786 -7106
rect 570022 -7342 570204 -7106
rect 569604 -7364 570204 -7342
rect 591760 -6786 592360 30698
rect 591760 -7022 591942 -6786
rect 592178 -7022 592360 -6786
rect 591760 -7106 592360 -7022
rect 591760 -7342 591942 -7106
rect 592178 -7342 592360 -7106
rect 591760 -7364 592360 -7342
<< via4 >>
rect -8254 711042 -8018 711278
rect -8254 710722 -8018 710958
rect -8254 679018 -8018 679254
rect -8254 678698 -8018 678934
rect -8254 643018 -8018 643254
rect -8254 642698 -8018 642934
rect -8254 607018 -8018 607254
rect -8254 606698 -8018 606934
rect -8254 571018 -8018 571254
rect -8254 570698 -8018 570934
rect -8254 535018 -8018 535254
rect -8254 534698 -8018 534934
rect -8254 499018 -8018 499254
rect -8254 498698 -8018 498934
rect -8254 463018 -8018 463254
rect -8254 462698 -8018 462934
rect -8254 427018 -8018 427254
rect -8254 426698 -8018 426934
rect -8254 391018 -8018 391254
rect -8254 390698 -8018 390934
rect -8254 355018 -8018 355254
rect -8254 354698 -8018 354934
rect -8254 319018 -8018 319254
rect -8254 318698 -8018 318934
rect -8254 283018 -8018 283254
rect -8254 282698 -8018 282934
rect -8254 247018 -8018 247254
rect -8254 246698 -8018 246934
rect -8254 211018 -8018 211254
rect -8254 210698 -8018 210934
rect -8254 175018 -8018 175254
rect -8254 174698 -8018 174934
rect -8254 139018 -8018 139254
rect -8254 138698 -8018 138934
rect -8254 103018 -8018 103254
rect -8254 102698 -8018 102934
rect -8254 67018 -8018 67254
rect -8254 66698 -8018 66934
rect -8254 31018 -8018 31254
rect -8254 30698 -8018 30934
rect -7334 710122 -7098 710358
rect -7334 709802 -7098 710038
rect 11786 710122 12022 710358
rect 11786 709802 12022 710038
rect -7334 697018 -7098 697254
rect -7334 696698 -7098 696934
rect -7334 661018 -7098 661254
rect -7334 660698 -7098 660934
rect -7334 625018 -7098 625254
rect -7334 624698 -7098 624934
rect -7334 589018 -7098 589254
rect -7334 588698 -7098 588934
rect -7334 553018 -7098 553254
rect -7334 552698 -7098 552934
rect -7334 517018 -7098 517254
rect -7334 516698 -7098 516934
rect -7334 481018 -7098 481254
rect -7334 480698 -7098 480934
rect -7334 445018 -7098 445254
rect -7334 444698 -7098 444934
rect -7334 409018 -7098 409254
rect -7334 408698 -7098 408934
rect -7334 373018 -7098 373254
rect -7334 372698 -7098 372934
rect -7334 337018 -7098 337254
rect -7334 336698 -7098 336934
rect -7334 301018 -7098 301254
rect -7334 300698 -7098 300934
rect -7334 265018 -7098 265254
rect -7334 264698 -7098 264934
rect -7334 229018 -7098 229254
rect -7334 228698 -7098 228934
rect -7334 193018 -7098 193254
rect -7334 192698 -7098 192934
rect -7334 157018 -7098 157254
rect -7334 156698 -7098 156934
rect -7334 121018 -7098 121254
rect -7334 120698 -7098 120934
rect -7334 85018 -7098 85254
rect -7334 84698 -7098 84934
rect -7334 49018 -7098 49254
rect -7334 48698 -7098 48934
rect -7334 13018 -7098 13254
rect -7334 12698 -7098 12934
rect -6414 709202 -6178 709438
rect -6414 708882 -6178 709118
rect -6414 675418 -6178 675654
rect -6414 675098 -6178 675334
rect -6414 639418 -6178 639654
rect -6414 639098 -6178 639334
rect -6414 603418 -6178 603654
rect -6414 603098 -6178 603334
rect -6414 567418 -6178 567654
rect -6414 567098 -6178 567334
rect -6414 531418 -6178 531654
rect -6414 531098 -6178 531334
rect -6414 495418 -6178 495654
rect -6414 495098 -6178 495334
rect -6414 459418 -6178 459654
rect -6414 459098 -6178 459334
rect -6414 423418 -6178 423654
rect -6414 423098 -6178 423334
rect -6414 387418 -6178 387654
rect -6414 387098 -6178 387334
rect -6414 351418 -6178 351654
rect -6414 351098 -6178 351334
rect -6414 315418 -6178 315654
rect -6414 315098 -6178 315334
rect -6414 279418 -6178 279654
rect -6414 279098 -6178 279334
rect -6414 243418 -6178 243654
rect -6414 243098 -6178 243334
rect -6414 207418 -6178 207654
rect -6414 207098 -6178 207334
rect -6414 171418 -6178 171654
rect -6414 171098 -6178 171334
rect -6414 135418 -6178 135654
rect -6414 135098 -6178 135334
rect -6414 99418 -6178 99654
rect -6414 99098 -6178 99334
rect -6414 63418 -6178 63654
rect -6414 63098 -6178 63334
rect -6414 27418 -6178 27654
rect -6414 27098 -6178 27334
rect -5494 708282 -5258 708518
rect -5494 707962 -5258 708198
rect 8186 708282 8422 708518
rect 8186 707962 8422 708198
rect -5494 693418 -5258 693654
rect -5494 693098 -5258 693334
rect -5494 657418 -5258 657654
rect -5494 657098 -5258 657334
rect -5494 621418 -5258 621654
rect -5494 621098 -5258 621334
rect -5494 585418 -5258 585654
rect -5494 585098 -5258 585334
rect -5494 549418 -5258 549654
rect -5494 549098 -5258 549334
rect -5494 513418 -5258 513654
rect -5494 513098 -5258 513334
rect -5494 477418 -5258 477654
rect -5494 477098 -5258 477334
rect -5494 441418 -5258 441654
rect -5494 441098 -5258 441334
rect -5494 405418 -5258 405654
rect -5494 405098 -5258 405334
rect -5494 369418 -5258 369654
rect -5494 369098 -5258 369334
rect -5494 333418 -5258 333654
rect -5494 333098 -5258 333334
rect -5494 297418 -5258 297654
rect -5494 297098 -5258 297334
rect -5494 261418 -5258 261654
rect -5494 261098 -5258 261334
rect -5494 225418 -5258 225654
rect -5494 225098 -5258 225334
rect -5494 189418 -5258 189654
rect -5494 189098 -5258 189334
rect -5494 153418 -5258 153654
rect -5494 153098 -5258 153334
rect -5494 117418 -5258 117654
rect -5494 117098 -5258 117334
rect -5494 81418 -5258 81654
rect -5494 81098 -5258 81334
rect -5494 45418 -5258 45654
rect -5494 45098 -5258 45334
rect -5494 9418 -5258 9654
rect -5494 9098 -5258 9334
rect -4574 707362 -4338 707598
rect -4574 707042 -4338 707278
rect -4574 671818 -4338 672054
rect -4574 671498 -4338 671734
rect -4574 635818 -4338 636054
rect -4574 635498 -4338 635734
rect -4574 599818 -4338 600054
rect -4574 599498 -4338 599734
rect -4574 563818 -4338 564054
rect -4574 563498 -4338 563734
rect -4574 527818 -4338 528054
rect -4574 527498 -4338 527734
rect -4574 491818 -4338 492054
rect -4574 491498 -4338 491734
rect -4574 455818 -4338 456054
rect -4574 455498 -4338 455734
rect -4574 419818 -4338 420054
rect -4574 419498 -4338 419734
rect -4574 383818 -4338 384054
rect -4574 383498 -4338 383734
rect -4574 347818 -4338 348054
rect -4574 347498 -4338 347734
rect -4574 311818 -4338 312054
rect -4574 311498 -4338 311734
rect -4574 275818 -4338 276054
rect -4574 275498 -4338 275734
rect -4574 239818 -4338 240054
rect -4574 239498 -4338 239734
rect -4574 203818 -4338 204054
rect -4574 203498 -4338 203734
rect -4574 167818 -4338 168054
rect -4574 167498 -4338 167734
rect -4574 131818 -4338 132054
rect -4574 131498 -4338 131734
rect -4574 95818 -4338 96054
rect -4574 95498 -4338 95734
rect -4574 59818 -4338 60054
rect -4574 59498 -4338 59734
rect -4574 23818 -4338 24054
rect -4574 23498 -4338 23734
rect -3654 706442 -3418 706678
rect -3654 706122 -3418 706358
rect 4586 706442 4822 706678
rect 4586 706122 4822 706358
rect -3654 689818 -3418 690054
rect -3654 689498 -3418 689734
rect -3654 653818 -3418 654054
rect -3654 653498 -3418 653734
rect -3654 617818 -3418 618054
rect -3654 617498 -3418 617734
rect -3654 581818 -3418 582054
rect -3654 581498 -3418 581734
rect -3654 545818 -3418 546054
rect -3654 545498 -3418 545734
rect -3654 509818 -3418 510054
rect -3654 509498 -3418 509734
rect -3654 473818 -3418 474054
rect -3654 473498 -3418 473734
rect -3654 437818 -3418 438054
rect -3654 437498 -3418 437734
rect -3654 401818 -3418 402054
rect -3654 401498 -3418 401734
rect -3654 365818 -3418 366054
rect -3654 365498 -3418 365734
rect -3654 329818 -3418 330054
rect -3654 329498 -3418 329734
rect -3654 293818 -3418 294054
rect -3654 293498 -3418 293734
rect -3654 257818 -3418 258054
rect -3654 257498 -3418 257734
rect -3654 221818 -3418 222054
rect -3654 221498 -3418 221734
rect -3654 185818 -3418 186054
rect -3654 185498 -3418 185734
rect -3654 149818 -3418 150054
rect -3654 149498 -3418 149734
rect -3654 113818 -3418 114054
rect -3654 113498 -3418 113734
rect -3654 77818 -3418 78054
rect -3654 77498 -3418 77734
rect -3654 41818 -3418 42054
rect -3654 41498 -3418 41734
rect -3654 5818 -3418 6054
rect -3654 5498 -3418 5734
rect -2734 705522 -2498 705758
rect -2734 705202 -2498 705438
rect -2734 668218 -2498 668454
rect -2734 667898 -2498 668134
rect -2734 632218 -2498 632454
rect -2734 631898 -2498 632134
rect -2734 596218 -2498 596454
rect -2734 595898 -2498 596134
rect -2734 560218 -2498 560454
rect -2734 559898 -2498 560134
rect -2734 524218 -2498 524454
rect -2734 523898 -2498 524134
rect -2734 488218 -2498 488454
rect -2734 487898 -2498 488134
rect -2734 452218 -2498 452454
rect -2734 451898 -2498 452134
rect -2734 416218 -2498 416454
rect -2734 415898 -2498 416134
rect -2734 380218 -2498 380454
rect -2734 379898 -2498 380134
rect -2734 344218 -2498 344454
rect -2734 343898 -2498 344134
rect -2734 308218 -2498 308454
rect -2734 307898 -2498 308134
rect -2734 272218 -2498 272454
rect -2734 271898 -2498 272134
rect -2734 236218 -2498 236454
rect -2734 235898 -2498 236134
rect -2734 200218 -2498 200454
rect -2734 199898 -2498 200134
rect -2734 164218 -2498 164454
rect -2734 163898 -2498 164134
rect -2734 128218 -2498 128454
rect -2734 127898 -2498 128134
rect -2734 92218 -2498 92454
rect -2734 91898 -2498 92134
rect -2734 56218 -2498 56454
rect -2734 55898 -2498 56134
rect -2734 20218 -2498 20454
rect -2734 19898 -2498 20134
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 686218 -1578 686454
rect -1814 685898 -1578 686134
rect -1814 650218 -1578 650454
rect -1814 649898 -1578 650134
rect -1814 614218 -1578 614454
rect -1814 613898 -1578 614134
rect -1814 578218 -1578 578454
rect -1814 577898 -1578 578134
rect -1814 542218 -1578 542454
rect -1814 541898 -1578 542134
rect -1814 506218 -1578 506454
rect -1814 505898 -1578 506134
rect -1814 470218 -1578 470454
rect -1814 469898 -1578 470134
rect -1814 434218 -1578 434454
rect -1814 433898 -1578 434134
rect -1814 398218 -1578 398454
rect -1814 397898 -1578 398134
rect -1814 362218 -1578 362454
rect -1814 361898 -1578 362134
rect -1814 326218 -1578 326454
rect -1814 325898 -1578 326134
rect -1814 290218 -1578 290454
rect -1814 289898 -1578 290134
rect -1814 254218 -1578 254454
rect -1814 253898 -1578 254134
rect -1814 218218 -1578 218454
rect -1814 217898 -1578 218134
rect -1814 182218 -1578 182454
rect -1814 181898 -1578 182134
rect -1814 146218 -1578 146454
rect -1814 145898 -1578 146134
rect -1814 110218 -1578 110454
rect -1814 109898 -1578 110134
rect -1814 74218 -1578 74454
rect -1814 73898 -1578 74134
rect -1814 38218 -1578 38454
rect -1814 37898 -1578 38134
rect -1814 2218 -1578 2454
rect -1814 1898 -1578 2134
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 986 704602 1222 704838
rect 986 704282 1222 704518
rect 986 686218 1222 686454
rect 986 685898 1222 686134
rect 986 650218 1222 650454
rect 986 649898 1222 650134
rect 986 614218 1222 614454
rect 986 613898 1222 614134
rect 986 578218 1222 578454
rect 986 577898 1222 578134
rect 986 542218 1222 542454
rect 986 541898 1222 542134
rect 986 506218 1222 506454
rect 986 505898 1222 506134
rect 986 470218 1222 470454
rect 986 469898 1222 470134
rect 986 434218 1222 434454
rect 986 433898 1222 434134
rect 986 398218 1222 398454
rect 986 397898 1222 398134
rect 986 362218 1222 362454
rect 986 361898 1222 362134
rect 986 326218 1222 326454
rect 986 325898 1222 326134
rect 986 290218 1222 290454
rect 986 289898 1222 290134
rect 986 254218 1222 254454
rect 986 253898 1222 254134
rect 986 218218 1222 218454
rect 986 217898 1222 218134
rect 986 182218 1222 182454
rect 986 181898 1222 182134
rect 986 146218 1222 146454
rect 986 145898 1222 146134
rect 986 110218 1222 110454
rect 986 109898 1222 110134
rect 986 74218 1222 74454
rect 986 73898 1222 74134
rect 986 38218 1222 38454
rect 986 37898 1222 38134
rect 986 2218 1222 2454
rect 986 1898 1222 2134
rect 986 -582 1222 -346
rect 986 -902 1222 -666
rect -2734 -1502 -2498 -1266
rect -2734 -1822 -2498 -1586
rect 4586 689818 4822 690054
rect 4586 689498 4822 689734
rect 4586 653818 4822 654054
rect 4586 653498 4822 653734
rect 4586 617818 4822 618054
rect 4586 617498 4822 617734
rect 4586 581818 4822 582054
rect 4586 581498 4822 581734
rect 8186 693418 8422 693654
rect 8186 693098 8422 693334
rect 8186 657418 8422 657654
rect 8186 657098 8422 657334
rect 8186 621418 8422 621654
rect 8186 621098 8422 621334
rect 8186 585418 8422 585654
rect 8186 585098 8422 585334
rect 5126 562732 5362 562818
rect 5126 562668 5212 562732
rect 5212 562668 5276 562732
rect 5276 562668 5362 562732
rect 5126 562582 5362 562668
rect 4586 545818 4822 546054
rect 4586 545498 4822 545734
rect 4586 509818 4822 510054
rect 4586 509498 4822 509734
rect 4586 473818 4822 474054
rect 4586 473498 4822 473734
rect 4586 437818 4822 438054
rect 4586 437498 4822 437734
rect 4586 401818 4822 402054
rect 4586 401498 4822 401734
rect 4586 365818 4822 366054
rect 4586 365498 4822 365734
rect 4586 329818 4822 330054
rect 4586 329498 4822 329734
rect 4586 293818 4822 294054
rect 4586 293498 4822 293734
rect 4586 257818 4822 258054
rect 4586 257498 4822 257734
rect 4586 221818 4822 222054
rect 4586 221498 4822 221734
rect 4586 185818 4822 186054
rect 4586 185498 4822 185734
rect 4586 149818 4822 150054
rect 4586 149498 4822 149734
rect 4586 113818 4822 114054
rect 4586 113498 4822 113734
rect 4586 77818 4822 78054
rect 4586 77498 4822 77734
rect 4586 41818 4822 42054
rect 4586 41498 4822 41734
rect 4586 5818 4822 6054
rect 4586 5498 4822 5734
rect -3654 -2422 -3418 -2186
rect -3654 -2742 -3418 -2506
rect 4586 -2422 4822 -2186
rect 4586 -2742 4822 -2506
rect -4574 -3342 -4338 -3106
rect -4574 -3662 -4338 -3426
rect 8186 549418 8422 549654
rect 8186 549098 8422 549334
rect 8186 513418 8422 513654
rect 8186 513098 8422 513334
rect 8186 477418 8422 477654
rect 8186 477098 8422 477334
rect 8186 441418 8422 441654
rect 8186 441098 8422 441334
rect 8186 405418 8422 405654
rect 8186 405098 8422 405334
rect 8186 369418 8422 369654
rect 8186 369098 8422 369334
rect 8186 333418 8422 333654
rect 8186 333098 8422 333334
rect 8186 297418 8422 297654
rect 8186 297098 8422 297334
rect 8186 261418 8422 261654
rect 8186 261098 8422 261334
rect 8186 225418 8422 225654
rect 8186 225098 8422 225334
rect 8186 189418 8422 189654
rect 8186 189098 8422 189334
rect 8186 153418 8422 153654
rect 8186 153098 8422 153334
rect 8186 117418 8422 117654
rect 8186 117098 8422 117334
rect 8186 81418 8422 81654
rect 8186 81098 8422 81334
rect 8186 45418 8422 45654
rect 8186 45098 8422 45334
rect 8186 9418 8422 9654
rect 8186 9098 8422 9334
rect -5494 -4262 -5258 -4026
rect -5494 -4582 -5258 -4346
rect 8186 -4262 8422 -4026
rect 8186 -4582 8422 -4346
rect -6414 -5182 -6178 -4946
rect -6414 -5502 -6178 -5266
rect 29786 711042 30022 711278
rect 29786 710722 30022 710958
rect 26186 709202 26422 709438
rect 26186 708882 26422 709118
rect 22586 707362 22822 707598
rect 22586 707042 22822 707278
rect 11786 697018 12022 697254
rect 11786 696698 12022 696934
rect 11786 661018 12022 661254
rect 11786 660698 12022 660934
rect 11786 625018 12022 625254
rect 11786 624698 12022 624934
rect 11786 589018 12022 589254
rect 11786 588698 12022 588934
rect 11786 553018 12022 553254
rect 11786 552698 12022 552934
rect 11786 517018 12022 517254
rect 11786 516698 12022 516934
rect 11786 481018 12022 481254
rect 11786 480698 12022 480934
rect 11786 445018 12022 445254
rect 11786 444698 12022 444934
rect 11786 409018 12022 409254
rect 11786 408698 12022 408934
rect 11786 373018 12022 373254
rect 11786 372698 12022 372934
rect 11786 337018 12022 337254
rect 11786 336698 12022 336934
rect 11786 301018 12022 301254
rect 11786 300698 12022 300934
rect 11786 265018 12022 265254
rect 11786 264698 12022 264934
rect 11786 229018 12022 229254
rect 11786 228698 12022 228934
rect 11786 193018 12022 193254
rect 11786 192698 12022 192934
rect 11786 157018 12022 157254
rect 11786 156698 12022 156934
rect 11786 121018 12022 121254
rect 11786 120698 12022 120934
rect 11786 85018 12022 85254
rect 11786 84698 12022 84934
rect 11786 49018 12022 49254
rect 11786 48698 12022 48934
rect 11786 13018 12022 13254
rect 11786 12698 12022 12934
rect -7334 -6102 -7098 -5866
rect -7334 -6422 -7098 -6186
rect 18986 705522 19222 705758
rect 18986 705202 19222 705438
rect 18986 668218 19222 668454
rect 18986 667898 19222 668134
rect 18986 632218 19222 632454
rect 18986 631898 19222 632134
rect 18986 596218 19222 596454
rect 18986 595898 19222 596134
rect 18986 560218 19222 560454
rect 18986 559898 19222 560134
rect 18986 524218 19222 524454
rect 18986 523898 19222 524134
rect 18986 488218 19222 488454
rect 18986 487898 19222 488134
rect 18986 452218 19222 452454
rect 18986 451898 19222 452134
rect 18986 416218 19222 416454
rect 18986 415898 19222 416134
rect 18986 380218 19222 380454
rect 18986 379898 19222 380134
rect 18986 344218 19222 344454
rect 18986 343898 19222 344134
rect 18986 308218 19222 308454
rect 18986 307898 19222 308134
rect 18986 272218 19222 272454
rect 18986 271898 19222 272134
rect 18986 236218 19222 236454
rect 18986 235898 19222 236134
rect 18986 200218 19222 200454
rect 18986 199898 19222 200134
rect 18986 164218 19222 164454
rect 18986 163898 19222 164134
rect 18986 128218 19222 128454
rect 18986 127898 19222 128134
rect 18986 92218 19222 92454
rect 18986 91898 19222 92134
rect 18986 56218 19222 56454
rect 18986 55898 19222 56134
rect 18986 20218 19222 20454
rect 18986 19898 19222 20134
rect 18986 -1502 19222 -1266
rect 18986 -1822 19222 -1586
rect 22586 671818 22822 672054
rect 22586 671498 22822 671734
rect 22586 635818 22822 636054
rect 22586 635498 22822 635734
rect 22586 599818 22822 600054
rect 22586 599498 22822 599734
rect 22586 563818 22822 564054
rect 22586 563498 22822 563734
rect 22586 527818 22822 528054
rect 22586 527498 22822 527734
rect 22586 491818 22822 492054
rect 22586 491498 22822 491734
rect 22586 455818 22822 456054
rect 22586 455498 22822 455734
rect 22586 419818 22822 420054
rect 22586 419498 22822 419734
rect 22586 383818 22822 384054
rect 22586 383498 22822 383734
rect 22586 347818 22822 348054
rect 22586 347498 22822 347734
rect 22586 311818 22822 312054
rect 22586 311498 22822 311734
rect 22586 275818 22822 276054
rect 22586 275498 22822 275734
rect 22586 239818 22822 240054
rect 22586 239498 22822 239734
rect 22586 203818 22822 204054
rect 22586 203498 22822 203734
rect 22586 167818 22822 168054
rect 22586 167498 22822 167734
rect 22586 131818 22822 132054
rect 22586 131498 22822 131734
rect 22586 95818 22822 96054
rect 22586 95498 22822 95734
rect 22586 59818 22822 60054
rect 22586 59498 22822 59734
rect 22586 23818 22822 24054
rect 22586 23498 22822 23734
rect 22586 -3342 22822 -3106
rect 22586 -3662 22822 -3426
rect 26186 675418 26422 675654
rect 26186 675098 26422 675334
rect 26186 639418 26422 639654
rect 26186 639098 26422 639334
rect 26186 603418 26422 603654
rect 26186 603098 26422 603334
rect 26186 567418 26422 567654
rect 26186 567098 26422 567334
rect 26186 531418 26422 531654
rect 26186 531098 26422 531334
rect 26186 495418 26422 495654
rect 26186 495098 26422 495334
rect 26186 459418 26422 459654
rect 26186 459098 26422 459334
rect 26186 423418 26422 423654
rect 26186 423098 26422 423334
rect 26186 387418 26422 387654
rect 26186 387098 26422 387334
rect 26186 351418 26422 351654
rect 26186 351098 26422 351334
rect 26186 315418 26422 315654
rect 26186 315098 26422 315334
rect 26186 279418 26422 279654
rect 26186 279098 26422 279334
rect 26186 243418 26422 243654
rect 26186 243098 26422 243334
rect 26186 207418 26422 207654
rect 26186 207098 26422 207334
rect 26186 171418 26422 171654
rect 26186 171098 26422 171334
rect 26186 135418 26422 135654
rect 26186 135098 26422 135334
rect 26186 99418 26422 99654
rect 26186 99098 26422 99334
rect 26186 63418 26422 63654
rect 26186 63098 26422 63334
rect 26186 27418 26422 27654
rect 26186 27098 26422 27334
rect 26186 -5182 26422 -4946
rect 26186 -5502 26422 -5266
rect 47786 710122 48022 710358
rect 47786 709802 48022 710038
rect 44186 708282 44422 708518
rect 44186 707962 44422 708198
rect 40586 706442 40822 706678
rect 40586 706122 40822 706358
rect 29786 679018 30022 679254
rect 29786 678698 30022 678934
rect 29786 643018 30022 643254
rect 29786 642698 30022 642934
rect 29786 607018 30022 607254
rect 29786 606698 30022 606934
rect 29786 571018 30022 571254
rect 29786 570698 30022 570934
rect 29786 535018 30022 535254
rect 29786 534698 30022 534934
rect 29786 499018 30022 499254
rect 29786 498698 30022 498934
rect 29786 463018 30022 463254
rect 29786 462698 30022 462934
rect 29786 427018 30022 427254
rect 29786 426698 30022 426934
rect 29786 391018 30022 391254
rect 29786 390698 30022 390934
rect 29786 355018 30022 355254
rect 29786 354698 30022 354934
rect 29786 319018 30022 319254
rect 29786 318698 30022 318934
rect 29786 283018 30022 283254
rect 29786 282698 30022 282934
rect 29786 247018 30022 247254
rect 29786 246698 30022 246934
rect 29786 211018 30022 211254
rect 29786 210698 30022 210934
rect 29786 175018 30022 175254
rect 29786 174698 30022 174934
rect 29786 139018 30022 139254
rect 29786 138698 30022 138934
rect 29786 103018 30022 103254
rect 29786 102698 30022 102934
rect 29786 67018 30022 67254
rect 29786 66698 30022 66934
rect 29786 31018 30022 31254
rect 29786 30698 30022 30934
rect 11786 -6102 12022 -5866
rect 11786 -6422 12022 -6186
rect -8254 -7022 -8018 -6786
rect -8254 -7342 -8018 -7106
rect 36986 704602 37222 704838
rect 36986 704282 37222 704518
rect 36986 686218 37222 686454
rect 36986 685898 37222 686134
rect 36986 650218 37222 650454
rect 36986 649898 37222 650134
rect 36986 614218 37222 614454
rect 36986 613898 37222 614134
rect 36986 578218 37222 578454
rect 36986 577898 37222 578134
rect 36986 542218 37222 542454
rect 36986 541898 37222 542134
rect 36986 506218 37222 506454
rect 36986 505898 37222 506134
rect 36986 470218 37222 470454
rect 36986 469898 37222 470134
rect 36986 434218 37222 434454
rect 36986 433898 37222 434134
rect 36986 398218 37222 398454
rect 36986 397898 37222 398134
rect 36986 362218 37222 362454
rect 36986 361898 37222 362134
rect 36986 326218 37222 326454
rect 36986 325898 37222 326134
rect 36986 290218 37222 290454
rect 36986 289898 37222 290134
rect 36986 254218 37222 254454
rect 36986 253898 37222 254134
rect 36986 218218 37222 218454
rect 36986 217898 37222 218134
rect 36986 182218 37222 182454
rect 36986 181898 37222 182134
rect 36986 146218 37222 146454
rect 36986 145898 37222 146134
rect 36986 110218 37222 110454
rect 36986 109898 37222 110134
rect 36986 74218 37222 74454
rect 36986 73898 37222 74134
rect 36986 38218 37222 38454
rect 36986 37898 37222 38134
rect 36986 2218 37222 2454
rect 36986 1898 37222 2134
rect 36986 -582 37222 -346
rect 36986 -902 37222 -666
rect 40586 689818 40822 690054
rect 40586 689498 40822 689734
rect 40586 653818 40822 654054
rect 40586 653498 40822 653734
rect 40586 617818 40822 618054
rect 40586 617498 40822 617734
rect 40586 581818 40822 582054
rect 40586 581498 40822 581734
rect 40586 545818 40822 546054
rect 40586 545498 40822 545734
rect 40586 509818 40822 510054
rect 40586 509498 40822 509734
rect 40586 473818 40822 474054
rect 40586 473498 40822 473734
rect 40586 437818 40822 438054
rect 40586 437498 40822 437734
rect 40586 401818 40822 402054
rect 40586 401498 40822 401734
rect 40586 365818 40822 366054
rect 40586 365498 40822 365734
rect 40586 329818 40822 330054
rect 40586 329498 40822 329734
rect 40586 293818 40822 294054
rect 40586 293498 40822 293734
rect 40586 257818 40822 258054
rect 40586 257498 40822 257734
rect 40586 221818 40822 222054
rect 40586 221498 40822 221734
rect 40586 185818 40822 186054
rect 40586 185498 40822 185734
rect 40586 149818 40822 150054
rect 40586 149498 40822 149734
rect 40586 113818 40822 114054
rect 40586 113498 40822 113734
rect 40586 77818 40822 78054
rect 40586 77498 40822 77734
rect 40586 41818 40822 42054
rect 40586 41498 40822 41734
rect 40586 5818 40822 6054
rect 40586 5498 40822 5734
rect 40586 -2422 40822 -2186
rect 40586 -2742 40822 -2506
rect 44186 693418 44422 693654
rect 44186 693098 44422 693334
rect 44186 657418 44422 657654
rect 44186 657098 44422 657334
rect 44186 621418 44422 621654
rect 44186 621098 44422 621334
rect 44186 585418 44422 585654
rect 44186 585098 44422 585334
rect 44186 549418 44422 549654
rect 44186 549098 44422 549334
rect 44186 513418 44422 513654
rect 44186 513098 44422 513334
rect 44186 477418 44422 477654
rect 44186 477098 44422 477334
rect 44186 441418 44422 441654
rect 44186 441098 44422 441334
rect 44186 405418 44422 405654
rect 44186 405098 44422 405334
rect 44186 369418 44422 369654
rect 44186 369098 44422 369334
rect 44186 333418 44422 333654
rect 44186 333098 44422 333334
rect 44186 297418 44422 297654
rect 44186 297098 44422 297334
rect 44186 261418 44422 261654
rect 44186 261098 44422 261334
rect 44186 225418 44422 225654
rect 44186 225098 44422 225334
rect 44186 189418 44422 189654
rect 44186 189098 44422 189334
rect 44186 153418 44422 153654
rect 44186 153098 44422 153334
rect 44186 117418 44422 117654
rect 44186 117098 44422 117334
rect 44186 81418 44422 81654
rect 44186 81098 44422 81334
rect 44186 45418 44422 45654
rect 44186 45098 44422 45334
rect 44186 9418 44422 9654
rect 44186 9098 44422 9334
rect 44186 -4262 44422 -4026
rect 44186 -4582 44422 -4346
rect 65786 711042 66022 711278
rect 65786 710722 66022 710958
rect 62186 709202 62422 709438
rect 62186 708882 62422 709118
rect 58586 707362 58822 707598
rect 58586 707042 58822 707278
rect 47786 697018 48022 697254
rect 47786 696698 48022 696934
rect 47786 661018 48022 661254
rect 47786 660698 48022 660934
rect 47786 625018 48022 625254
rect 47786 624698 48022 624934
rect 47786 589018 48022 589254
rect 47786 588698 48022 588934
rect 54986 705522 55222 705758
rect 54986 705202 55222 705438
rect 54986 668218 55222 668454
rect 54986 667898 55222 668134
rect 54986 632218 55222 632454
rect 54986 631898 55222 632134
rect 54986 596218 55222 596454
rect 54986 595898 55222 596134
rect 50390 561372 50626 561458
rect 50390 561308 50476 561372
rect 50476 561308 50540 561372
rect 50540 561308 50626 561372
rect 50390 561222 50626 561308
rect 51494 561372 51730 561458
rect 51494 561308 51580 561372
rect 51580 561308 51644 561372
rect 51644 561308 51730 561372
rect 51494 561222 51730 561308
rect 47786 553018 48022 553254
rect 47786 552698 48022 552934
rect 47786 517018 48022 517254
rect 47786 516698 48022 516934
rect 47786 481018 48022 481254
rect 47786 480698 48022 480934
rect 47786 445018 48022 445254
rect 47786 444698 48022 444934
rect 47786 409018 48022 409254
rect 47786 408698 48022 408934
rect 47786 373018 48022 373254
rect 47786 372698 48022 372934
rect 47786 337018 48022 337254
rect 47786 336698 48022 336934
rect 47786 301018 48022 301254
rect 47786 300698 48022 300934
rect 47786 265018 48022 265254
rect 47786 264698 48022 264934
rect 47786 229018 48022 229254
rect 47786 228698 48022 228934
rect 47786 193018 48022 193254
rect 47786 192698 48022 192934
rect 47786 157018 48022 157254
rect 47786 156698 48022 156934
rect 47786 121018 48022 121254
rect 47786 120698 48022 120934
rect 47786 85018 48022 85254
rect 47786 84698 48022 84934
rect 47786 49018 48022 49254
rect 47786 48698 48022 48934
rect 47786 13018 48022 13254
rect 47786 12698 48022 12934
rect 29786 -7022 30022 -6786
rect 29786 -7342 30022 -7106
rect 54986 560218 55222 560454
rect 54986 559898 55222 560134
rect 54986 524218 55222 524454
rect 54986 523898 55222 524134
rect 54986 488218 55222 488454
rect 54986 487898 55222 488134
rect 54986 452218 55222 452454
rect 54986 451898 55222 452134
rect 54986 416218 55222 416454
rect 54986 415898 55222 416134
rect 54986 380218 55222 380454
rect 54986 379898 55222 380134
rect 54986 344218 55222 344454
rect 54986 343898 55222 344134
rect 54986 308218 55222 308454
rect 54986 307898 55222 308134
rect 54986 272218 55222 272454
rect 54986 271898 55222 272134
rect 54986 236218 55222 236454
rect 54986 235898 55222 236134
rect 54986 200218 55222 200454
rect 54986 199898 55222 200134
rect 54986 164218 55222 164454
rect 54986 163898 55222 164134
rect 54986 128218 55222 128454
rect 54986 127898 55222 128134
rect 54986 92218 55222 92454
rect 54986 91898 55222 92134
rect 54986 56218 55222 56454
rect 54986 55898 55222 56134
rect 54986 20218 55222 20454
rect 54986 19898 55222 20134
rect 54986 -1502 55222 -1266
rect 54986 -1822 55222 -1586
rect 58586 671818 58822 672054
rect 58586 671498 58822 671734
rect 58586 635818 58822 636054
rect 58586 635498 58822 635734
rect 58586 599818 58822 600054
rect 58586 599498 58822 599734
rect 58586 563818 58822 564054
rect 58586 563498 58822 563734
rect 58586 527818 58822 528054
rect 58586 527498 58822 527734
rect 58586 491818 58822 492054
rect 58586 491498 58822 491734
rect 58586 455818 58822 456054
rect 58586 455498 58822 455734
rect 58586 419818 58822 420054
rect 58586 419498 58822 419734
rect 58586 383818 58822 384054
rect 58586 383498 58822 383734
rect 58586 347818 58822 348054
rect 58586 347498 58822 347734
rect 58586 311818 58822 312054
rect 58586 311498 58822 311734
rect 58586 275818 58822 276054
rect 58586 275498 58822 275734
rect 58586 239818 58822 240054
rect 58586 239498 58822 239734
rect 58586 203818 58822 204054
rect 58586 203498 58822 203734
rect 58586 167818 58822 168054
rect 58586 167498 58822 167734
rect 58586 131818 58822 132054
rect 58586 131498 58822 131734
rect 58586 95818 58822 96054
rect 58586 95498 58822 95734
rect 58586 59818 58822 60054
rect 58586 59498 58822 59734
rect 58586 23818 58822 24054
rect 58586 23498 58822 23734
rect 58586 -3342 58822 -3106
rect 58586 -3662 58822 -3426
rect 62186 675418 62422 675654
rect 62186 675098 62422 675334
rect 62186 639418 62422 639654
rect 62186 639098 62422 639334
rect 62186 603418 62422 603654
rect 62186 603098 62422 603334
rect 62186 567418 62422 567654
rect 62186 567098 62422 567334
rect 62186 531418 62422 531654
rect 62186 531098 62422 531334
rect 62186 495418 62422 495654
rect 62186 495098 62422 495334
rect 62186 459418 62422 459654
rect 62186 459098 62422 459334
rect 62186 423418 62422 423654
rect 62186 423098 62422 423334
rect 62186 387418 62422 387654
rect 62186 387098 62422 387334
rect 62186 351418 62422 351654
rect 62186 351098 62422 351334
rect 62186 315418 62422 315654
rect 62186 315098 62422 315334
rect 62186 279418 62422 279654
rect 62186 279098 62422 279334
rect 62186 243418 62422 243654
rect 62186 243098 62422 243334
rect 62186 207418 62422 207654
rect 62186 207098 62422 207334
rect 62186 171418 62422 171654
rect 62186 171098 62422 171334
rect 62186 135418 62422 135654
rect 62186 135098 62422 135334
rect 62186 99418 62422 99654
rect 62186 99098 62422 99334
rect 62186 63418 62422 63654
rect 62186 63098 62422 63334
rect 62186 27418 62422 27654
rect 62186 27098 62422 27334
rect 62186 -5182 62422 -4946
rect 62186 -5502 62422 -5266
rect 83786 710122 84022 710358
rect 83786 709802 84022 710038
rect 80186 708282 80422 708518
rect 80186 707962 80422 708198
rect 76586 706442 76822 706678
rect 76586 706122 76822 706358
rect 65786 679018 66022 679254
rect 65786 678698 66022 678934
rect 65786 643018 66022 643254
rect 65786 642698 66022 642934
rect 65786 607018 66022 607254
rect 65786 606698 66022 606934
rect 65786 571018 66022 571254
rect 65786 570698 66022 570934
rect 65786 535018 66022 535254
rect 65786 534698 66022 534934
rect 65786 499018 66022 499254
rect 65786 498698 66022 498934
rect 65786 463018 66022 463254
rect 65786 462698 66022 462934
rect 65786 427018 66022 427254
rect 65786 426698 66022 426934
rect 65786 391018 66022 391254
rect 65786 390698 66022 390934
rect 65786 355018 66022 355254
rect 65786 354698 66022 354934
rect 65786 319018 66022 319254
rect 65786 318698 66022 318934
rect 65786 283018 66022 283254
rect 65786 282698 66022 282934
rect 65786 247018 66022 247254
rect 65786 246698 66022 246934
rect 65786 211018 66022 211254
rect 65786 210698 66022 210934
rect 65786 175018 66022 175254
rect 65786 174698 66022 174934
rect 65786 139018 66022 139254
rect 65786 138698 66022 138934
rect 65786 103018 66022 103254
rect 65786 102698 66022 102934
rect 65786 67018 66022 67254
rect 65786 66698 66022 66934
rect 65786 31018 66022 31254
rect 65786 30698 66022 30934
rect 47786 -6102 48022 -5866
rect 47786 -6422 48022 -6186
rect 72986 704602 73222 704838
rect 72986 704282 73222 704518
rect 72986 686218 73222 686454
rect 72986 685898 73222 686134
rect 72986 650218 73222 650454
rect 72986 649898 73222 650134
rect 72986 614218 73222 614454
rect 72986 613898 73222 614134
rect 72986 578218 73222 578454
rect 72986 577898 73222 578134
rect 72986 542218 73222 542454
rect 72986 541898 73222 542134
rect 72986 506218 73222 506454
rect 72986 505898 73222 506134
rect 72986 470218 73222 470454
rect 72986 469898 73222 470134
rect 72986 434218 73222 434454
rect 72986 433898 73222 434134
rect 72986 398218 73222 398454
rect 72986 397898 73222 398134
rect 72986 362218 73222 362454
rect 72986 361898 73222 362134
rect 72986 326218 73222 326454
rect 72986 325898 73222 326134
rect 72986 290218 73222 290454
rect 72986 289898 73222 290134
rect 72986 254218 73222 254454
rect 72986 253898 73222 254134
rect 72986 218218 73222 218454
rect 72986 217898 73222 218134
rect 72986 182218 73222 182454
rect 72986 181898 73222 182134
rect 72986 146218 73222 146454
rect 72986 145898 73222 146134
rect 72986 110218 73222 110454
rect 72986 109898 73222 110134
rect 72986 74218 73222 74454
rect 72986 73898 73222 74134
rect 72986 38218 73222 38454
rect 72986 37898 73222 38134
rect 72986 2218 73222 2454
rect 72986 1898 73222 2134
rect 72986 -582 73222 -346
rect 72986 -902 73222 -666
rect 76586 689818 76822 690054
rect 76586 689498 76822 689734
rect 76586 653818 76822 654054
rect 76586 653498 76822 653734
rect 76586 617818 76822 618054
rect 76586 617498 76822 617734
rect 76586 581818 76822 582054
rect 76586 581498 76822 581734
rect 76586 545818 76822 546054
rect 76586 545498 76822 545734
rect 76586 509818 76822 510054
rect 76586 509498 76822 509734
rect 76586 473818 76822 474054
rect 76586 473498 76822 473734
rect 76586 437818 76822 438054
rect 76586 437498 76822 437734
rect 76586 401818 76822 402054
rect 76586 401498 76822 401734
rect 76586 365818 76822 366054
rect 76586 365498 76822 365734
rect 76586 329818 76822 330054
rect 76586 329498 76822 329734
rect 76586 293818 76822 294054
rect 76586 293498 76822 293734
rect 76586 257818 76822 258054
rect 76586 257498 76822 257734
rect 76586 221818 76822 222054
rect 76586 221498 76822 221734
rect 76586 185818 76822 186054
rect 76586 185498 76822 185734
rect 76586 149818 76822 150054
rect 76586 149498 76822 149734
rect 76586 113818 76822 114054
rect 76586 113498 76822 113734
rect 76586 77818 76822 78054
rect 76586 77498 76822 77734
rect 76586 41818 76822 42054
rect 76586 41498 76822 41734
rect 76586 5818 76822 6054
rect 76586 5498 76822 5734
rect 76586 -2422 76822 -2186
rect 76586 -2742 76822 -2506
rect 80186 693418 80422 693654
rect 80186 693098 80422 693334
rect 80186 657418 80422 657654
rect 80186 657098 80422 657334
rect 80186 621418 80422 621654
rect 80186 621098 80422 621334
rect 80186 585418 80422 585654
rect 80186 585098 80422 585334
rect 80186 549418 80422 549654
rect 80186 549098 80422 549334
rect 80186 513418 80422 513654
rect 80186 513098 80422 513334
rect 80186 477418 80422 477654
rect 80186 477098 80422 477334
rect 80186 441418 80422 441654
rect 80186 441098 80422 441334
rect 80186 405418 80422 405654
rect 80186 405098 80422 405334
rect 80186 369418 80422 369654
rect 80186 369098 80422 369334
rect 80186 333418 80422 333654
rect 80186 333098 80422 333334
rect 80186 297418 80422 297654
rect 80186 297098 80422 297334
rect 80186 261418 80422 261654
rect 80186 261098 80422 261334
rect 80186 225418 80422 225654
rect 80186 225098 80422 225334
rect 80186 189418 80422 189654
rect 80186 189098 80422 189334
rect 80186 153418 80422 153654
rect 80186 153098 80422 153334
rect 80186 117418 80422 117654
rect 80186 117098 80422 117334
rect 80186 81418 80422 81654
rect 80186 81098 80422 81334
rect 80186 45418 80422 45654
rect 80186 45098 80422 45334
rect 80186 9418 80422 9654
rect 80186 9098 80422 9334
rect 80186 -4262 80422 -4026
rect 80186 -4582 80422 -4346
rect 101786 711042 102022 711278
rect 101786 710722 102022 710958
rect 98186 709202 98422 709438
rect 98186 708882 98422 709118
rect 94586 707362 94822 707598
rect 94586 707042 94822 707278
rect 83786 697018 84022 697254
rect 83786 696698 84022 696934
rect 83786 661018 84022 661254
rect 83786 660698 84022 660934
rect 83786 625018 84022 625254
rect 83786 624698 84022 624934
rect 83786 589018 84022 589254
rect 83786 588698 84022 588934
rect 90986 705522 91222 705758
rect 90986 705202 91222 705438
rect 90986 668218 91222 668454
rect 90986 667898 91222 668134
rect 90986 632218 91222 632454
rect 90986 631898 91222 632134
rect 90986 596218 91222 596454
rect 90986 595898 91222 596134
rect 85534 561372 85770 561458
rect 85534 561308 85620 561372
rect 85620 561308 85684 561372
rect 85684 561308 85770 561372
rect 85534 561222 85770 561308
rect 90134 561372 90370 561458
rect 90134 561308 90220 561372
rect 90220 561308 90284 561372
rect 90284 561308 90370 561372
rect 90134 561222 90370 561308
rect 83786 553018 84022 553254
rect 83786 552698 84022 552934
rect 83786 517018 84022 517254
rect 83786 516698 84022 516934
rect 83786 481018 84022 481254
rect 83786 480698 84022 480934
rect 83786 445018 84022 445254
rect 83786 444698 84022 444934
rect 83786 409018 84022 409254
rect 83786 408698 84022 408934
rect 83786 373018 84022 373254
rect 83786 372698 84022 372934
rect 83786 337018 84022 337254
rect 83786 336698 84022 336934
rect 83786 301018 84022 301254
rect 83786 300698 84022 300934
rect 83786 265018 84022 265254
rect 83786 264698 84022 264934
rect 83786 229018 84022 229254
rect 83786 228698 84022 228934
rect 83786 193018 84022 193254
rect 83786 192698 84022 192934
rect 83786 157018 84022 157254
rect 83786 156698 84022 156934
rect 83786 121018 84022 121254
rect 83786 120698 84022 120934
rect 83786 85018 84022 85254
rect 83786 84698 84022 84934
rect 83786 49018 84022 49254
rect 83786 48698 84022 48934
rect 83786 13018 84022 13254
rect 83786 12698 84022 12934
rect 65786 -7022 66022 -6786
rect 65786 -7342 66022 -7106
rect 90986 560218 91222 560454
rect 90986 559898 91222 560134
rect 90986 524218 91222 524454
rect 90986 523898 91222 524134
rect 90986 488218 91222 488454
rect 90986 487898 91222 488134
rect 90986 452218 91222 452454
rect 90986 451898 91222 452134
rect 90986 416218 91222 416454
rect 90986 415898 91222 416134
rect 90986 380218 91222 380454
rect 90986 379898 91222 380134
rect 90986 344218 91222 344454
rect 90986 343898 91222 344134
rect 90986 308218 91222 308454
rect 90986 307898 91222 308134
rect 90986 272218 91222 272454
rect 90986 271898 91222 272134
rect 90986 236218 91222 236454
rect 90986 235898 91222 236134
rect 90986 200218 91222 200454
rect 90986 199898 91222 200134
rect 90986 164218 91222 164454
rect 90986 163898 91222 164134
rect 90986 128218 91222 128454
rect 90986 127898 91222 128134
rect 90986 92218 91222 92454
rect 90986 91898 91222 92134
rect 90986 56218 91222 56454
rect 90986 55898 91222 56134
rect 90986 20218 91222 20454
rect 90986 19898 91222 20134
rect 90986 -1502 91222 -1266
rect 90986 -1822 91222 -1586
rect 94586 671818 94822 672054
rect 94586 671498 94822 671734
rect 94586 635818 94822 636054
rect 94586 635498 94822 635734
rect 94586 599818 94822 600054
rect 94586 599498 94822 599734
rect 94586 563818 94822 564054
rect 94586 563498 94822 563734
rect 94586 527818 94822 528054
rect 94586 527498 94822 527734
rect 94586 491818 94822 492054
rect 94586 491498 94822 491734
rect 94586 455818 94822 456054
rect 94586 455498 94822 455734
rect 94586 419818 94822 420054
rect 94586 419498 94822 419734
rect 94586 383818 94822 384054
rect 94586 383498 94822 383734
rect 94586 347818 94822 348054
rect 94586 347498 94822 347734
rect 94586 311818 94822 312054
rect 94586 311498 94822 311734
rect 94586 275818 94822 276054
rect 94586 275498 94822 275734
rect 94586 239818 94822 240054
rect 94586 239498 94822 239734
rect 94586 203818 94822 204054
rect 94586 203498 94822 203734
rect 94586 167818 94822 168054
rect 94586 167498 94822 167734
rect 94586 131818 94822 132054
rect 94586 131498 94822 131734
rect 94586 95818 94822 96054
rect 94586 95498 94822 95734
rect 94586 59818 94822 60054
rect 94586 59498 94822 59734
rect 94586 23818 94822 24054
rect 94586 23498 94822 23734
rect 94586 -3342 94822 -3106
rect 94586 -3662 94822 -3426
rect 98186 675418 98422 675654
rect 98186 675098 98422 675334
rect 98186 639418 98422 639654
rect 98186 639098 98422 639334
rect 98186 603418 98422 603654
rect 98186 603098 98422 603334
rect 98186 567418 98422 567654
rect 98186 567098 98422 567334
rect 98186 531418 98422 531654
rect 98186 531098 98422 531334
rect 98186 495418 98422 495654
rect 98186 495098 98422 495334
rect 98186 459418 98422 459654
rect 98186 459098 98422 459334
rect 98186 423418 98422 423654
rect 98186 423098 98422 423334
rect 98186 387418 98422 387654
rect 98186 387098 98422 387334
rect 98186 351418 98422 351654
rect 98186 351098 98422 351334
rect 98186 315418 98422 315654
rect 98186 315098 98422 315334
rect 98186 279418 98422 279654
rect 98186 279098 98422 279334
rect 98186 243418 98422 243654
rect 98186 243098 98422 243334
rect 98186 207418 98422 207654
rect 98186 207098 98422 207334
rect 98186 171418 98422 171654
rect 98186 171098 98422 171334
rect 98186 135418 98422 135654
rect 98186 135098 98422 135334
rect 98186 99418 98422 99654
rect 98186 99098 98422 99334
rect 98186 63418 98422 63654
rect 98186 63098 98422 63334
rect 98186 27418 98422 27654
rect 98186 27098 98422 27334
rect 98186 -5182 98422 -4946
rect 98186 -5502 98422 -5266
rect 119786 710122 120022 710358
rect 119786 709802 120022 710038
rect 116186 708282 116422 708518
rect 116186 707962 116422 708198
rect 112586 706442 112822 706678
rect 112586 706122 112822 706358
rect 101786 679018 102022 679254
rect 101786 678698 102022 678934
rect 101786 643018 102022 643254
rect 101786 642698 102022 642934
rect 101786 607018 102022 607254
rect 101786 606698 102022 606934
rect 101786 571018 102022 571254
rect 101786 570698 102022 570934
rect 108986 704602 109222 704838
rect 108986 704282 109222 704518
rect 108986 686218 109222 686454
rect 108986 685898 109222 686134
rect 108986 650218 109222 650454
rect 108986 649898 109222 650134
rect 108986 614218 109222 614454
rect 108986 613898 109222 614134
rect 108986 578218 109222 578454
rect 108986 577898 109222 578134
rect 108350 561372 108586 561458
rect 108350 561308 108436 561372
rect 108436 561308 108500 561372
rect 108500 561308 108586 561372
rect 108350 561222 108586 561308
rect 101786 535018 102022 535254
rect 101786 534698 102022 534934
rect 101786 499018 102022 499254
rect 101786 498698 102022 498934
rect 101786 463018 102022 463254
rect 101786 462698 102022 462934
rect 101786 427018 102022 427254
rect 101786 426698 102022 426934
rect 101786 391018 102022 391254
rect 101786 390698 102022 390934
rect 101786 355018 102022 355254
rect 101786 354698 102022 354934
rect 101786 319018 102022 319254
rect 101786 318698 102022 318934
rect 101786 283018 102022 283254
rect 101786 282698 102022 282934
rect 101786 247018 102022 247254
rect 101786 246698 102022 246934
rect 101786 211018 102022 211254
rect 101786 210698 102022 210934
rect 101786 175018 102022 175254
rect 101786 174698 102022 174934
rect 101786 139018 102022 139254
rect 101786 138698 102022 138934
rect 101786 103018 102022 103254
rect 101786 102698 102022 102934
rect 101786 67018 102022 67254
rect 101786 66698 102022 66934
rect 101786 31018 102022 31254
rect 101786 30698 102022 30934
rect 83786 -6102 84022 -5866
rect 83786 -6422 84022 -6186
rect 112586 689818 112822 690054
rect 112586 689498 112822 689734
rect 112586 653818 112822 654054
rect 112586 653498 112822 653734
rect 112586 617818 112822 618054
rect 112586 617498 112822 617734
rect 112586 581818 112822 582054
rect 112586 581498 112822 581734
rect 109638 561372 109874 561458
rect 109638 561308 109724 561372
rect 109724 561308 109788 561372
rect 109788 561308 109874 561372
rect 109638 561222 109874 561308
rect 108986 542218 109222 542454
rect 108986 541898 109222 542134
rect 108986 506218 109222 506454
rect 108986 505898 109222 506134
rect 108986 470218 109222 470454
rect 108986 469898 109222 470134
rect 108986 434218 109222 434454
rect 108986 433898 109222 434134
rect 108986 398218 109222 398454
rect 108986 397898 109222 398134
rect 108986 362218 109222 362454
rect 108986 361898 109222 362134
rect 108986 326218 109222 326454
rect 108986 325898 109222 326134
rect 108986 290218 109222 290454
rect 108986 289898 109222 290134
rect 108986 254218 109222 254454
rect 108986 253898 109222 254134
rect 108986 218218 109222 218454
rect 108986 217898 109222 218134
rect 108986 182218 109222 182454
rect 108986 181898 109222 182134
rect 108986 146218 109222 146454
rect 108986 145898 109222 146134
rect 108986 110218 109222 110454
rect 108986 109898 109222 110134
rect 108986 74218 109222 74454
rect 108986 73898 109222 74134
rect 108986 38218 109222 38454
rect 108986 37898 109222 38134
rect 108986 2218 109222 2454
rect 108986 1898 109222 2134
rect 108986 -582 109222 -346
rect 108986 -902 109222 -666
rect 112586 545818 112822 546054
rect 112586 545498 112822 545734
rect 112586 509818 112822 510054
rect 112586 509498 112822 509734
rect 112586 473818 112822 474054
rect 112586 473498 112822 473734
rect 112586 437818 112822 438054
rect 112586 437498 112822 437734
rect 112586 401818 112822 402054
rect 112586 401498 112822 401734
rect 112586 365818 112822 366054
rect 112586 365498 112822 365734
rect 112586 329818 112822 330054
rect 112586 329498 112822 329734
rect 112586 293818 112822 294054
rect 112586 293498 112822 293734
rect 112586 257818 112822 258054
rect 112586 257498 112822 257734
rect 112586 221818 112822 222054
rect 112586 221498 112822 221734
rect 112586 185818 112822 186054
rect 112586 185498 112822 185734
rect 112586 149818 112822 150054
rect 112586 149498 112822 149734
rect 112586 113818 112822 114054
rect 112586 113498 112822 113734
rect 112586 77818 112822 78054
rect 112586 77498 112822 77734
rect 112586 41818 112822 42054
rect 112586 41498 112822 41734
rect 112586 5818 112822 6054
rect 112586 5498 112822 5734
rect 112586 -2422 112822 -2186
rect 112586 -2742 112822 -2506
rect 116186 693418 116422 693654
rect 116186 693098 116422 693334
rect 116186 657418 116422 657654
rect 116186 657098 116422 657334
rect 116186 621418 116422 621654
rect 116186 621098 116422 621334
rect 116186 585418 116422 585654
rect 116186 585098 116422 585334
rect 137786 711042 138022 711278
rect 137786 710722 138022 710958
rect 134186 709202 134422 709438
rect 134186 708882 134422 709118
rect 130586 707362 130822 707598
rect 130586 707042 130822 707278
rect 119786 697018 120022 697254
rect 119786 696698 120022 696934
rect 119786 661018 120022 661254
rect 119786 660698 120022 660934
rect 119786 625018 120022 625254
rect 119786 624698 120022 624934
rect 119786 589018 120022 589254
rect 119786 588698 120022 588934
rect 117550 561372 117786 561458
rect 117550 561308 117636 561372
rect 117636 561308 117700 561372
rect 117700 561308 117786 561372
rect 117550 561222 117786 561308
rect 116186 549418 116422 549654
rect 116186 549098 116422 549334
rect 116186 513418 116422 513654
rect 116186 513098 116422 513334
rect 116186 477418 116422 477654
rect 116186 477098 116422 477334
rect 116186 441418 116422 441654
rect 116186 441098 116422 441334
rect 116186 405418 116422 405654
rect 116186 405098 116422 405334
rect 116186 369418 116422 369654
rect 116186 369098 116422 369334
rect 116186 333418 116422 333654
rect 116186 333098 116422 333334
rect 116186 297418 116422 297654
rect 116186 297098 116422 297334
rect 116186 261418 116422 261654
rect 116186 261098 116422 261334
rect 116186 225418 116422 225654
rect 116186 225098 116422 225334
rect 116186 189418 116422 189654
rect 116186 189098 116422 189334
rect 116186 153418 116422 153654
rect 116186 153098 116422 153334
rect 116186 117418 116422 117654
rect 116186 117098 116422 117334
rect 116186 81418 116422 81654
rect 116186 81098 116422 81334
rect 116186 45418 116422 45654
rect 116186 45098 116422 45334
rect 116186 9418 116422 9654
rect 116186 9098 116422 9334
rect 116186 -4262 116422 -4026
rect 116186 -4582 116422 -4346
rect 126986 705522 127222 705758
rect 126986 705202 127222 705438
rect 126986 668218 127222 668454
rect 126986 667898 127222 668134
rect 126986 632218 127222 632454
rect 126986 631898 127222 632134
rect 126986 596218 127222 596454
rect 126986 595898 127222 596134
rect 120678 562582 120914 562818
rect 125462 562732 125698 562818
rect 125462 562668 125548 562732
rect 125548 562668 125612 562732
rect 125612 562668 125698 562732
rect 125462 562582 125698 562668
rect 119786 553018 120022 553254
rect 119786 552698 120022 552934
rect 119786 517018 120022 517254
rect 119786 516698 120022 516934
rect 119786 481018 120022 481254
rect 119786 480698 120022 480934
rect 119786 445018 120022 445254
rect 119786 444698 120022 444934
rect 119786 409018 120022 409254
rect 119786 408698 120022 408934
rect 119786 373018 120022 373254
rect 119786 372698 120022 372934
rect 119786 337018 120022 337254
rect 119786 336698 120022 336934
rect 119786 301018 120022 301254
rect 119786 300698 120022 300934
rect 119786 265018 120022 265254
rect 119786 264698 120022 264934
rect 119786 229018 120022 229254
rect 119786 228698 120022 228934
rect 119786 193018 120022 193254
rect 119786 192698 120022 192934
rect 119786 157018 120022 157254
rect 119786 156698 120022 156934
rect 119786 121018 120022 121254
rect 119786 120698 120022 120934
rect 119786 85018 120022 85254
rect 119786 84698 120022 84934
rect 119786 49018 120022 49254
rect 119786 48698 120022 48934
rect 119786 13018 120022 13254
rect 119786 12698 120022 12934
rect 101786 -7022 102022 -6786
rect 101786 -7342 102022 -7106
rect 126986 560218 127222 560454
rect 126986 559898 127222 560134
rect 126986 524218 127222 524454
rect 126986 523898 127222 524134
rect 126986 488218 127222 488454
rect 126986 487898 127222 488134
rect 126986 452218 127222 452454
rect 126986 451898 127222 452134
rect 126986 416218 127222 416454
rect 126986 415898 127222 416134
rect 126986 380218 127222 380454
rect 126986 379898 127222 380134
rect 126986 344218 127222 344454
rect 126986 343898 127222 344134
rect 126986 308218 127222 308454
rect 126986 307898 127222 308134
rect 126986 272218 127222 272454
rect 126986 271898 127222 272134
rect 126986 236218 127222 236454
rect 126986 235898 127222 236134
rect 126986 200218 127222 200454
rect 126986 199898 127222 200134
rect 126986 164218 127222 164454
rect 126986 163898 127222 164134
rect 126986 128218 127222 128454
rect 126986 127898 127222 128134
rect 126986 92218 127222 92454
rect 126986 91898 127222 92134
rect 126986 56218 127222 56454
rect 126986 55898 127222 56134
rect 126986 20218 127222 20454
rect 126986 19898 127222 20134
rect 126986 -1502 127222 -1266
rect 126986 -1822 127222 -1586
rect 130586 671818 130822 672054
rect 130586 671498 130822 671734
rect 130586 635818 130822 636054
rect 130586 635498 130822 635734
rect 130586 599818 130822 600054
rect 130586 599498 130822 599734
rect 130586 563818 130822 564054
rect 130586 563498 130822 563734
rect 130586 527818 130822 528054
rect 130586 527498 130822 527734
rect 130586 491818 130822 492054
rect 130586 491498 130822 491734
rect 130586 455818 130822 456054
rect 130586 455498 130822 455734
rect 130586 419818 130822 420054
rect 130586 419498 130822 419734
rect 130586 383818 130822 384054
rect 130586 383498 130822 383734
rect 130586 347818 130822 348054
rect 130586 347498 130822 347734
rect 130586 311818 130822 312054
rect 130586 311498 130822 311734
rect 130586 275818 130822 276054
rect 130586 275498 130822 275734
rect 130586 239818 130822 240054
rect 130586 239498 130822 239734
rect 130586 203818 130822 204054
rect 130586 203498 130822 203734
rect 130586 167818 130822 168054
rect 130586 167498 130822 167734
rect 130586 131818 130822 132054
rect 130586 131498 130822 131734
rect 130586 95818 130822 96054
rect 130586 95498 130822 95734
rect 130586 59818 130822 60054
rect 130586 59498 130822 59734
rect 130586 23818 130822 24054
rect 130586 23498 130822 23734
rect 130586 -3342 130822 -3106
rect 130586 -3662 130822 -3426
rect 134186 675418 134422 675654
rect 134186 675098 134422 675334
rect 134186 639418 134422 639654
rect 134186 639098 134422 639334
rect 134186 603418 134422 603654
rect 134186 603098 134422 603334
rect 134186 567418 134422 567654
rect 134186 567098 134422 567334
rect 155786 710122 156022 710358
rect 155786 709802 156022 710038
rect 152186 708282 152422 708518
rect 152186 707962 152422 708198
rect 148586 706442 148822 706678
rect 148586 706122 148822 706358
rect 137786 679018 138022 679254
rect 137786 678698 138022 678934
rect 137786 643018 138022 643254
rect 137786 642698 138022 642934
rect 137786 607018 138022 607254
rect 137786 606698 138022 606934
rect 137786 571018 138022 571254
rect 137786 570698 138022 570934
rect 135030 561222 135266 561458
rect 135582 561372 135818 561458
rect 135582 561308 135668 561372
rect 135668 561308 135732 561372
rect 135732 561308 135818 561372
rect 135582 561222 135818 561308
rect 134186 531418 134422 531654
rect 134186 531098 134422 531334
rect 134186 495418 134422 495654
rect 134186 495098 134422 495334
rect 134186 459418 134422 459654
rect 134186 459098 134422 459334
rect 134186 423418 134422 423654
rect 134186 423098 134422 423334
rect 134186 387418 134422 387654
rect 134186 387098 134422 387334
rect 134186 351418 134422 351654
rect 134186 351098 134422 351334
rect 134186 315418 134422 315654
rect 134186 315098 134422 315334
rect 134186 279418 134422 279654
rect 134186 279098 134422 279334
rect 134186 243418 134422 243654
rect 134186 243098 134422 243334
rect 134186 207418 134422 207654
rect 134186 207098 134422 207334
rect 134186 171418 134422 171654
rect 134186 171098 134422 171334
rect 134186 135418 134422 135654
rect 134186 135098 134422 135334
rect 134186 99418 134422 99654
rect 134186 99098 134422 99334
rect 134186 63418 134422 63654
rect 134186 63098 134422 63334
rect 134186 27418 134422 27654
rect 134186 27098 134422 27334
rect 134186 -5182 134422 -4946
rect 134186 -5502 134422 -5266
rect 144986 704602 145222 704838
rect 144986 704282 145222 704518
rect 144986 686218 145222 686454
rect 144986 685898 145222 686134
rect 144986 650218 145222 650454
rect 144986 649898 145222 650134
rect 144986 614218 145222 614454
rect 144986 613898 145222 614134
rect 144986 578218 145222 578454
rect 144986 577898 145222 578134
rect 139998 562582 140234 562818
rect 137786 535018 138022 535254
rect 137786 534698 138022 534934
rect 137786 499018 138022 499254
rect 137786 498698 138022 498934
rect 137786 463018 138022 463254
rect 137786 462698 138022 462934
rect 137786 427018 138022 427254
rect 137786 426698 138022 426934
rect 137786 391018 138022 391254
rect 137786 390698 138022 390934
rect 137786 355018 138022 355254
rect 137786 354698 138022 354934
rect 137786 319018 138022 319254
rect 137786 318698 138022 318934
rect 137786 283018 138022 283254
rect 137786 282698 138022 282934
rect 137786 247018 138022 247254
rect 137786 246698 138022 246934
rect 137786 211018 138022 211254
rect 137786 210698 138022 210934
rect 137786 175018 138022 175254
rect 137786 174698 138022 174934
rect 137786 139018 138022 139254
rect 137786 138698 138022 138934
rect 137786 103018 138022 103254
rect 137786 102698 138022 102934
rect 137786 67018 138022 67254
rect 137786 66698 138022 66934
rect 137786 31018 138022 31254
rect 137786 30698 138022 30934
rect 119786 -6102 120022 -5866
rect 119786 -6422 120022 -6186
rect 148586 689818 148822 690054
rect 148586 689498 148822 689734
rect 148586 653818 148822 654054
rect 148586 653498 148822 653734
rect 148586 617818 148822 618054
rect 148586 617498 148822 617734
rect 148586 581818 148822 582054
rect 148586 581498 148822 581734
rect 147358 561372 147594 561458
rect 147358 561308 147444 561372
rect 147444 561308 147508 561372
rect 147508 561308 147594 561372
rect 147358 561222 147594 561308
rect 144986 542218 145222 542454
rect 144986 541898 145222 542134
rect 144986 506218 145222 506454
rect 144986 505898 145222 506134
rect 144986 470218 145222 470454
rect 144986 469898 145222 470134
rect 144986 434218 145222 434454
rect 144986 433898 145222 434134
rect 144986 398218 145222 398454
rect 144986 397898 145222 398134
rect 144986 362218 145222 362454
rect 144986 361898 145222 362134
rect 144986 326218 145222 326454
rect 144986 325898 145222 326134
rect 144986 290218 145222 290454
rect 144986 289898 145222 290134
rect 144986 254218 145222 254454
rect 144986 253898 145222 254134
rect 144986 218218 145222 218454
rect 144986 217898 145222 218134
rect 144986 182218 145222 182454
rect 144986 181898 145222 182134
rect 144986 146218 145222 146454
rect 144986 145898 145222 146134
rect 144986 110218 145222 110454
rect 144986 109898 145222 110134
rect 144986 74218 145222 74454
rect 144986 73898 145222 74134
rect 144986 38218 145222 38454
rect 144986 37898 145222 38134
rect 144986 2218 145222 2454
rect 144986 1898 145222 2134
rect 144986 -582 145222 -346
rect 144986 -902 145222 -666
rect 148586 545818 148822 546054
rect 148586 545498 148822 545734
rect 148586 509818 148822 510054
rect 148586 509498 148822 509734
rect 148586 473818 148822 474054
rect 148586 473498 148822 473734
rect 148586 437818 148822 438054
rect 148586 437498 148822 437734
rect 148586 401818 148822 402054
rect 148586 401498 148822 401734
rect 148586 365818 148822 366054
rect 148586 365498 148822 365734
rect 148586 329818 148822 330054
rect 148586 329498 148822 329734
rect 148586 293818 148822 294054
rect 148586 293498 148822 293734
rect 148586 257818 148822 258054
rect 148586 257498 148822 257734
rect 148586 221818 148822 222054
rect 148586 221498 148822 221734
rect 148586 185818 148822 186054
rect 148586 185498 148822 185734
rect 148586 149818 148822 150054
rect 148586 149498 148822 149734
rect 148586 113818 148822 114054
rect 148586 113498 148822 113734
rect 148586 77818 148822 78054
rect 148586 77498 148822 77734
rect 148586 41818 148822 42054
rect 148586 41498 148822 41734
rect 148586 5818 148822 6054
rect 148586 5498 148822 5734
rect 148586 -2422 148822 -2186
rect 148586 -2742 148822 -2506
rect 152186 693418 152422 693654
rect 152186 693098 152422 693334
rect 152186 657418 152422 657654
rect 152186 657098 152422 657334
rect 152186 621418 152422 621654
rect 152186 621098 152422 621334
rect 152186 585418 152422 585654
rect 152186 585098 152422 585334
rect 173786 711042 174022 711278
rect 173786 710722 174022 710958
rect 170186 709202 170422 709438
rect 170186 708882 170422 709118
rect 166586 707362 166822 707598
rect 166586 707042 166822 707278
rect 155786 697018 156022 697254
rect 155786 696698 156022 696934
rect 155786 661018 156022 661254
rect 155786 660698 156022 660934
rect 155786 625018 156022 625254
rect 155786 624698 156022 624934
rect 155786 589018 156022 589254
rect 155786 588698 156022 588934
rect 154350 561372 154586 561458
rect 154350 561308 154436 561372
rect 154436 561308 154500 561372
rect 154500 561308 154586 561372
rect 154350 561222 154586 561308
rect 154902 561372 155138 561458
rect 154902 561308 154988 561372
rect 154988 561308 155052 561372
rect 155052 561308 155138 561372
rect 154902 561222 155138 561308
rect 152186 549418 152422 549654
rect 152186 549098 152422 549334
rect 152186 513418 152422 513654
rect 152186 513098 152422 513334
rect 152186 477418 152422 477654
rect 152186 477098 152422 477334
rect 152186 441418 152422 441654
rect 152186 441098 152422 441334
rect 152186 405418 152422 405654
rect 152186 405098 152422 405334
rect 152186 369418 152422 369654
rect 152186 369098 152422 369334
rect 152186 333418 152422 333654
rect 152186 333098 152422 333334
rect 152186 297418 152422 297654
rect 152186 297098 152422 297334
rect 152186 261418 152422 261654
rect 152186 261098 152422 261334
rect 152186 225418 152422 225654
rect 152186 225098 152422 225334
rect 152186 189418 152422 189654
rect 152186 189098 152422 189334
rect 152186 153418 152422 153654
rect 152186 153098 152422 153334
rect 152186 117418 152422 117654
rect 152186 117098 152422 117334
rect 152186 81418 152422 81654
rect 152186 81098 152422 81334
rect 152186 45418 152422 45654
rect 152186 45098 152422 45334
rect 152186 9418 152422 9654
rect 152186 9098 152422 9334
rect 152186 -4262 152422 -4026
rect 152186 -4582 152422 -4346
rect 162986 705522 163222 705758
rect 162986 705202 163222 705438
rect 162986 668218 163222 668454
rect 162986 667898 163222 668134
rect 162986 632218 163222 632454
rect 162986 631898 163222 632134
rect 162986 596218 163222 596454
rect 162986 595898 163222 596134
rect 159318 562582 159554 562818
rect 155786 553018 156022 553254
rect 155786 552698 156022 552934
rect 155786 517018 156022 517254
rect 155786 516698 156022 516934
rect 155786 481018 156022 481254
rect 155786 480698 156022 480934
rect 155786 445018 156022 445254
rect 155786 444698 156022 444934
rect 155786 409018 156022 409254
rect 155786 408698 156022 408934
rect 155786 373018 156022 373254
rect 155786 372698 156022 372934
rect 155786 337018 156022 337254
rect 155786 336698 156022 336934
rect 155786 301018 156022 301254
rect 155786 300698 156022 300934
rect 155786 265018 156022 265254
rect 155786 264698 156022 264934
rect 155786 229018 156022 229254
rect 155786 228698 156022 228934
rect 155786 193018 156022 193254
rect 155786 192698 156022 192934
rect 155786 157018 156022 157254
rect 155786 156698 156022 156934
rect 155786 121018 156022 121254
rect 155786 120698 156022 120934
rect 155786 85018 156022 85254
rect 155786 84698 156022 84934
rect 155786 49018 156022 49254
rect 155786 48698 156022 48934
rect 155786 13018 156022 13254
rect 155786 12698 156022 12934
rect 137786 -7022 138022 -6786
rect 137786 -7342 138022 -7106
rect 166586 671818 166822 672054
rect 166586 671498 166822 671734
rect 166586 635818 166822 636054
rect 166586 635498 166822 635734
rect 166586 599818 166822 600054
rect 166586 599498 166822 599734
rect 166586 563818 166822 564054
rect 166586 563498 166822 563734
rect 164102 562732 164338 562818
rect 164102 562668 164188 562732
rect 164188 562668 164252 562732
rect 164252 562668 164338 562732
rect 164102 562582 164338 562668
rect 162986 560218 163222 560454
rect 162986 559898 163222 560134
rect 162986 524218 163222 524454
rect 162986 523898 163222 524134
rect 162986 488218 163222 488454
rect 162986 487898 163222 488134
rect 162986 452218 163222 452454
rect 162986 451898 163222 452134
rect 162986 416218 163222 416454
rect 162986 415898 163222 416134
rect 162986 380218 163222 380454
rect 162986 379898 163222 380134
rect 162986 344218 163222 344454
rect 162986 343898 163222 344134
rect 162986 308218 163222 308454
rect 162986 307898 163222 308134
rect 162986 272218 163222 272454
rect 162986 271898 163222 272134
rect 162986 236218 163222 236454
rect 162986 235898 163222 236134
rect 162986 200218 163222 200454
rect 162986 199898 163222 200134
rect 162986 164218 163222 164454
rect 162986 163898 163222 164134
rect 162986 128218 163222 128454
rect 162986 127898 163222 128134
rect 162986 92218 163222 92454
rect 162986 91898 163222 92134
rect 162986 56218 163222 56454
rect 162986 55898 163222 56134
rect 162986 20218 163222 20454
rect 162986 19898 163222 20134
rect 162986 -1502 163222 -1266
rect 162986 -1822 163222 -1586
rect 170186 675418 170422 675654
rect 170186 675098 170422 675334
rect 170186 639418 170422 639654
rect 170186 639098 170422 639334
rect 170186 603418 170422 603654
rect 170186 603098 170422 603334
rect 170186 567418 170422 567654
rect 170186 567098 170422 567334
rect 167230 562732 167466 562818
rect 167230 562668 167316 562732
rect 167316 562668 167380 562732
rect 167380 562668 167466 562732
rect 167230 562582 167466 562668
rect 166586 527818 166822 528054
rect 166586 527498 166822 527734
rect 166586 491818 166822 492054
rect 166586 491498 166822 491734
rect 166586 455818 166822 456054
rect 166586 455498 166822 455734
rect 166586 419818 166822 420054
rect 166586 419498 166822 419734
rect 166586 383818 166822 384054
rect 166586 383498 166822 383734
rect 166586 347818 166822 348054
rect 166586 347498 166822 347734
rect 166586 311818 166822 312054
rect 166586 311498 166822 311734
rect 166586 275818 166822 276054
rect 166586 275498 166822 275734
rect 166586 239818 166822 240054
rect 166586 239498 166822 239734
rect 166586 203818 166822 204054
rect 166586 203498 166822 203734
rect 166586 167818 166822 168054
rect 166586 167498 166822 167734
rect 166586 131818 166822 132054
rect 166586 131498 166822 131734
rect 166586 95818 166822 96054
rect 166586 95498 166822 95734
rect 166586 59818 166822 60054
rect 166586 59498 166822 59734
rect 166586 23818 166822 24054
rect 166586 23498 166822 23734
rect 166586 -3342 166822 -3106
rect 166586 -3662 166822 -3426
rect 170186 531418 170422 531654
rect 170186 531098 170422 531334
rect 170186 495418 170422 495654
rect 170186 495098 170422 495334
rect 170186 459418 170422 459654
rect 170186 459098 170422 459334
rect 170186 423418 170422 423654
rect 170186 423098 170422 423334
rect 170186 387418 170422 387654
rect 170186 387098 170422 387334
rect 170186 351418 170422 351654
rect 170186 351098 170422 351334
rect 170186 315418 170422 315654
rect 170186 315098 170422 315334
rect 170186 279418 170422 279654
rect 170186 279098 170422 279334
rect 170186 243418 170422 243654
rect 170186 243098 170422 243334
rect 170186 207418 170422 207654
rect 170186 207098 170422 207334
rect 170186 171418 170422 171654
rect 170186 171098 170422 171334
rect 170186 135418 170422 135654
rect 170186 135098 170422 135334
rect 170186 99418 170422 99654
rect 170186 99098 170422 99334
rect 170186 63418 170422 63654
rect 170186 63098 170422 63334
rect 170186 27418 170422 27654
rect 170186 27098 170422 27334
rect 170186 -5182 170422 -4946
rect 170186 -5502 170422 -5266
rect 191786 710122 192022 710358
rect 191786 709802 192022 710038
rect 188186 708282 188422 708518
rect 188186 707962 188422 708198
rect 184586 706442 184822 706678
rect 184586 706122 184822 706358
rect 173786 679018 174022 679254
rect 173786 678698 174022 678934
rect 173786 643018 174022 643254
rect 173786 642698 174022 642934
rect 173786 607018 174022 607254
rect 173786 606698 174022 606934
rect 173786 571018 174022 571254
rect 173786 570698 174022 570934
rect 180986 704602 181222 704838
rect 180986 704282 181222 704518
rect 180986 686218 181222 686454
rect 180986 685898 181222 686134
rect 180986 650218 181222 650454
rect 180986 649898 181222 650134
rect 180986 614218 181222 614454
rect 180986 613898 181222 614134
rect 180986 578218 181222 578454
rect 180986 577898 181222 578134
rect 178638 562582 178874 562818
rect 176062 561372 176298 561458
rect 176062 561308 176148 561372
rect 176148 561308 176212 561372
rect 176212 561308 176298 561372
rect 176062 561222 176298 561308
rect 173786 535018 174022 535254
rect 173786 534698 174022 534934
rect 173786 499018 174022 499254
rect 173786 498698 174022 498934
rect 173786 463018 174022 463254
rect 173786 462698 174022 462934
rect 173786 427018 174022 427254
rect 173786 426698 174022 426934
rect 173786 391018 174022 391254
rect 173786 390698 174022 390934
rect 173786 355018 174022 355254
rect 173786 354698 174022 354934
rect 173786 319018 174022 319254
rect 173786 318698 174022 318934
rect 173786 283018 174022 283254
rect 173786 282698 174022 282934
rect 173786 247018 174022 247254
rect 173786 246698 174022 246934
rect 173786 211018 174022 211254
rect 173786 210698 174022 210934
rect 173786 175018 174022 175254
rect 173786 174698 174022 174934
rect 173786 139018 174022 139254
rect 173786 138698 174022 138934
rect 173786 103018 174022 103254
rect 173786 102698 174022 102934
rect 173786 67018 174022 67254
rect 173786 66698 174022 66934
rect 173786 31018 174022 31254
rect 173786 30698 174022 30934
rect 155786 -6102 156022 -5866
rect 155786 -6422 156022 -6186
rect 184586 689818 184822 690054
rect 184586 689498 184822 689734
rect 184586 653818 184822 654054
rect 184586 653498 184822 653734
rect 184586 617818 184822 618054
rect 184586 617498 184822 617734
rect 184586 581818 184822 582054
rect 184586 581498 184822 581734
rect 183422 562732 183658 562818
rect 183422 562668 183508 562732
rect 183508 562668 183572 562732
rect 183572 562668 183658 562732
rect 183422 562582 183658 562668
rect 180986 542218 181222 542454
rect 180986 541898 181222 542134
rect 180986 506218 181222 506454
rect 180986 505898 181222 506134
rect 180986 470218 181222 470454
rect 180986 469898 181222 470134
rect 180986 434218 181222 434454
rect 180986 433898 181222 434134
rect 180986 398218 181222 398454
rect 180986 397898 181222 398134
rect 180986 362218 181222 362454
rect 180986 361898 181222 362134
rect 180986 326218 181222 326454
rect 180986 325898 181222 326134
rect 180986 290218 181222 290454
rect 180986 289898 181222 290134
rect 180986 254218 181222 254454
rect 180986 253898 181222 254134
rect 180986 218218 181222 218454
rect 180986 217898 181222 218134
rect 180986 182218 181222 182454
rect 180986 181898 181222 182134
rect 180986 146218 181222 146454
rect 180986 145898 181222 146134
rect 180986 110218 181222 110454
rect 180986 109898 181222 110134
rect 180986 74218 181222 74454
rect 180986 73898 181222 74134
rect 180986 38218 181222 38454
rect 180986 37898 181222 38134
rect 180986 2218 181222 2454
rect 180986 1898 181222 2134
rect 180986 -582 181222 -346
rect 180986 -902 181222 -666
rect 184586 545818 184822 546054
rect 184586 545498 184822 545734
rect 184586 509818 184822 510054
rect 184586 509498 184822 509734
rect 184586 473818 184822 474054
rect 184586 473498 184822 473734
rect 184586 437818 184822 438054
rect 184586 437498 184822 437734
rect 184586 401818 184822 402054
rect 184586 401498 184822 401734
rect 184586 365818 184822 366054
rect 184586 365498 184822 365734
rect 184586 329818 184822 330054
rect 184586 329498 184822 329734
rect 184586 293818 184822 294054
rect 184586 293498 184822 293734
rect 184586 257818 184822 258054
rect 184586 257498 184822 257734
rect 184586 221818 184822 222054
rect 184586 221498 184822 221734
rect 184586 185818 184822 186054
rect 184586 185498 184822 185734
rect 184586 149818 184822 150054
rect 184586 149498 184822 149734
rect 184586 113818 184822 114054
rect 184586 113498 184822 113734
rect 184586 77818 184822 78054
rect 184586 77498 184822 77734
rect 184586 41818 184822 42054
rect 184586 41498 184822 41734
rect 184586 5818 184822 6054
rect 184586 5498 184822 5734
rect 184586 -2422 184822 -2186
rect 184586 -2742 184822 -2506
rect 188186 693418 188422 693654
rect 188186 693098 188422 693334
rect 188186 657418 188422 657654
rect 188186 657098 188422 657334
rect 188186 621418 188422 621654
rect 188186 621098 188422 621334
rect 188186 585418 188422 585654
rect 188186 585098 188422 585334
rect 188186 549418 188422 549654
rect 188186 549098 188422 549334
rect 188186 513418 188422 513654
rect 188186 513098 188422 513334
rect 188186 477418 188422 477654
rect 188186 477098 188422 477334
rect 188186 441418 188422 441654
rect 188186 441098 188422 441334
rect 188186 405418 188422 405654
rect 188186 405098 188422 405334
rect 188186 369418 188422 369654
rect 188186 369098 188422 369334
rect 188186 333418 188422 333654
rect 188186 333098 188422 333334
rect 188186 297418 188422 297654
rect 188186 297098 188422 297334
rect 188186 261418 188422 261654
rect 188186 261098 188422 261334
rect 188186 225418 188422 225654
rect 188186 225098 188422 225334
rect 188186 189418 188422 189654
rect 188186 189098 188422 189334
rect 188186 153418 188422 153654
rect 188186 153098 188422 153334
rect 188186 117418 188422 117654
rect 188186 117098 188422 117334
rect 188186 81418 188422 81654
rect 188186 81098 188422 81334
rect 188186 45418 188422 45654
rect 188186 45098 188422 45334
rect 188186 9418 188422 9654
rect 188186 9098 188422 9334
rect 188186 -4262 188422 -4026
rect 188186 -4582 188422 -4346
rect 209786 711042 210022 711278
rect 209786 710722 210022 710958
rect 206186 709202 206422 709438
rect 206186 708882 206422 709118
rect 202586 707362 202822 707598
rect 202586 707042 202822 707278
rect 191786 697018 192022 697254
rect 191786 696698 192022 696934
rect 191786 661018 192022 661254
rect 191786 660698 192022 660934
rect 191786 625018 192022 625254
rect 191786 624698 192022 624934
rect 191786 589018 192022 589254
rect 191786 588698 192022 588934
rect 198986 705522 199222 705758
rect 198986 705202 199222 705438
rect 198986 668218 199222 668454
rect 198986 667898 199222 668134
rect 198986 632218 199222 632454
rect 198986 631898 199222 632134
rect 198986 596218 199222 596454
rect 198986 595898 199222 596134
rect 196670 562582 196906 562818
rect 192990 561222 193226 561458
rect 193542 561372 193778 561458
rect 193542 561308 193628 561372
rect 193628 561308 193692 561372
rect 193692 561308 193778 561372
rect 193542 561222 193778 561308
rect 191786 553018 192022 553254
rect 191786 552698 192022 552934
rect 191786 517018 192022 517254
rect 191786 516698 192022 516934
rect 191786 481018 192022 481254
rect 191786 480698 192022 480934
rect 191786 445018 192022 445254
rect 191786 444698 192022 444934
rect 191786 409018 192022 409254
rect 191786 408698 192022 408934
rect 191786 373018 192022 373254
rect 191786 372698 192022 372934
rect 191786 337018 192022 337254
rect 191786 336698 192022 336934
rect 191786 301018 192022 301254
rect 191786 300698 192022 300934
rect 191786 265018 192022 265254
rect 191786 264698 192022 264934
rect 191786 229018 192022 229254
rect 191786 228698 192022 228934
rect 191786 193018 192022 193254
rect 191786 192698 192022 192934
rect 191786 157018 192022 157254
rect 191786 156698 192022 156934
rect 191786 121018 192022 121254
rect 191786 120698 192022 120934
rect 191786 85018 192022 85254
rect 191786 84698 192022 84934
rect 191786 49018 192022 49254
rect 191786 48698 192022 48934
rect 191786 13018 192022 13254
rect 191786 12698 192022 12934
rect 173786 -7022 174022 -6786
rect 173786 -7342 174022 -7106
rect 198986 560218 199222 560454
rect 198986 559898 199222 560134
rect 198986 524218 199222 524454
rect 198986 523898 199222 524134
rect 198986 488218 199222 488454
rect 198986 487898 199222 488134
rect 198986 452218 199222 452454
rect 198986 451898 199222 452134
rect 198986 416218 199222 416454
rect 198986 415898 199222 416134
rect 198986 380218 199222 380454
rect 198986 379898 199222 380134
rect 198986 344218 199222 344454
rect 198986 343898 199222 344134
rect 198986 308218 199222 308454
rect 198986 307898 199222 308134
rect 198986 272218 199222 272454
rect 198986 271898 199222 272134
rect 198986 236218 199222 236454
rect 198986 235898 199222 236134
rect 198986 200218 199222 200454
rect 198986 199898 199222 200134
rect 198986 164218 199222 164454
rect 198986 163898 199222 164134
rect 198986 128218 199222 128454
rect 198986 127898 199222 128134
rect 198986 92218 199222 92454
rect 198986 91898 199222 92134
rect 198986 56218 199222 56454
rect 198986 55898 199222 56134
rect 198986 20218 199222 20454
rect 198986 19898 199222 20134
rect 198986 -1502 199222 -1266
rect 198986 -1822 199222 -1586
rect 202586 671818 202822 672054
rect 202586 671498 202822 671734
rect 202586 635818 202822 636054
rect 202586 635498 202822 635734
rect 202586 599818 202822 600054
rect 202586 599498 202822 599734
rect 202586 563818 202822 564054
rect 202586 563498 202822 563734
rect 206186 675418 206422 675654
rect 206186 675098 206422 675334
rect 206186 639418 206422 639654
rect 206186 639098 206422 639334
rect 206186 603418 206422 603654
rect 206186 603098 206422 603334
rect 206186 567418 206422 567654
rect 206186 567098 206422 567334
rect 204950 562732 205186 562818
rect 204950 562668 205036 562732
rect 205036 562668 205100 562732
rect 205100 562668 205186 562732
rect 204950 562582 205186 562668
rect 202586 527818 202822 528054
rect 202586 527498 202822 527734
rect 202586 491818 202822 492054
rect 202586 491498 202822 491734
rect 202586 455818 202822 456054
rect 202586 455498 202822 455734
rect 202586 419818 202822 420054
rect 202586 419498 202822 419734
rect 202586 383818 202822 384054
rect 202586 383498 202822 383734
rect 202586 347818 202822 348054
rect 202586 347498 202822 347734
rect 202586 311818 202822 312054
rect 202586 311498 202822 311734
rect 202586 275818 202822 276054
rect 202586 275498 202822 275734
rect 202586 239818 202822 240054
rect 202586 239498 202822 239734
rect 202586 203818 202822 204054
rect 202586 203498 202822 203734
rect 202586 167818 202822 168054
rect 202586 167498 202822 167734
rect 202586 131818 202822 132054
rect 202586 131498 202822 131734
rect 202586 95818 202822 96054
rect 202586 95498 202822 95734
rect 202586 59818 202822 60054
rect 202586 59498 202822 59734
rect 202586 23818 202822 24054
rect 202586 23498 202822 23734
rect 202586 -3342 202822 -3106
rect 202586 -3662 202822 -3426
rect 227786 710122 228022 710358
rect 227786 709802 228022 710038
rect 224186 708282 224422 708518
rect 224186 707962 224422 708198
rect 220586 706442 220822 706678
rect 220586 706122 220822 706358
rect 209786 679018 210022 679254
rect 209786 678698 210022 678934
rect 209786 643018 210022 643254
rect 209786 642698 210022 642934
rect 209786 607018 210022 607254
rect 209786 606698 210022 606934
rect 209786 571018 210022 571254
rect 209786 570698 210022 570934
rect 207526 561222 207762 561458
rect 206186 531418 206422 531654
rect 206186 531098 206422 531334
rect 206186 495418 206422 495654
rect 206186 495098 206422 495334
rect 206186 459418 206422 459654
rect 206186 459098 206422 459334
rect 206186 423418 206422 423654
rect 206186 423098 206422 423334
rect 206186 387418 206422 387654
rect 206186 387098 206422 387334
rect 206186 351418 206422 351654
rect 206186 351098 206422 351334
rect 206186 315418 206422 315654
rect 206186 315098 206422 315334
rect 206186 279418 206422 279654
rect 206186 279098 206422 279334
rect 206186 243418 206422 243654
rect 206186 243098 206422 243334
rect 206186 207418 206422 207654
rect 206186 207098 206422 207334
rect 206186 171418 206422 171654
rect 206186 171098 206422 171334
rect 206186 135418 206422 135654
rect 206186 135098 206422 135334
rect 206186 99418 206422 99654
rect 206186 99098 206422 99334
rect 206186 63418 206422 63654
rect 206186 63098 206422 63334
rect 206186 27418 206422 27654
rect 206186 27098 206422 27334
rect 206186 -5182 206422 -4946
rect 206186 -5502 206422 -5266
rect 209786 535018 210022 535254
rect 209786 534698 210022 534934
rect 209786 499018 210022 499254
rect 209786 498698 210022 498934
rect 209786 463018 210022 463254
rect 209786 462698 210022 462934
rect 209786 427018 210022 427254
rect 209786 426698 210022 426934
rect 209786 391018 210022 391254
rect 209786 390698 210022 390934
rect 209786 355018 210022 355254
rect 209786 354698 210022 354934
rect 209786 319018 210022 319254
rect 209786 318698 210022 318934
rect 209786 283018 210022 283254
rect 209786 282698 210022 282934
rect 209786 247018 210022 247254
rect 209786 246698 210022 246934
rect 209786 211018 210022 211254
rect 209786 210698 210022 210934
rect 209786 175018 210022 175254
rect 209786 174698 210022 174934
rect 209786 139018 210022 139254
rect 209786 138698 210022 138934
rect 209786 103018 210022 103254
rect 209786 102698 210022 102934
rect 209786 67018 210022 67254
rect 209786 66698 210022 66934
rect 209786 31018 210022 31254
rect 209786 30698 210022 30934
rect 191786 -6102 192022 -5866
rect 191786 -6422 192022 -6186
rect 216986 704602 217222 704838
rect 216986 704282 217222 704518
rect 216986 686218 217222 686454
rect 216986 685898 217222 686134
rect 216986 650218 217222 650454
rect 216986 649898 217222 650134
rect 216986 614218 217222 614454
rect 216986 613898 217222 614134
rect 216986 578218 217222 578454
rect 216986 577898 217222 578134
rect 216986 542218 217222 542454
rect 216986 541898 217222 542134
rect 216986 506218 217222 506454
rect 216986 505898 217222 506134
rect 216986 470218 217222 470454
rect 216986 469898 217222 470134
rect 216986 434218 217222 434454
rect 216986 433898 217222 434134
rect 216986 398218 217222 398454
rect 216986 397898 217222 398134
rect 216986 362218 217222 362454
rect 216986 361898 217222 362134
rect 216986 326218 217222 326454
rect 216986 325898 217222 326134
rect 216986 290218 217222 290454
rect 216986 289898 217222 290134
rect 216986 254218 217222 254454
rect 216986 253898 217222 254134
rect 216986 218218 217222 218454
rect 216986 217898 217222 218134
rect 216986 182218 217222 182454
rect 216986 181898 217222 182134
rect 216986 146218 217222 146454
rect 216986 145898 217222 146134
rect 216986 110218 217222 110454
rect 216986 109898 217222 110134
rect 216986 74218 217222 74454
rect 216986 73898 217222 74134
rect 216986 38218 217222 38454
rect 216986 37898 217222 38134
rect 216986 2218 217222 2454
rect 216986 1898 217222 2134
rect 216986 -582 217222 -346
rect 216986 -902 217222 -666
rect 220586 689818 220822 690054
rect 220586 689498 220822 689734
rect 220586 653818 220822 654054
rect 220586 653498 220822 653734
rect 220586 617818 220822 618054
rect 220586 617498 220822 617734
rect 220586 581818 220822 582054
rect 220586 581498 220822 581734
rect 224186 693418 224422 693654
rect 224186 693098 224422 693334
rect 224186 657418 224422 657654
rect 224186 657098 224422 657334
rect 224186 621418 224422 621654
rect 224186 621098 224422 621334
rect 224186 585418 224422 585654
rect 224186 585098 224422 585334
rect 223534 561372 223770 561458
rect 223534 561308 223620 561372
rect 223620 561308 223684 561372
rect 223684 561308 223770 561372
rect 223534 561222 223770 561308
rect 220586 545818 220822 546054
rect 220586 545498 220822 545734
rect 220586 509818 220822 510054
rect 220586 509498 220822 509734
rect 220586 473818 220822 474054
rect 220586 473498 220822 473734
rect 220586 437818 220822 438054
rect 220586 437498 220822 437734
rect 220586 401818 220822 402054
rect 220586 401498 220822 401734
rect 220586 365818 220822 366054
rect 220586 365498 220822 365734
rect 220586 329818 220822 330054
rect 220586 329498 220822 329734
rect 220586 293818 220822 294054
rect 220586 293498 220822 293734
rect 220586 257818 220822 258054
rect 220586 257498 220822 257734
rect 220586 221818 220822 222054
rect 220586 221498 220822 221734
rect 220586 185818 220822 186054
rect 220586 185498 220822 185734
rect 220586 149818 220822 150054
rect 220586 149498 220822 149734
rect 220586 113818 220822 114054
rect 220586 113498 220822 113734
rect 220586 77818 220822 78054
rect 220586 77498 220822 77734
rect 220586 41818 220822 42054
rect 220586 41498 220822 41734
rect 220586 5818 220822 6054
rect 220586 5498 220822 5734
rect 220586 -2422 220822 -2186
rect 220586 -2742 220822 -2506
rect 245786 711042 246022 711278
rect 245786 710722 246022 710958
rect 242186 709202 242422 709438
rect 242186 708882 242422 709118
rect 238586 707362 238822 707598
rect 238586 707042 238822 707278
rect 227786 697018 228022 697254
rect 227786 696698 228022 696934
rect 227786 661018 228022 661254
rect 227786 660698 228022 660934
rect 227786 625018 228022 625254
rect 227786 624698 228022 624934
rect 227786 589018 228022 589254
rect 227786 588698 228022 588934
rect 225374 561902 225610 562138
rect 224186 549418 224422 549654
rect 224186 549098 224422 549334
rect 224186 513418 224422 513654
rect 224186 513098 224422 513334
rect 224186 477418 224422 477654
rect 224186 477098 224422 477334
rect 224186 441418 224422 441654
rect 224186 441098 224422 441334
rect 224186 405418 224422 405654
rect 224186 405098 224422 405334
rect 224186 369418 224422 369654
rect 224186 369098 224422 369334
rect 224186 333418 224422 333654
rect 224186 333098 224422 333334
rect 224186 297418 224422 297654
rect 224186 297098 224422 297334
rect 224186 261418 224422 261654
rect 224186 261098 224422 261334
rect 224186 225418 224422 225654
rect 224186 225098 224422 225334
rect 224186 189418 224422 189654
rect 224186 189098 224422 189334
rect 224186 153418 224422 153654
rect 224186 153098 224422 153334
rect 224186 117418 224422 117654
rect 224186 117098 224422 117334
rect 224186 81418 224422 81654
rect 224186 81098 224422 81334
rect 224186 45418 224422 45654
rect 224186 45098 224422 45334
rect 224186 9418 224422 9654
rect 224186 9098 224422 9334
rect 224186 -4262 224422 -4026
rect 224186 -4582 224422 -4346
rect 234986 705522 235222 705758
rect 234986 705202 235222 705438
rect 234986 668218 235222 668454
rect 234986 667898 235222 668134
rect 234986 632218 235222 632454
rect 234986 631898 235222 632134
rect 234986 596218 235222 596454
rect 234986 595898 235222 596134
rect 238586 671818 238822 672054
rect 238586 671498 238822 671734
rect 238586 635818 238822 636054
rect 238586 635498 238822 635734
rect 238586 599818 238822 600054
rect 238586 599498 238822 599734
rect 238586 563818 238822 564054
rect 238586 563498 238822 563734
rect 234986 560218 235222 560454
rect 234986 559898 235222 560134
rect 227786 553018 228022 553254
rect 227786 552698 228022 552934
rect 227786 517018 228022 517254
rect 227786 516698 228022 516934
rect 227786 481018 228022 481254
rect 227786 480698 228022 480934
rect 227786 445018 228022 445254
rect 227786 444698 228022 444934
rect 227786 409018 228022 409254
rect 227786 408698 228022 408934
rect 227786 373018 228022 373254
rect 227786 372698 228022 372934
rect 227786 337018 228022 337254
rect 227786 336698 228022 336934
rect 227786 301018 228022 301254
rect 227786 300698 228022 300934
rect 227786 265018 228022 265254
rect 227786 264698 228022 264934
rect 227786 229018 228022 229254
rect 227786 228698 228022 228934
rect 227786 193018 228022 193254
rect 227786 192698 228022 192934
rect 227786 157018 228022 157254
rect 227786 156698 228022 156934
rect 227786 121018 228022 121254
rect 227786 120698 228022 120934
rect 227786 85018 228022 85254
rect 227786 84698 228022 84934
rect 227786 49018 228022 49254
rect 227786 48698 228022 48934
rect 234986 524218 235222 524454
rect 234986 523898 235222 524134
rect 234986 488218 235222 488454
rect 234986 487898 235222 488134
rect 234986 452218 235222 452454
rect 234986 451898 235222 452134
rect 234986 416218 235222 416454
rect 234986 415898 235222 416134
rect 234986 380218 235222 380454
rect 234986 379898 235222 380134
rect 234986 344218 235222 344454
rect 234986 343898 235222 344134
rect 234986 308218 235222 308454
rect 234986 307898 235222 308134
rect 234986 272218 235222 272454
rect 234986 271898 235222 272134
rect 234986 236218 235222 236454
rect 234986 235898 235222 236134
rect 234986 200218 235222 200454
rect 234986 199898 235222 200134
rect 234986 164218 235222 164454
rect 234986 163898 235222 164134
rect 234986 128218 235222 128454
rect 234986 127898 235222 128134
rect 234986 92218 235222 92454
rect 234986 91898 235222 92134
rect 238586 527818 238822 528054
rect 238586 527498 238822 527734
rect 238586 491818 238822 492054
rect 238586 491498 238822 491734
rect 238586 455818 238822 456054
rect 238586 455498 238822 455734
rect 238586 419818 238822 420054
rect 238586 419498 238822 419734
rect 238586 383818 238822 384054
rect 238586 383498 238822 383734
rect 238586 347818 238822 348054
rect 238586 347498 238822 347734
rect 238586 311818 238822 312054
rect 238586 311498 238822 311734
rect 238586 275818 238822 276054
rect 238586 275498 238822 275734
rect 238586 239818 238822 240054
rect 238586 239498 238822 239734
rect 238586 203818 238822 204054
rect 238586 203498 238822 203734
rect 242186 675418 242422 675654
rect 242186 675098 242422 675334
rect 242186 639418 242422 639654
rect 242186 639098 242422 639334
rect 242186 603418 242422 603654
rect 242186 603098 242422 603334
rect 242186 567418 242422 567654
rect 242186 567098 242422 567334
rect 263786 710122 264022 710358
rect 263786 709802 264022 710038
rect 260186 708282 260422 708518
rect 260186 707962 260422 708198
rect 256586 706442 256822 706678
rect 256586 706122 256822 706358
rect 245786 679018 246022 679254
rect 245786 678698 246022 678934
rect 245786 643018 246022 643254
rect 245786 642698 246022 642934
rect 245786 607018 246022 607254
rect 245786 606698 246022 606934
rect 245786 571018 246022 571254
rect 245786 570698 246022 570934
rect 242186 531418 242422 531654
rect 242186 531098 242422 531334
rect 242186 495418 242422 495654
rect 242186 495098 242422 495334
rect 242186 459418 242422 459654
rect 242186 459098 242422 459334
rect 242186 423418 242422 423654
rect 242186 423098 242422 423334
rect 242186 387418 242422 387654
rect 242186 387098 242422 387334
rect 242186 351418 242422 351654
rect 242186 351098 242422 351334
rect 242186 315418 242422 315654
rect 242186 315098 242422 315334
rect 242186 279418 242422 279654
rect 242186 279098 242422 279334
rect 242186 243418 242422 243654
rect 242186 243098 242422 243334
rect 242186 207418 242422 207654
rect 242186 207098 242422 207334
rect 238586 167818 238822 168054
rect 238586 167498 238822 167734
rect 238586 131818 238822 132054
rect 238586 131498 238822 131734
rect 238586 95818 238822 96054
rect 238586 95498 238822 95734
rect 234986 56218 235222 56454
rect 234986 55898 235222 56134
rect 234986 20218 235222 20454
rect 234986 19898 235222 20134
rect 227786 13018 228022 13254
rect 227786 12698 228022 12934
rect 209786 -7022 210022 -6786
rect 209786 -7342 210022 -7106
rect 234986 -1502 235222 -1266
rect 234986 -1822 235222 -1586
rect 238586 59818 238822 60054
rect 238586 59498 238822 59734
rect 238586 23818 238822 24054
rect 238586 23498 238822 23734
rect 238586 -3342 238822 -3106
rect 238586 -3662 238822 -3426
rect 242186 171418 242422 171654
rect 242186 171098 242422 171334
rect 242186 135418 242422 135654
rect 242186 135098 242422 135334
rect 242186 99418 242422 99654
rect 242186 99098 242422 99334
rect 242186 63418 242422 63654
rect 242186 63098 242422 63334
rect 242186 27418 242422 27654
rect 242186 27098 242422 27334
rect 242186 -5182 242422 -4946
rect 242186 -5502 242422 -5266
rect 252986 704602 253222 704838
rect 252986 704282 253222 704518
rect 252986 686218 253222 686454
rect 252986 685898 253222 686134
rect 252986 650218 253222 650454
rect 252986 649898 253222 650134
rect 252986 614218 253222 614454
rect 252986 613898 253222 614134
rect 252986 578218 253222 578454
rect 252986 577898 253222 578134
rect 252422 561902 252658 562138
rect 245786 535018 246022 535254
rect 245786 534698 246022 534934
rect 245786 499018 246022 499254
rect 245786 498698 246022 498934
rect 245786 463018 246022 463254
rect 245786 462698 246022 462934
rect 245786 427018 246022 427254
rect 245786 426698 246022 426934
rect 245786 391018 246022 391254
rect 245786 390698 246022 390934
rect 245786 355018 246022 355254
rect 245786 354698 246022 354934
rect 245786 319018 246022 319254
rect 245786 318698 246022 318934
rect 245786 283018 246022 283254
rect 245786 282698 246022 282934
rect 245786 247018 246022 247254
rect 245786 246698 246022 246934
rect 245786 211018 246022 211254
rect 245786 210698 246022 210934
rect 245786 175018 246022 175254
rect 245786 174698 246022 174934
rect 245786 139018 246022 139254
rect 245786 138698 246022 138934
rect 245786 103018 246022 103254
rect 245786 102698 246022 102934
rect 245786 67018 246022 67254
rect 245786 66698 246022 66934
rect 256586 689818 256822 690054
rect 256586 689498 256822 689734
rect 256586 653818 256822 654054
rect 256586 653498 256822 653734
rect 256586 617818 256822 618054
rect 256586 617498 256822 617734
rect 256586 581818 256822 582054
rect 256586 581498 256822 581734
rect 253526 562582 253762 562818
rect 252986 542218 253222 542454
rect 252986 541898 253222 542134
rect 252986 506218 253222 506454
rect 252986 505898 253222 506134
rect 252986 470218 253222 470454
rect 252986 469898 253222 470134
rect 252986 434218 253222 434454
rect 252986 433898 253222 434134
rect 252986 398218 253222 398454
rect 252986 397898 253222 398134
rect 252986 362218 253222 362454
rect 252986 361898 253222 362134
rect 252986 326218 253222 326454
rect 252986 325898 253222 326134
rect 252986 290218 253222 290454
rect 252986 289898 253222 290134
rect 252986 254218 253222 254454
rect 252986 253898 253222 254134
rect 252986 218218 253222 218454
rect 252986 217898 253222 218134
rect 252986 182218 253222 182454
rect 252986 181898 253222 182134
rect 252986 146218 253222 146454
rect 252986 145898 253222 146134
rect 252986 110218 253222 110454
rect 252986 109898 253222 110134
rect 252986 74218 253222 74454
rect 252986 73898 253222 74134
rect 245786 31018 246022 31254
rect 245786 30698 246022 30934
rect 227786 -6102 228022 -5866
rect 227786 -6422 228022 -6186
rect 252986 38218 253222 38454
rect 252986 37898 253222 38134
rect 252986 2218 253222 2454
rect 252986 1898 253222 2134
rect 252986 -582 253222 -346
rect 252986 -902 253222 -666
rect 256586 545818 256822 546054
rect 256586 545498 256822 545734
rect 256586 509818 256822 510054
rect 256586 509498 256822 509734
rect 256586 473818 256822 474054
rect 256586 473498 256822 473734
rect 256586 437818 256822 438054
rect 256586 437498 256822 437734
rect 256586 401818 256822 402054
rect 256586 401498 256822 401734
rect 256586 365818 256822 366054
rect 256586 365498 256822 365734
rect 256586 329818 256822 330054
rect 256586 329498 256822 329734
rect 256586 293818 256822 294054
rect 256586 293498 256822 293734
rect 256586 257818 256822 258054
rect 256586 257498 256822 257734
rect 256586 221818 256822 222054
rect 256586 221498 256822 221734
rect 256586 185818 256822 186054
rect 256586 185498 256822 185734
rect 256586 149818 256822 150054
rect 256586 149498 256822 149734
rect 256586 113818 256822 114054
rect 256586 113498 256822 113734
rect 256586 77818 256822 78054
rect 256586 77498 256822 77734
rect 256586 41818 256822 42054
rect 256586 41498 256822 41734
rect 256586 5818 256822 6054
rect 256586 5498 256822 5734
rect 256586 -2422 256822 -2186
rect 256586 -2742 256822 -2506
rect 260186 693418 260422 693654
rect 260186 693098 260422 693334
rect 260186 657418 260422 657654
rect 260186 657098 260422 657334
rect 260186 621418 260422 621654
rect 260186 621098 260422 621334
rect 260186 585418 260422 585654
rect 260186 585098 260422 585334
rect 260186 549418 260422 549654
rect 260186 549098 260422 549334
rect 260186 513418 260422 513654
rect 260186 513098 260422 513334
rect 260186 477418 260422 477654
rect 260186 477098 260422 477334
rect 260186 441418 260422 441654
rect 260186 441098 260422 441334
rect 260186 405418 260422 405654
rect 260186 405098 260422 405334
rect 260186 369418 260422 369654
rect 260186 369098 260422 369334
rect 260186 333418 260422 333654
rect 260186 333098 260422 333334
rect 260186 297418 260422 297654
rect 260186 297098 260422 297334
rect 260186 261418 260422 261654
rect 260186 261098 260422 261334
rect 260186 225418 260422 225654
rect 260186 225098 260422 225334
rect 260186 189418 260422 189654
rect 260186 189098 260422 189334
rect 260186 153418 260422 153654
rect 260186 153098 260422 153334
rect 260186 117418 260422 117654
rect 260186 117098 260422 117334
rect 260186 81418 260422 81654
rect 260186 81098 260422 81334
rect 260186 45418 260422 45654
rect 260186 45098 260422 45334
rect 260186 9418 260422 9654
rect 260186 9098 260422 9334
rect 260186 -4262 260422 -4026
rect 260186 -4582 260422 -4346
rect 281786 711042 282022 711278
rect 281786 710722 282022 710958
rect 278186 709202 278422 709438
rect 278186 708882 278422 709118
rect 274586 707362 274822 707598
rect 274586 707042 274822 707278
rect 263786 697018 264022 697254
rect 263786 696698 264022 696934
rect 263786 661018 264022 661254
rect 263786 660698 264022 660934
rect 263786 625018 264022 625254
rect 263786 624698 264022 624934
rect 263786 589018 264022 589254
rect 263786 588698 264022 588934
rect 270986 705522 271222 705758
rect 270986 705202 271222 705438
rect 270986 668218 271222 668454
rect 270986 667898 271222 668134
rect 270986 632218 271222 632454
rect 270986 631898 271222 632134
rect 270986 596218 271222 596454
rect 270986 595898 271222 596134
rect 266222 561902 266458 562138
rect 263786 553018 264022 553254
rect 263786 552698 264022 552934
rect 263786 517018 264022 517254
rect 263786 516698 264022 516934
rect 263786 481018 264022 481254
rect 263786 480698 264022 480934
rect 263786 445018 264022 445254
rect 263786 444698 264022 444934
rect 263786 409018 264022 409254
rect 263786 408698 264022 408934
rect 263786 373018 264022 373254
rect 263786 372698 264022 372934
rect 263786 337018 264022 337254
rect 263786 336698 264022 336934
rect 263786 301018 264022 301254
rect 263786 300698 264022 300934
rect 263786 265018 264022 265254
rect 263786 264698 264022 264934
rect 263786 229018 264022 229254
rect 263786 228698 264022 228934
rect 263786 193018 264022 193254
rect 263786 192698 264022 192934
rect 263786 157018 264022 157254
rect 263786 156698 264022 156934
rect 263786 121018 264022 121254
rect 263786 120698 264022 120934
rect 270986 560218 271222 560454
rect 270986 559898 271222 560134
rect 270986 524218 271222 524454
rect 270986 523898 271222 524134
rect 270986 488218 271222 488454
rect 270986 487898 271222 488134
rect 270986 452218 271222 452454
rect 270986 451898 271222 452134
rect 270986 416218 271222 416454
rect 270986 415898 271222 416134
rect 270986 380218 271222 380454
rect 270986 379898 271222 380134
rect 270986 344218 271222 344454
rect 270986 343898 271222 344134
rect 270986 308218 271222 308454
rect 270986 307898 271222 308134
rect 270986 272218 271222 272454
rect 270986 271898 271222 272134
rect 270986 236218 271222 236454
rect 270986 235898 271222 236134
rect 270986 200218 271222 200454
rect 270986 199898 271222 200134
rect 270986 164218 271222 164454
rect 270986 163898 271222 164134
rect 270986 128218 271222 128454
rect 270986 127898 271222 128134
rect 270986 92218 271222 92454
rect 270986 91898 271222 92134
rect 263786 85018 264022 85254
rect 263786 84698 264022 84934
rect 263786 49018 264022 49254
rect 263786 48698 264022 48934
rect 263786 13018 264022 13254
rect 263786 12698 264022 12934
rect 245786 -7022 246022 -6786
rect 245786 -7342 246022 -7106
rect 270986 56218 271222 56454
rect 270986 55898 271222 56134
rect 270986 20218 271222 20454
rect 270986 19898 271222 20134
rect 270986 -1502 271222 -1266
rect 270986 -1822 271222 -1586
rect 274586 671818 274822 672054
rect 274586 671498 274822 671734
rect 274586 635818 274822 636054
rect 274586 635498 274822 635734
rect 274586 599818 274822 600054
rect 274586 599498 274822 599734
rect 274586 563818 274822 564054
rect 274586 563498 274822 563734
rect 278186 675418 278422 675654
rect 278186 675098 278422 675334
rect 278186 639418 278422 639654
rect 278186 639098 278422 639334
rect 278186 603418 278422 603654
rect 278186 603098 278422 603334
rect 278186 567418 278422 567654
rect 278186 567098 278422 567334
rect 275790 562582 276026 562818
rect 274586 527818 274822 528054
rect 274586 527498 274822 527734
rect 274586 491818 274822 492054
rect 274586 491498 274822 491734
rect 274586 455818 274822 456054
rect 274586 455498 274822 455734
rect 274586 419818 274822 420054
rect 274586 419498 274822 419734
rect 274586 383818 274822 384054
rect 274586 383498 274822 383734
rect 274586 347818 274822 348054
rect 274586 347498 274822 347734
rect 274586 311818 274822 312054
rect 274586 311498 274822 311734
rect 274586 275818 274822 276054
rect 274586 275498 274822 275734
rect 274586 239818 274822 240054
rect 274586 239498 274822 239734
rect 274586 203818 274822 204054
rect 274586 203498 274822 203734
rect 274586 167818 274822 168054
rect 274586 167498 274822 167734
rect 274586 131818 274822 132054
rect 274586 131498 274822 131734
rect 274586 95818 274822 96054
rect 274586 95498 274822 95734
rect 274586 59818 274822 60054
rect 274586 59498 274822 59734
rect 274586 23818 274822 24054
rect 274586 23498 274822 23734
rect 274586 -3342 274822 -3106
rect 274586 -3662 274822 -3426
rect 299786 710122 300022 710358
rect 299786 709802 300022 710038
rect 296186 708282 296422 708518
rect 296186 707962 296422 708198
rect 292586 706442 292822 706678
rect 292586 706122 292822 706358
rect 281786 679018 282022 679254
rect 281786 678698 282022 678934
rect 281786 643018 282022 643254
rect 281786 642698 282022 642934
rect 281786 607018 282022 607254
rect 281786 606698 282022 606934
rect 281786 571018 282022 571254
rect 281786 570698 282022 570934
rect 278186 531418 278422 531654
rect 278186 531098 278422 531334
rect 278186 495418 278422 495654
rect 278186 495098 278422 495334
rect 278186 459418 278422 459654
rect 278186 459098 278422 459334
rect 278186 423418 278422 423654
rect 278186 423098 278422 423334
rect 278186 387418 278422 387654
rect 278186 387098 278422 387334
rect 278186 351418 278422 351654
rect 278186 351098 278422 351334
rect 278186 315418 278422 315654
rect 278186 315098 278422 315334
rect 278186 279418 278422 279654
rect 278186 279098 278422 279334
rect 278186 243418 278422 243654
rect 278186 243098 278422 243334
rect 278186 207418 278422 207654
rect 278186 207098 278422 207334
rect 278186 171418 278422 171654
rect 278186 171098 278422 171334
rect 278186 135418 278422 135654
rect 278186 135098 278422 135334
rect 278186 99418 278422 99654
rect 278186 99098 278422 99334
rect 278186 63418 278422 63654
rect 278186 63098 278422 63334
rect 278186 27418 278422 27654
rect 278186 27098 278422 27334
rect 278186 -5182 278422 -4946
rect 278186 -5502 278422 -5266
rect 288986 704602 289222 704838
rect 288986 704282 289222 704518
rect 288986 686218 289222 686454
rect 288986 685898 289222 686134
rect 288986 650218 289222 650454
rect 288986 649898 289222 650134
rect 288986 614218 289222 614454
rect 288986 613898 289222 614134
rect 288986 578218 289222 578454
rect 288986 577898 289222 578134
rect 288302 561902 288538 562138
rect 281786 535018 282022 535254
rect 281786 534698 282022 534934
rect 281786 499018 282022 499254
rect 281786 498698 282022 498934
rect 281786 463018 282022 463254
rect 281786 462698 282022 462934
rect 281786 427018 282022 427254
rect 281786 426698 282022 426934
rect 281786 391018 282022 391254
rect 281786 390698 282022 390934
rect 281786 355018 282022 355254
rect 281786 354698 282022 354934
rect 281786 319018 282022 319254
rect 281786 318698 282022 318934
rect 281786 283018 282022 283254
rect 281786 282698 282022 282934
rect 281786 247018 282022 247254
rect 281786 246698 282022 246934
rect 281786 211018 282022 211254
rect 281786 210698 282022 210934
rect 281786 175018 282022 175254
rect 281786 174698 282022 174934
rect 281786 139018 282022 139254
rect 281786 138698 282022 138934
rect 281786 103018 282022 103254
rect 281786 102698 282022 102934
rect 281786 67018 282022 67254
rect 281786 66698 282022 66934
rect 281786 31018 282022 31254
rect 281786 30698 282022 30934
rect 263786 -6102 264022 -5866
rect 263786 -6422 264022 -6186
rect 288986 542218 289222 542454
rect 288986 541898 289222 542134
rect 288986 506218 289222 506454
rect 288986 505898 289222 506134
rect 288986 470218 289222 470454
rect 288986 469898 289222 470134
rect 288986 434218 289222 434454
rect 288986 433898 289222 434134
rect 288986 398218 289222 398454
rect 288986 397898 289222 398134
rect 288986 362218 289222 362454
rect 288986 361898 289222 362134
rect 288986 326218 289222 326454
rect 288986 325898 289222 326134
rect 288986 290218 289222 290454
rect 288986 289898 289222 290134
rect 288986 254218 289222 254454
rect 288986 253898 289222 254134
rect 288986 218218 289222 218454
rect 288986 217898 289222 218134
rect 288986 182218 289222 182454
rect 288986 181898 289222 182134
rect 288986 146218 289222 146454
rect 288986 145898 289222 146134
rect 288986 110218 289222 110454
rect 288986 109898 289222 110134
rect 288986 74218 289222 74454
rect 288986 73898 289222 74134
rect 288986 38218 289222 38454
rect 288986 37898 289222 38134
rect 288986 2218 289222 2454
rect 288986 1898 289222 2134
rect 288986 -582 289222 -346
rect 288986 -902 289222 -666
rect 292586 689818 292822 690054
rect 292586 689498 292822 689734
rect 292586 653818 292822 654054
rect 292586 653498 292822 653734
rect 292586 617818 292822 618054
rect 292586 617498 292822 617734
rect 292586 581818 292822 582054
rect 292586 581498 292822 581734
rect 296186 693418 296422 693654
rect 296186 693098 296422 693334
rect 296186 657418 296422 657654
rect 296186 657098 296422 657334
rect 296186 621418 296422 621654
rect 296186 621098 296422 621334
rect 296186 585418 296422 585654
rect 296186 585098 296422 585334
rect 293086 562582 293322 562818
rect 292586 545818 292822 546054
rect 292586 545498 292822 545734
rect 292586 509818 292822 510054
rect 292586 509498 292822 509734
rect 292586 473818 292822 474054
rect 292586 473498 292822 473734
rect 292586 437818 292822 438054
rect 292586 437498 292822 437734
rect 292586 401818 292822 402054
rect 292586 401498 292822 401734
rect 292586 365818 292822 366054
rect 292586 365498 292822 365734
rect 292586 329818 292822 330054
rect 292586 329498 292822 329734
rect 292586 293818 292822 294054
rect 292586 293498 292822 293734
rect 292586 257818 292822 258054
rect 292586 257498 292822 257734
rect 292586 221818 292822 222054
rect 292586 221498 292822 221734
rect 292586 185818 292822 186054
rect 292586 185498 292822 185734
rect 292586 149818 292822 150054
rect 292586 149498 292822 149734
rect 292586 113818 292822 114054
rect 292586 113498 292822 113734
rect 292586 77818 292822 78054
rect 292586 77498 292822 77734
rect 292586 41818 292822 42054
rect 292586 41498 292822 41734
rect 292586 5818 292822 6054
rect 292586 5498 292822 5734
rect 292586 -2422 292822 -2186
rect 292586 -2742 292822 -2506
rect 317786 711042 318022 711278
rect 317786 710722 318022 710958
rect 314186 709202 314422 709438
rect 314186 708882 314422 709118
rect 310586 707362 310822 707598
rect 310586 707042 310822 707278
rect 299786 697018 300022 697254
rect 299786 696698 300022 696934
rect 299786 661018 300022 661254
rect 299786 660698 300022 660934
rect 299786 625018 300022 625254
rect 299786 624698 300022 624934
rect 299786 589018 300022 589254
rect 299786 588698 300022 588934
rect 296186 549418 296422 549654
rect 296186 549098 296422 549334
rect 296186 513418 296422 513654
rect 296186 513098 296422 513334
rect 296186 477418 296422 477654
rect 296186 477098 296422 477334
rect 296186 441418 296422 441654
rect 296186 441098 296422 441334
rect 296186 405418 296422 405654
rect 296186 405098 296422 405334
rect 296186 369418 296422 369654
rect 296186 369098 296422 369334
rect 296186 333418 296422 333654
rect 296186 333098 296422 333334
rect 296186 297418 296422 297654
rect 296186 297098 296422 297334
rect 296186 261418 296422 261654
rect 296186 261098 296422 261334
rect 296186 225418 296422 225654
rect 296186 225098 296422 225334
rect 296186 189418 296422 189654
rect 296186 189098 296422 189334
rect 299786 553018 300022 553254
rect 299786 552698 300022 552934
rect 299786 517018 300022 517254
rect 299786 516698 300022 516934
rect 299786 481018 300022 481254
rect 299786 480698 300022 480934
rect 299786 445018 300022 445254
rect 299786 444698 300022 444934
rect 299786 409018 300022 409254
rect 299786 408698 300022 408934
rect 299786 373018 300022 373254
rect 299786 372698 300022 372934
rect 299786 337018 300022 337254
rect 299786 336698 300022 336934
rect 299786 301018 300022 301254
rect 299786 300698 300022 300934
rect 299786 265018 300022 265254
rect 299786 264698 300022 264934
rect 299786 229018 300022 229254
rect 299786 228698 300022 228934
rect 299786 193018 300022 193254
rect 299786 192698 300022 192934
rect 296186 153418 296422 153654
rect 296186 153098 296422 153334
rect 296186 117418 296422 117654
rect 296186 117098 296422 117334
rect 299786 157018 300022 157254
rect 299786 156698 300022 156934
rect 299786 121018 300022 121254
rect 299786 120698 300022 120934
rect 296186 81418 296422 81654
rect 296186 81098 296422 81334
rect 296186 45418 296422 45654
rect 296186 45098 296422 45334
rect 296186 9418 296422 9654
rect 296186 9098 296422 9334
rect 296186 -4262 296422 -4026
rect 296186 -4582 296422 -4346
rect 299786 85018 300022 85254
rect 299786 84698 300022 84934
rect 299786 49018 300022 49254
rect 299786 48698 300022 48934
rect 299786 13018 300022 13254
rect 299786 12698 300022 12934
rect 281786 -7022 282022 -6786
rect 281786 -7342 282022 -7106
rect 306986 705522 307222 705758
rect 306986 705202 307222 705438
rect 306986 668218 307222 668454
rect 306986 667898 307222 668134
rect 306986 632218 307222 632454
rect 306986 631898 307222 632134
rect 306986 596218 307222 596454
rect 306986 595898 307222 596134
rect 310586 671818 310822 672054
rect 310586 671498 310822 671734
rect 310586 635818 310822 636054
rect 310586 635498 310822 635734
rect 310586 599818 310822 600054
rect 310586 599498 310822 599734
rect 310586 563818 310822 564054
rect 310586 563498 310822 563734
rect 306986 560218 307222 560454
rect 306986 559898 307222 560134
rect 306986 524218 307222 524454
rect 306986 523898 307222 524134
rect 306986 488218 307222 488454
rect 306986 487898 307222 488134
rect 306986 452218 307222 452454
rect 306986 451898 307222 452134
rect 306986 416218 307222 416454
rect 306986 415898 307222 416134
rect 306986 380218 307222 380454
rect 306986 379898 307222 380134
rect 306986 344218 307222 344454
rect 306986 343898 307222 344134
rect 306986 308218 307222 308454
rect 306986 307898 307222 308134
rect 306986 272218 307222 272454
rect 306986 271898 307222 272134
rect 306986 236218 307222 236454
rect 306986 235898 307222 236134
rect 306986 200218 307222 200454
rect 306986 199898 307222 200134
rect 306986 164218 307222 164454
rect 306986 163898 307222 164134
rect 306986 128218 307222 128454
rect 306986 127898 307222 128134
rect 306986 92218 307222 92454
rect 306986 91898 307222 92134
rect 306986 56218 307222 56454
rect 306986 55898 307222 56134
rect 306986 20218 307222 20454
rect 306986 19898 307222 20134
rect 306986 -1502 307222 -1266
rect 306986 -1822 307222 -1586
rect 314186 675418 314422 675654
rect 314186 675098 314422 675334
rect 314186 639418 314422 639654
rect 314186 639098 314422 639334
rect 314186 603418 314422 603654
rect 314186 603098 314422 603334
rect 314186 567418 314422 567654
rect 314186 567098 314422 567334
rect 310586 527818 310822 528054
rect 310586 527498 310822 527734
rect 310586 491818 310822 492054
rect 310586 491498 310822 491734
rect 310586 455818 310822 456054
rect 310586 455498 310822 455734
rect 310586 419818 310822 420054
rect 310586 419498 310822 419734
rect 310586 383818 310822 384054
rect 310586 383498 310822 383734
rect 310586 347818 310822 348054
rect 310586 347498 310822 347734
rect 310586 311818 310822 312054
rect 310586 311498 310822 311734
rect 310586 275818 310822 276054
rect 310586 275498 310822 275734
rect 310586 239818 310822 240054
rect 310586 239498 310822 239734
rect 310586 203818 310822 204054
rect 310586 203498 310822 203734
rect 310586 167818 310822 168054
rect 310586 167498 310822 167734
rect 310586 131818 310822 132054
rect 310586 131498 310822 131734
rect 310586 95818 310822 96054
rect 310586 95498 310822 95734
rect 310586 59818 310822 60054
rect 310586 59498 310822 59734
rect 310586 23818 310822 24054
rect 310586 23498 310822 23734
rect 310586 -3342 310822 -3106
rect 310586 -3662 310822 -3426
rect 314186 531418 314422 531654
rect 314186 531098 314422 531334
rect 314186 495418 314422 495654
rect 314186 495098 314422 495334
rect 314186 459418 314422 459654
rect 314186 459098 314422 459334
rect 314186 423418 314422 423654
rect 314186 423098 314422 423334
rect 314186 387418 314422 387654
rect 314186 387098 314422 387334
rect 314186 351418 314422 351654
rect 314186 351098 314422 351334
rect 314186 315418 314422 315654
rect 314186 315098 314422 315334
rect 314186 279418 314422 279654
rect 314186 279098 314422 279334
rect 314186 243418 314422 243654
rect 314186 243098 314422 243334
rect 314186 207418 314422 207654
rect 314186 207098 314422 207334
rect 314186 171418 314422 171654
rect 314186 171098 314422 171334
rect 314186 135418 314422 135654
rect 314186 135098 314422 135334
rect 314186 99418 314422 99654
rect 314186 99098 314422 99334
rect 335786 710122 336022 710358
rect 335786 709802 336022 710038
rect 332186 708282 332422 708518
rect 332186 707962 332422 708198
rect 328586 706442 328822 706678
rect 328586 706122 328822 706358
rect 317786 679018 318022 679254
rect 317786 678698 318022 678934
rect 317786 643018 318022 643254
rect 317786 642698 318022 642934
rect 317786 607018 318022 607254
rect 317786 606698 318022 606934
rect 317786 571018 318022 571254
rect 317786 570698 318022 570934
rect 324986 704602 325222 704838
rect 324986 704282 325222 704518
rect 324986 686218 325222 686454
rect 324986 685898 325222 686134
rect 324986 650218 325222 650454
rect 324986 649898 325222 650134
rect 324986 614218 325222 614454
rect 324986 613898 325222 614134
rect 324986 578218 325222 578454
rect 324986 577898 325222 578134
rect 318478 561222 318714 561458
rect 319214 561222 319450 561458
rect 317786 535018 318022 535254
rect 317786 534698 318022 534934
rect 317786 499018 318022 499254
rect 317786 498698 318022 498934
rect 317786 463018 318022 463254
rect 317786 462698 318022 462934
rect 317786 427018 318022 427254
rect 317786 426698 318022 426934
rect 317786 391018 318022 391254
rect 317786 390698 318022 390934
rect 317786 355018 318022 355254
rect 317786 354698 318022 354934
rect 317786 319018 318022 319254
rect 317786 318698 318022 318934
rect 317786 283018 318022 283254
rect 317786 282698 318022 282934
rect 317786 247018 318022 247254
rect 317786 246698 318022 246934
rect 317786 211018 318022 211254
rect 317786 210698 318022 210934
rect 317786 175018 318022 175254
rect 317786 174698 318022 174934
rect 317786 139018 318022 139254
rect 317786 138698 318022 138934
rect 317786 103018 318022 103254
rect 317786 102698 318022 102934
rect 314186 63418 314422 63654
rect 314186 63098 314422 63334
rect 317786 67018 318022 67254
rect 317786 66698 318022 66934
rect 317786 31018 318022 31254
rect 317786 30698 318022 30934
rect 314186 27418 314422 27654
rect 314186 27098 314422 27334
rect 314186 -5182 314422 -4946
rect 314186 -5502 314422 -5266
rect 299786 -6102 300022 -5866
rect 299786 -6422 300022 -6186
rect 328586 689818 328822 690054
rect 328586 689498 328822 689734
rect 328586 653818 328822 654054
rect 328586 653498 328822 653734
rect 328586 617818 328822 618054
rect 328586 617498 328822 617734
rect 328586 581818 328822 582054
rect 328586 581498 328822 581734
rect 325654 561372 325890 561458
rect 325654 561308 325740 561372
rect 325740 561308 325804 561372
rect 325804 561308 325890 561372
rect 325654 561222 325890 561308
rect 324986 542218 325222 542454
rect 324986 541898 325222 542134
rect 324986 506218 325222 506454
rect 324986 505898 325222 506134
rect 324986 470218 325222 470454
rect 324986 469898 325222 470134
rect 324986 434218 325222 434454
rect 324986 433898 325222 434134
rect 324986 398218 325222 398454
rect 324986 397898 325222 398134
rect 324986 362218 325222 362454
rect 324986 361898 325222 362134
rect 324986 326218 325222 326454
rect 324986 325898 325222 326134
rect 324986 290218 325222 290454
rect 324986 289898 325222 290134
rect 324986 254218 325222 254454
rect 324986 253898 325222 254134
rect 324986 218218 325222 218454
rect 324986 217898 325222 218134
rect 324986 182218 325222 182454
rect 324986 181898 325222 182134
rect 324986 146218 325222 146454
rect 324986 145898 325222 146134
rect 328586 545818 328822 546054
rect 328586 545498 328822 545734
rect 328586 509818 328822 510054
rect 328586 509498 328822 509734
rect 328586 473818 328822 474054
rect 328586 473498 328822 473734
rect 328586 437818 328822 438054
rect 328586 437498 328822 437734
rect 328586 401818 328822 402054
rect 328586 401498 328822 401734
rect 328586 365818 328822 366054
rect 328586 365498 328822 365734
rect 328586 329818 328822 330054
rect 328586 329498 328822 329734
rect 328586 293818 328822 294054
rect 328586 293498 328822 293734
rect 328586 257818 328822 258054
rect 328586 257498 328822 257734
rect 328586 221818 328822 222054
rect 328586 221498 328822 221734
rect 328586 185818 328822 186054
rect 328586 185498 328822 185734
rect 328586 149818 328822 150054
rect 328586 149498 328822 149734
rect 324986 110218 325222 110454
rect 324986 109898 325222 110134
rect 324986 74218 325222 74454
rect 324986 73898 325222 74134
rect 324986 38218 325222 38454
rect 324986 37898 325222 38134
rect 328586 113818 328822 114054
rect 328586 113498 328822 113734
rect 328586 77818 328822 78054
rect 328586 77498 328822 77734
rect 328586 41818 328822 42054
rect 328586 41498 328822 41734
rect 324986 2218 325222 2454
rect 324986 1898 325222 2134
rect 324986 -582 325222 -346
rect 324986 -902 325222 -666
rect 328586 5818 328822 6054
rect 328586 5498 328822 5734
rect 328586 -2422 328822 -2186
rect 328586 -2742 328822 -2506
rect 332186 693418 332422 693654
rect 332186 693098 332422 693334
rect 332186 657418 332422 657654
rect 332186 657098 332422 657334
rect 332186 621418 332422 621654
rect 332186 621098 332422 621334
rect 332186 585418 332422 585654
rect 332186 585098 332422 585334
rect 353786 711042 354022 711278
rect 353786 710722 354022 710958
rect 350186 709202 350422 709438
rect 350186 708882 350422 709118
rect 346586 707362 346822 707598
rect 346586 707042 346822 707278
rect 335786 697018 336022 697254
rect 335786 696698 336022 696934
rect 335786 661018 336022 661254
rect 335786 660698 336022 660934
rect 335786 625018 336022 625254
rect 335786 624698 336022 624934
rect 335786 589018 336022 589254
rect 335786 588698 336022 588934
rect 335038 562582 335274 562818
rect 332186 549418 332422 549654
rect 332186 549098 332422 549334
rect 332186 513418 332422 513654
rect 332186 513098 332422 513334
rect 332186 477418 332422 477654
rect 332186 477098 332422 477334
rect 332186 441418 332422 441654
rect 332186 441098 332422 441334
rect 332186 405418 332422 405654
rect 332186 405098 332422 405334
rect 332186 369418 332422 369654
rect 332186 369098 332422 369334
rect 332186 333418 332422 333654
rect 332186 333098 332422 333334
rect 332186 297418 332422 297654
rect 332186 297098 332422 297334
rect 332186 261418 332422 261654
rect 332186 261098 332422 261334
rect 332186 225418 332422 225654
rect 332186 225098 332422 225334
rect 332186 189418 332422 189654
rect 332186 189098 332422 189334
rect 332186 153418 332422 153654
rect 332186 153098 332422 153334
rect 332186 117418 332422 117654
rect 332186 117098 332422 117334
rect 332186 81418 332422 81654
rect 332186 81098 332422 81334
rect 332186 45418 332422 45654
rect 332186 45098 332422 45334
rect 332186 9418 332422 9654
rect 332186 9098 332422 9334
rect 332186 -4262 332422 -4026
rect 332186 -4582 332422 -4346
rect 342986 705522 343222 705758
rect 342986 705202 343222 705438
rect 342986 668218 343222 668454
rect 342986 667898 343222 668134
rect 342986 632218 343222 632454
rect 342986 631898 343222 632134
rect 342986 596218 343222 596454
rect 342986 595898 343222 596134
rect 336694 562582 336930 562818
rect 337246 561902 337482 562138
rect 342986 560218 343222 560454
rect 342986 559898 343222 560134
rect 335786 553018 336022 553254
rect 335786 552698 336022 552934
rect 335786 517018 336022 517254
rect 335786 516698 336022 516934
rect 335786 481018 336022 481254
rect 335786 480698 336022 480934
rect 335786 445018 336022 445254
rect 335786 444698 336022 444934
rect 335786 409018 336022 409254
rect 335786 408698 336022 408934
rect 335786 373018 336022 373254
rect 335786 372698 336022 372934
rect 335786 337018 336022 337254
rect 335786 336698 336022 336934
rect 335786 301018 336022 301254
rect 335786 300698 336022 300934
rect 335786 265018 336022 265254
rect 335786 264698 336022 264934
rect 335786 229018 336022 229254
rect 335786 228698 336022 228934
rect 335786 193018 336022 193254
rect 335786 192698 336022 192934
rect 335786 157018 336022 157254
rect 335786 156698 336022 156934
rect 335786 121018 336022 121254
rect 335786 120698 336022 120934
rect 335786 85018 336022 85254
rect 335786 84698 336022 84934
rect 335786 49018 336022 49254
rect 335786 48698 336022 48934
rect 335786 13018 336022 13254
rect 335786 12698 336022 12934
rect 317786 -7022 318022 -6786
rect 317786 -7342 318022 -7106
rect 342986 524218 343222 524454
rect 342986 523898 343222 524134
rect 342986 488218 343222 488454
rect 342986 487898 343222 488134
rect 342986 452218 343222 452454
rect 342986 451898 343222 452134
rect 342986 416218 343222 416454
rect 342986 415898 343222 416134
rect 342986 380218 343222 380454
rect 342986 379898 343222 380134
rect 342986 344218 343222 344454
rect 342986 343898 343222 344134
rect 342986 308218 343222 308454
rect 342986 307898 343222 308134
rect 342986 272218 343222 272454
rect 342986 271898 343222 272134
rect 342986 236218 343222 236454
rect 342986 235898 343222 236134
rect 342986 200218 343222 200454
rect 342986 199898 343222 200134
rect 342986 164218 343222 164454
rect 342986 163898 343222 164134
rect 342986 128218 343222 128454
rect 342986 127898 343222 128134
rect 342986 92218 343222 92454
rect 342986 91898 343222 92134
rect 346586 671818 346822 672054
rect 346586 671498 346822 671734
rect 346586 635818 346822 636054
rect 346586 635498 346822 635734
rect 346586 599818 346822 600054
rect 346586 599498 346822 599734
rect 346586 563818 346822 564054
rect 346586 563498 346822 563734
rect 346586 527818 346822 528054
rect 346586 527498 346822 527734
rect 346586 491818 346822 492054
rect 346586 491498 346822 491734
rect 346586 455818 346822 456054
rect 346586 455498 346822 455734
rect 346586 419818 346822 420054
rect 346586 419498 346822 419734
rect 346586 383818 346822 384054
rect 346586 383498 346822 383734
rect 346586 347818 346822 348054
rect 346586 347498 346822 347734
rect 346586 311818 346822 312054
rect 346586 311498 346822 311734
rect 346586 275818 346822 276054
rect 346586 275498 346822 275734
rect 346586 239818 346822 240054
rect 346586 239498 346822 239734
rect 346586 203818 346822 204054
rect 346586 203498 346822 203734
rect 346586 167818 346822 168054
rect 346586 167498 346822 167734
rect 346586 131818 346822 132054
rect 346586 131498 346822 131734
rect 346586 95818 346822 96054
rect 346586 95498 346822 95734
rect 342986 56218 343222 56454
rect 342986 55898 343222 56134
rect 342986 20218 343222 20454
rect 342986 19898 343222 20134
rect 342986 -1502 343222 -1266
rect 342986 -1822 343222 -1586
rect 346586 59818 346822 60054
rect 346586 59498 346822 59734
rect 346586 23818 346822 24054
rect 346586 23498 346822 23734
rect 346586 -3342 346822 -3106
rect 346586 -3662 346822 -3426
rect 350186 675418 350422 675654
rect 350186 675098 350422 675334
rect 350186 639418 350422 639654
rect 350186 639098 350422 639334
rect 350186 603418 350422 603654
rect 350186 603098 350422 603334
rect 350186 567418 350422 567654
rect 350186 567098 350422 567334
rect 371786 710122 372022 710358
rect 371786 709802 372022 710038
rect 368186 708282 368422 708518
rect 368186 707962 368422 708198
rect 364586 706442 364822 706678
rect 364586 706122 364822 706358
rect 353786 679018 354022 679254
rect 353786 678698 354022 678934
rect 353786 643018 354022 643254
rect 353786 642698 354022 642934
rect 353786 607018 354022 607254
rect 353786 606698 354022 606934
rect 353786 571018 354022 571254
rect 353786 570698 354022 570934
rect 350186 531418 350422 531654
rect 350186 531098 350422 531334
rect 350186 495418 350422 495654
rect 350186 495098 350422 495334
rect 350186 459418 350422 459654
rect 350186 459098 350422 459334
rect 350186 423418 350422 423654
rect 350186 423098 350422 423334
rect 350186 387418 350422 387654
rect 350186 387098 350422 387334
rect 350186 351418 350422 351654
rect 350186 351098 350422 351334
rect 350186 315418 350422 315654
rect 350186 315098 350422 315334
rect 350186 279418 350422 279654
rect 350186 279098 350422 279334
rect 350186 243418 350422 243654
rect 350186 243098 350422 243334
rect 350186 207418 350422 207654
rect 350186 207098 350422 207334
rect 350186 171418 350422 171654
rect 350186 171098 350422 171334
rect 350186 135418 350422 135654
rect 350186 135098 350422 135334
rect 350186 99418 350422 99654
rect 350186 99098 350422 99334
rect 350186 63418 350422 63654
rect 350186 63098 350422 63334
rect 350186 27418 350422 27654
rect 350186 27098 350422 27334
rect 350186 -5182 350422 -4946
rect 350186 -5502 350422 -5266
rect 360986 704602 361222 704838
rect 360986 704282 361222 704518
rect 360986 686218 361222 686454
rect 360986 685898 361222 686134
rect 360986 650218 361222 650454
rect 360986 649898 361222 650134
rect 360986 614218 361222 614454
rect 360986 613898 361222 614134
rect 360986 578218 361222 578454
rect 360986 577898 361222 578134
rect 357302 562582 357538 562818
rect 353786 535018 354022 535254
rect 353786 534698 354022 534934
rect 353786 499018 354022 499254
rect 353786 498698 354022 498934
rect 353786 463018 354022 463254
rect 353786 462698 354022 462934
rect 353786 427018 354022 427254
rect 353786 426698 354022 426934
rect 353786 391018 354022 391254
rect 353786 390698 354022 390934
rect 353786 355018 354022 355254
rect 353786 354698 354022 354934
rect 353786 319018 354022 319254
rect 353786 318698 354022 318934
rect 353786 283018 354022 283254
rect 353786 282698 354022 282934
rect 353786 247018 354022 247254
rect 353786 246698 354022 246934
rect 353786 211018 354022 211254
rect 353786 210698 354022 210934
rect 360986 542218 361222 542454
rect 360986 541898 361222 542134
rect 360986 506218 361222 506454
rect 360986 505898 361222 506134
rect 360986 470218 361222 470454
rect 360986 469898 361222 470134
rect 360986 434218 361222 434454
rect 360986 433898 361222 434134
rect 360986 398218 361222 398454
rect 360986 397898 361222 398134
rect 360986 362218 361222 362454
rect 360986 361898 361222 362134
rect 360986 326218 361222 326454
rect 360986 325898 361222 326134
rect 360986 290218 361222 290454
rect 360986 289898 361222 290134
rect 360986 254218 361222 254454
rect 360986 253898 361222 254134
rect 360986 218218 361222 218454
rect 360986 217898 361222 218134
rect 360986 182218 361222 182454
rect 360986 181898 361222 182134
rect 353786 175018 354022 175254
rect 353786 174698 354022 174934
rect 353786 139018 354022 139254
rect 353786 138698 354022 138934
rect 353786 103018 354022 103254
rect 353786 102698 354022 102934
rect 353786 67018 354022 67254
rect 353786 66698 354022 66934
rect 353786 31018 354022 31254
rect 353786 30698 354022 30934
rect 335786 -6102 336022 -5866
rect 335786 -6422 336022 -6186
rect 360986 146218 361222 146454
rect 360986 145898 361222 146134
rect 360986 110218 361222 110454
rect 360986 109898 361222 110134
rect 360986 74218 361222 74454
rect 360986 73898 361222 74134
rect 360986 38218 361222 38454
rect 360986 37898 361222 38134
rect 360986 2218 361222 2454
rect 360986 1898 361222 2134
rect 360986 -582 361222 -346
rect 360986 -902 361222 -666
rect 364586 689818 364822 690054
rect 364586 689498 364822 689734
rect 364586 653818 364822 654054
rect 364586 653498 364822 653734
rect 364586 617818 364822 618054
rect 364586 617498 364822 617734
rect 364586 581818 364822 582054
rect 364586 581498 364822 581734
rect 368186 693418 368422 693654
rect 368186 693098 368422 693334
rect 368186 657418 368422 657654
rect 368186 657098 368422 657334
rect 368186 621418 368422 621654
rect 368186 621098 368422 621334
rect 368186 585418 368422 585654
rect 368186 585098 368422 585334
rect 366870 561902 367106 562138
rect 364586 545818 364822 546054
rect 364586 545498 364822 545734
rect 364586 509818 364822 510054
rect 364586 509498 364822 509734
rect 364586 473818 364822 474054
rect 364586 473498 364822 473734
rect 364586 437818 364822 438054
rect 364586 437498 364822 437734
rect 364586 401818 364822 402054
rect 364586 401498 364822 401734
rect 364586 365818 364822 366054
rect 364586 365498 364822 365734
rect 364586 329818 364822 330054
rect 364586 329498 364822 329734
rect 364586 293818 364822 294054
rect 364586 293498 364822 293734
rect 364586 257818 364822 258054
rect 364586 257498 364822 257734
rect 364586 221818 364822 222054
rect 364586 221498 364822 221734
rect 364586 185818 364822 186054
rect 364586 185498 364822 185734
rect 364586 149818 364822 150054
rect 364586 149498 364822 149734
rect 364586 113818 364822 114054
rect 364586 113498 364822 113734
rect 389786 711042 390022 711278
rect 389786 710722 390022 710958
rect 386186 709202 386422 709438
rect 386186 708882 386422 709118
rect 382586 707362 382822 707598
rect 382586 707042 382822 707278
rect 371786 697018 372022 697254
rect 371786 696698 372022 696934
rect 371786 661018 372022 661254
rect 371786 660698 372022 660934
rect 371786 625018 372022 625254
rect 371786 624698 372022 624934
rect 371786 589018 372022 589254
rect 371786 588698 372022 588934
rect 370366 562582 370602 562818
rect 369262 561902 369498 562138
rect 368186 549418 368422 549654
rect 368186 549098 368422 549334
rect 368186 513418 368422 513654
rect 368186 513098 368422 513334
rect 368186 477418 368422 477654
rect 368186 477098 368422 477334
rect 368186 441418 368422 441654
rect 368186 441098 368422 441334
rect 368186 405418 368422 405654
rect 368186 405098 368422 405334
rect 368186 369418 368422 369654
rect 368186 369098 368422 369334
rect 368186 333418 368422 333654
rect 368186 333098 368422 333334
rect 368186 297418 368422 297654
rect 368186 297098 368422 297334
rect 368186 261418 368422 261654
rect 368186 261098 368422 261334
rect 368186 225418 368422 225654
rect 368186 225098 368422 225334
rect 368186 189418 368422 189654
rect 368186 189098 368422 189334
rect 368186 153418 368422 153654
rect 368186 153098 368422 153334
rect 368186 117418 368422 117654
rect 368186 117098 368422 117334
rect 364586 77818 364822 78054
rect 364586 77498 364822 77734
rect 364586 41818 364822 42054
rect 364586 41498 364822 41734
rect 368186 81418 368422 81654
rect 368186 81098 368422 81334
rect 368186 45418 368422 45654
rect 368186 45098 368422 45334
rect 364586 5818 364822 6054
rect 364586 5498 364822 5734
rect 364586 -2422 364822 -2186
rect 364586 -2742 364822 -2506
rect 368186 9418 368422 9654
rect 368186 9098 368422 9334
rect 368186 -4262 368422 -4026
rect 368186 -4582 368422 -4346
rect 378986 705522 379222 705758
rect 378986 705202 379222 705438
rect 378986 668218 379222 668454
rect 378986 667898 379222 668134
rect 378986 632218 379222 632454
rect 378986 631898 379222 632134
rect 378986 596218 379222 596454
rect 378986 595898 379222 596134
rect 371786 553018 372022 553254
rect 371786 552698 372022 552934
rect 371786 517018 372022 517254
rect 371786 516698 372022 516934
rect 371786 481018 372022 481254
rect 371786 480698 372022 480934
rect 371786 445018 372022 445254
rect 371786 444698 372022 444934
rect 371786 409018 372022 409254
rect 371786 408698 372022 408934
rect 371786 373018 372022 373254
rect 371786 372698 372022 372934
rect 371786 337018 372022 337254
rect 371786 336698 372022 336934
rect 371786 301018 372022 301254
rect 371786 300698 372022 300934
rect 371786 265018 372022 265254
rect 371786 264698 372022 264934
rect 371786 229018 372022 229254
rect 371786 228698 372022 228934
rect 371786 193018 372022 193254
rect 371786 192698 372022 192934
rect 371786 157018 372022 157254
rect 371786 156698 372022 156934
rect 371786 121018 372022 121254
rect 371786 120698 372022 120934
rect 371786 85018 372022 85254
rect 371786 84698 372022 84934
rect 371786 49018 372022 49254
rect 371786 48698 372022 48934
rect 371786 13018 372022 13254
rect 371786 12698 372022 12934
rect 353786 -7022 354022 -6786
rect 353786 -7342 354022 -7106
rect 378986 560218 379222 560454
rect 378986 559898 379222 560134
rect 378986 524218 379222 524454
rect 378986 523898 379222 524134
rect 378986 488218 379222 488454
rect 378986 487898 379222 488134
rect 378986 452218 379222 452454
rect 378986 451898 379222 452134
rect 378986 416218 379222 416454
rect 378986 415898 379222 416134
rect 378986 380218 379222 380454
rect 378986 379898 379222 380134
rect 378986 344218 379222 344454
rect 378986 343898 379222 344134
rect 378986 308218 379222 308454
rect 378986 307898 379222 308134
rect 378986 272218 379222 272454
rect 378986 271898 379222 272134
rect 378986 236218 379222 236454
rect 378986 235898 379222 236134
rect 378986 200218 379222 200454
rect 378986 199898 379222 200134
rect 378986 164218 379222 164454
rect 378986 163898 379222 164134
rect 378986 128218 379222 128454
rect 378986 127898 379222 128134
rect 378986 92218 379222 92454
rect 378986 91898 379222 92134
rect 378986 56218 379222 56454
rect 378986 55898 379222 56134
rect 378986 20218 379222 20454
rect 378986 19898 379222 20134
rect 378986 -1502 379222 -1266
rect 378986 -1822 379222 -1586
rect 382586 671818 382822 672054
rect 382586 671498 382822 671734
rect 382586 635818 382822 636054
rect 382586 635498 382822 635734
rect 382586 599818 382822 600054
rect 382586 599498 382822 599734
rect 382586 563818 382822 564054
rect 382586 563498 382822 563734
rect 386186 675418 386422 675654
rect 386186 675098 386422 675334
rect 386186 639418 386422 639654
rect 386186 639098 386422 639334
rect 386186 603418 386422 603654
rect 386186 603098 386422 603334
rect 386186 567418 386422 567654
rect 386186 567098 386422 567334
rect 382586 527818 382822 528054
rect 382586 527498 382822 527734
rect 382586 491818 382822 492054
rect 382586 491498 382822 491734
rect 382586 455818 382822 456054
rect 382586 455498 382822 455734
rect 382586 419818 382822 420054
rect 382586 419498 382822 419734
rect 382586 383818 382822 384054
rect 382586 383498 382822 383734
rect 382586 347818 382822 348054
rect 382586 347498 382822 347734
rect 382586 311818 382822 312054
rect 382586 311498 382822 311734
rect 382586 275818 382822 276054
rect 382586 275498 382822 275734
rect 382586 239818 382822 240054
rect 382586 239498 382822 239734
rect 382586 203818 382822 204054
rect 382586 203498 382822 203734
rect 382586 167818 382822 168054
rect 382586 167498 382822 167734
rect 382586 131818 382822 132054
rect 382586 131498 382822 131734
rect 382586 95818 382822 96054
rect 382586 95498 382822 95734
rect 382586 59818 382822 60054
rect 382586 59498 382822 59734
rect 382586 23818 382822 24054
rect 382586 23498 382822 23734
rect 382586 -3342 382822 -3106
rect 382586 -3662 382822 -3426
rect 386186 531418 386422 531654
rect 386186 531098 386422 531334
rect 386186 495418 386422 495654
rect 386186 495098 386422 495334
rect 386186 459418 386422 459654
rect 386186 459098 386422 459334
rect 386186 423418 386422 423654
rect 386186 423098 386422 423334
rect 386186 387418 386422 387654
rect 386186 387098 386422 387334
rect 386186 351418 386422 351654
rect 386186 351098 386422 351334
rect 386186 315418 386422 315654
rect 386186 315098 386422 315334
rect 386186 279418 386422 279654
rect 386186 279098 386422 279334
rect 386186 243418 386422 243654
rect 386186 243098 386422 243334
rect 386186 207418 386422 207654
rect 386186 207098 386422 207334
rect 386186 171418 386422 171654
rect 386186 171098 386422 171334
rect 386186 135418 386422 135654
rect 386186 135098 386422 135334
rect 386186 99418 386422 99654
rect 386186 99098 386422 99334
rect 386186 63418 386422 63654
rect 386186 63098 386422 63334
rect 386186 27418 386422 27654
rect 386186 27098 386422 27334
rect 386186 -5182 386422 -4946
rect 386186 -5502 386422 -5266
rect 407786 710122 408022 710358
rect 407786 709802 408022 710038
rect 404186 708282 404422 708518
rect 404186 707962 404422 708198
rect 400586 706442 400822 706678
rect 400586 706122 400822 706358
rect 389786 679018 390022 679254
rect 389786 678698 390022 678934
rect 389786 643018 390022 643254
rect 389786 642698 390022 642934
rect 389786 607018 390022 607254
rect 389786 606698 390022 606934
rect 389786 571018 390022 571254
rect 389786 570698 390022 570934
rect 396986 704602 397222 704838
rect 396986 704282 397222 704518
rect 396986 686218 397222 686454
rect 396986 685898 397222 686134
rect 396986 650218 397222 650454
rect 396986 649898 397222 650134
rect 396986 614218 397222 614454
rect 396986 613898 397222 614134
rect 396986 578218 397222 578454
rect 396986 577898 397222 578134
rect 393182 562582 393418 562818
rect 389786 535018 390022 535254
rect 389786 534698 390022 534934
rect 389786 499018 390022 499254
rect 389786 498698 390022 498934
rect 389786 463018 390022 463254
rect 389786 462698 390022 462934
rect 389786 427018 390022 427254
rect 389786 426698 390022 426934
rect 389786 391018 390022 391254
rect 389786 390698 390022 390934
rect 389786 355018 390022 355254
rect 389786 354698 390022 354934
rect 389786 319018 390022 319254
rect 389786 318698 390022 318934
rect 389786 283018 390022 283254
rect 389786 282698 390022 282934
rect 389786 247018 390022 247254
rect 389786 246698 390022 246934
rect 389786 211018 390022 211254
rect 389786 210698 390022 210934
rect 389786 175018 390022 175254
rect 389786 174698 390022 174934
rect 389786 139018 390022 139254
rect 389786 138698 390022 138934
rect 389786 103018 390022 103254
rect 389786 102698 390022 102934
rect 389786 67018 390022 67254
rect 389786 66698 390022 66934
rect 389786 31018 390022 31254
rect 389786 30698 390022 30934
rect 371786 -6102 372022 -5866
rect 371786 -6422 372022 -6186
rect 396986 542218 397222 542454
rect 396986 541898 397222 542134
rect 396986 506218 397222 506454
rect 396986 505898 397222 506134
rect 396986 470218 397222 470454
rect 396986 469898 397222 470134
rect 396986 434218 397222 434454
rect 396986 433898 397222 434134
rect 396986 398218 397222 398454
rect 396986 397898 397222 398134
rect 396986 362218 397222 362454
rect 396986 361898 397222 362134
rect 396986 326218 397222 326454
rect 396986 325898 397222 326134
rect 396986 290218 397222 290454
rect 396986 289898 397222 290134
rect 396986 254218 397222 254454
rect 396986 253898 397222 254134
rect 396986 218218 397222 218454
rect 396986 217898 397222 218134
rect 396986 182218 397222 182454
rect 396986 181898 397222 182134
rect 396986 146218 397222 146454
rect 396986 145898 397222 146134
rect 396986 110218 397222 110454
rect 396986 109898 397222 110134
rect 396986 74218 397222 74454
rect 396986 73898 397222 74134
rect 396986 38218 397222 38454
rect 396986 37898 397222 38134
rect 396986 2218 397222 2454
rect 396986 1898 397222 2134
rect 396986 -582 397222 -346
rect 396986 -902 397222 -666
rect 400586 689818 400822 690054
rect 400586 689498 400822 689734
rect 400586 653818 400822 654054
rect 400586 653498 400822 653734
rect 400586 617818 400822 618054
rect 400586 617498 400822 617734
rect 400586 581818 400822 582054
rect 400586 581498 400822 581734
rect 400586 545818 400822 546054
rect 400586 545498 400822 545734
rect 400586 509818 400822 510054
rect 400586 509498 400822 509734
rect 400586 473818 400822 474054
rect 400586 473498 400822 473734
rect 400586 437818 400822 438054
rect 400586 437498 400822 437734
rect 400586 401818 400822 402054
rect 400586 401498 400822 401734
rect 400586 365818 400822 366054
rect 400586 365498 400822 365734
rect 400586 329818 400822 330054
rect 400586 329498 400822 329734
rect 400586 293818 400822 294054
rect 400586 293498 400822 293734
rect 400586 257818 400822 258054
rect 400586 257498 400822 257734
rect 400586 221818 400822 222054
rect 400586 221498 400822 221734
rect 400586 185818 400822 186054
rect 400586 185498 400822 185734
rect 400586 149818 400822 150054
rect 400586 149498 400822 149734
rect 400586 113818 400822 114054
rect 400586 113498 400822 113734
rect 400586 77818 400822 78054
rect 400586 77498 400822 77734
rect 400586 41818 400822 42054
rect 400586 41498 400822 41734
rect 400586 5818 400822 6054
rect 400586 5498 400822 5734
rect 400586 -2422 400822 -2186
rect 400586 -2742 400822 -2506
rect 404186 693418 404422 693654
rect 404186 693098 404422 693334
rect 404186 657418 404422 657654
rect 404186 657098 404422 657334
rect 404186 621418 404422 621654
rect 404186 621098 404422 621334
rect 404186 585418 404422 585654
rect 404186 585098 404422 585334
rect 425786 711042 426022 711278
rect 425786 710722 426022 710958
rect 422186 709202 422422 709438
rect 422186 708882 422422 709118
rect 418586 707362 418822 707598
rect 418586 707042 418822 707278
rect 407786 697018 408022 697254
rect 407786 696698 408022 696934
rect 407786 661018 408022 661254
rect 407786 660698 408022 660934
rect 407786 625018 408022 625254
rect 407786 624698 408022 624934
rect 407786 589018 408022 589254
rect 407786 588698 408022 588934
rect 406246 561902 406482 562138
rect 404186 549418 404422 549654
rect 404186 549098 404422 549334
rect 404186 513418 404422 513654
rect 404186 513098 404422 513334
rect 404186 477418 404422 477654
rect 404186 477098 404422 477334
rect 404186 441418 404422 441654
rect 404186 441098 404422 441334
rect 404186 405418 404422 405654
rect 404186 405098 404422 405334
rect 404186 369418 404422 369654
rect 404186 369098 404422 369334
rect 404186 333418 404422 333654
rect 404186 333098 404422 333334
rect 404186 297418 404422 297654
rect 404186 297098 404422 297334
rect 404186 261418 404422 261654
rect 404186 261098 404422 261334
rect 404186 225418 404422 225654
rect 404186 225098 404422 225334
rect 404186 189418 404422 189654
rect 404186 189098 404422 189334
rect 404186 153418 404422 153654
rect 404186 153098 404422 153334
rect 404186 117418 404422 117654
rect 404186 117098 404422 117334
rect 404186 81418 404422 81654
rect 404186 81098 404422 81334
rect 404186 45418 404422 45654
rect 404186 45098 404422 45334
rect 404186 9418 404422 9654
rect 404186 9098 404422 9334
rect 404186 -4262 404422 -4026
rect 404186 -4582 404422 -4346
rect 414986 705522 415222 705758
rect 414986 705202 415222 705438
rect 414986 668218 415222 668454
rect 414986 667898 415222 668134
rect 414986 632218 415222 632454
rect 414986 631898 415222 632134
rect 414986 596218 415222 596454
rect 414986 595898 415222 596134
rect 414986 560218 415222 560454
rect 414986 559898 415222 560134
rect 407786 553018 408022 553254
rect 407786 552698 408022 552934
rect 407786 517018 408022 517254
rect 407786 516698 408022 516934
rect 407786 481018 408022 481254
rect 407786 480698 408022 480934
rect 407786 445018 408022 445254
rect 407786 444698 408022 444934
rect 407786 409018 408022 409254
rect 407786 408698 408022 408934
rect 407786 373018 408022 373254
rect 407786 372698 408022 372934
rect 407786 337018 408022 337254
rect 407786 336698 408022 336934
rect 407786 301018 408022 301254
rect 407786 300698 408022 300934
rect 407786 265018 408022 265254
rect 407786 264698 408022 264934
rect 407786 229018 408022 229254
rect 407786 228698 408022 228934
rect 407786 193018 408022 193254
rect 407786 192698 408022 192934
rect 407786 157018 408022 157254
rect 407786 156698 408022 156934
rect 407786 121018 408022 121254
rect 407786 120698 408022 120934
rect 407786 85018 408022 85254
rect 407786 84698 408022 84934
rect 407786 49018 408022 49254
rect 407786 48698 408022 48934
rect 407786 13018 408022 13254
rect 407786 12698 408022 12934
rect 389786 -7022 390022 -6786
rect 389786 -7342 390022 -7106
rect 414986 524218 415222 524454
rect 414986 523898 415222 524134
rect 414986 488218 415222 488454
rect 414986 487898 415222 488134
rect 414986 452218 415222 452454
rect 414986 451898 415222 452134
rect 414986 416218 415222 416454
rect 414986 415898 415222 416134
rect 414986 380218 415222 380454
rect 414986 379898 415222 380134
rect 414986 344218 415222 344454
rect 414986 343898 415222 344134
rect 414986 308218 415222 308454
rect 414986 307898 415222 308134
rect 414986 272218 415222 272454
rect 414986 271898 415222 272134
rect 414986 236218 415222 236454
rect 414986 235898 415222 236134
rect 414986 200218 415222 200454
rect 414986 199898 415222 200134
rect 414986 164218 415222 164454
rect 414986 163898 415222 164134
rect 414986 128218 415222 128454
rect 414986 127898 415222 128134
rect 414986 92218 415222 92454
rect 414986 91898 415222 92134
rect 414986 56218 415222 56454
rect 414986 55898 415222 56134
rect 414986 20218 415222 20454
rect 414986 19898 415222 20134
rect 414986 -1502 415222 -1266
rect 414986 -1822 415222 -1586
rect 418586 671818 418822 672054
rect 418586 671498 418822 671734
rect 418586 635818 418822 636054
rect 418586 635498 418822 635734
rect 418586 599818 418822 600054
rect 418586 599498 418822 599734
rect 418586 563818 418822 564054
rect 418586 563498 418822 563734
rect 418586 527818 418822 528054
rect 418586 527498 418822 527734
rect 418586 491818 418822 492054
rect 418586 491498 418822 491734
rect 418586 455818 418822 456054
rect 418586 455498 418822 455734
rect 418586 419818 418822 420054
rect 418586 419498 418822 419734
rect 418586 383818 418822 384054
rect 418586 383498 418822 383734
rect 418586 347818 418822 348054
rect 418586 347498 418822 347734
rect 418586 311818 418822 312054
rect 418586 311498 418822 311734
rect 418586 275818 418822 276054
rect 418586 275498 418822 275734
rect 418586 239818 418822 240054
rect 418586 239498 418822 239734
rect 418586 203818 418822 204054
rect 418586 203498 418822 203734
rect 418586 167818 418822 168054
rect 418586 167498 418822 167734
rect 418586 131818 418822 132054
rect 418586 131498 418822 131734
rect 418586 95818 418822 96054
rect 418586 95498 418822 95734
rect 418586 59818 418822 60054
rect 418586 59498 418822 59734
rect 418586 23818 418822 24054
rect 418586 23498 418822 23734
rect 418586 -3342 418822 -3106
rect 418586 -3662 418822 -3426
rect 422186 675418 422422 675654
rect 422186 675098 422422 675334
rect 422186 639418 422422 639654
rect 422186 639098 422422 639334
rect 422186 603418 422422 603654
rect 422186 603098 422422 603334
rect 422186 567418 422422 567654
rect 422186 567098 422422 567334
rect 443786 710122 444022 710358
rect 443786 709802 444022 710038
rect 440186 708282 440422 708518
rect 440186 707962 440422 708198
rect 436586 706442 436822 706678
rect 436586 706122 436822 706358
rect 425786 679018 426022 679254
rect 425786 678698 426022 678934
rect 425786 643018 426022 643254
rect 425786 642698 426022 642934
rect 425786 607018 426022 607254
rect 425786 606698 426022 606934
rect 425786 571018 426022 571254
rect 425786 570698 426022 570934
rect 424278 562732 424514 562818
rect 424278 562668 424364 562732
rect 424364 562668 424428 562732
rect 424428 562668 424514 562732
rect 424278 562582 424514 562668
rect 422186 531418 422422 531654
rect 422186 531098 422422 531334
rect 422186 495418 422422 495654
rect 422186 495098 422422 495334
rect 422186 459418 422422 459654
rect 422186 459098 422422 459334
rect 422186 423418 422422 423654
rect 422186 423098 422422 423334
rect 422186 387418 422422 387654
rect 422186 387098 422422 387334
rect 422186 351418 422422 351654
rect 422186 351098 422422 351334
rect 422186 315418 422422 315654
rect 422186 315098 422422 315334
rect 422186 279418 422422 279654
rect 422186 279098 422422 279334
rect 422186 243418 422422 243654
rect 422186 243098 422422 243334
rect 422186 207418 422422 207654
rect 422186 207098 422422 207334
rect 422186 171418 422422 171654
rect 422186 171098 422422 171334
rect 422186 135418 422422 135654
rect 422186 135098 422422 135334
rect 422186 99418 422422 99654
rect 422186 99098 422422 99334
rect 422186 63418 422422 63654
rect 422186 63098 422422 63334
rect 422186 27418 422422 27654
rect 422186 27098 422422 27334
rect 422186 -5182 422422 -4946
rect 422186 -5502 422422 -5266
rect 432986 704602 433222 704838
rect 432986 704282 433222 704518
rect 432986 686218 433222 686454
rect 432986 685898 433222 686134
rect 432986 650218 433222 650454
rect 432986 649898 433222 650134
rect 432986 614218 433222 614454
rect 432986 613898 433222 614134
rect 432986 578218 433222 578454
rect 432986 577898 433222 578134
rect 428326 562732 428562 562818
rect 428326 562668 428412 562732
rect 428412 562668 428476 562732
rect 428476 562668 428562 562732
rect 428326 562582 428562 562668
rect 425786 535018 426022 535254
rect 425786 534698 426022 534934
rect 425786 499018 426022 499254
rect 425786 498698 426022 498934
rect 425786 463018 426022 463254
rect 425786 462698 426022 462934
rect 425786 427018 426022 427254
rect 425786 426698 426022 426934
rect 425786 391018 426022 391254
rect 425786 390698 426022 390934
rect 425786 355018 426022 355254
rect 425786 354698 426022 354934
rect 425786 319018 426022 319254
rect 425786 318698 426022 318934
rect 425786 283018 426022 283254
rect 425786 282698 426022 282934
rect 425786 247018 426022 247254
rect 425786 246698 426022 246934
rect 425786 211018 426022 211254
rect 425786 210698 426022 210934
rect 425786 175018 426022 175254
rect 425786 174698 426022 174934
rect 425786 139018 426022 139254
rect 425786 138698 426022 138934
rect 425786 103018 426022 103254
rect 425786 102698 426022 102934
rect 425786 67018 426022 67254
rect 425786 66698 426022 66934
rect 425786 31018 426022 31254
rect 425786 30698 426022 30934
rect 407786 -6102 408022 -5866
rect 407786 -6422 408022 -6186
rect 436586 689818 436822 690054
rect 436586 689498 436822 689734
rect 436586 653818 436822 654054
rect 436586 653498 436822 653734
rect 436586 617818 436822 618054
rect 436586 617498 436822 617734
rect 436586 581818 436822 582054
rect 436586 581498 436822 581734
rect 436054 562732 436290 562818
rect 436054 562668 436140 562732
rect 436140 562668 436204 562732
rect 436204 562668 436290 562732
rect 436054 562582 436290 562668
rect 432986 542218 433222 542454
rect 432986 541898 433222 542134
rect 432986 506218 433222 506454
rect 432986 505898 433222 506134
rect 432986 470218 433222 470454
rect 432986 469898 433222 470134
rect 432986 434218 433222 434454
rect 432986 433898 433222 434134
rect 432986 398218 433222 398454
rect 432986 397898 433222 398134
rect 432986 362218 433222 362454
rect 432986 361898 433222 362134
rect 432986 326218 433222 326454
rect 432986 325898 433222 326134
rect 436586 545818 436822 546054
rect 436586 545498 436822 545734
rect 436586 509818 436822 510054
rect 436586 509498 436822 509734
rect 436586 473818 436822 474054
rect 436586 473498 436822 473734
rect 436586 437818 436822 438054
rect 436586 437498 436822 437734
rect 436586 401818 436822 402054
rect 436586 401498 436822 401734
rect 436586 365818 436822 366054
rect 436586 365498 436822 365734
rect 436586 329818 436822 330054
rect 436586 329498 436822 329734
rect 432986 290218 433222 290454
rect 432986 289898 433222 290134
rect 436586 293818 436822 294054
rect 436586 293498 436822 293734
rect 432986 254218 433222 254454
rect 432986 253898 433222 254134
rect 436586 257818 436822 258054
rect 436586 257498 436822 257734
rect 432986 218218 433222 218454
rect 432986 217898 433222 218134
rect 432986 182218 433222 182454
rect 432986 181898 433222 182134
rect 436586 221818 436822 222054
rect 436586 221498 436822 221734
rect 436586 185818 436822 186054
rect 436586 185498 436822 185734
rect 432986 146218 433222 146454
rect 432986 145898 433222 146134
rect 432986 110218 433222 110454
rect 432986 109898 433222 110134
rect 432986 74218 433222 74454
rect 432986 73898 433222 74134
rect 436586 149818 436822 150054
rect 436586 149498 436822 149734
rect 436586 113818 436822 114054
rect 436586 113498 436822 113734
rect 436586 77818 436822 78054
rect 436586 77498 436822 77734
rect 436586 41818 436822 42054
rect 436586 41498 436822 41734
rect 432986 38218 433222 38454
rect 432986 37898 433222 38134
rect 432986 2218 433222 2454
rect 432986 1898 433222 2134
rect 432986 -582 433222 -346
rect 432986 -902 433222 -666
rect 436586 5818 436822 6054
rect 436586 5498 436822 5734
rect 436586 -2422 436822 -2186
rect 436586 -2742 436822 -2506
rect 440186 693418 440422 693654
rect 440186 693098 440422 693334
rect 440186 657418 440422 657654
rect 440186 657098 440422 657334
rect 440186 621418 440422 621654
rect 440186 621098 440422 621334
rect 440186 585418 440422 585654
rect 440186 585098 440422 585334
rect 440186 549418 440422 549654
rect 440186 549098 440422 549334
rect 440186 513418 440422 513654
rect 440186 513098 440422 513334
rect 440186 477418 440422 477654
rect 440186 477098 440422 477334
rect 440186 441418 440422 441654
rect 440186 441098 440422 441334
rect 440186 405418 440422 405654
rect 440186 405098 440422 405334
rect 440186 369418 440422 369654
rect 440186 369098 440422 369334
rect 440186 333418 440422 333654
rect 440186 333098 440422 333334
rect 440186 297418 440422 297654
rect 440186 297098 440422 297334
rect 440186 261418 440422 261654
rect 440186 261098 440422 261334
rect 440186 225418 440422 225654
rect 440186 225098 440422 225334
rect 440186 189418 440422 189654
rect 440186 189098 440422 189334
rect 440186 153418 440422 153654
rect 440186 153098 440422 153334
rect 440186 117418 440422 117654
rect 440186 117098 440422 117334
rect 440186 81418 440422 81654
rect 440186 81098 440422 81334
rect 440186 45418 440422 45654
rect 440186 45098 440422 45334
rect 440186 9418 440422 9654
rect 440186 9098 440422 9334
rect 440186 -4262 440422 -4026
rect 440186 -4582 440422 -4346
rect 461786 711042 462022 711278
rect 461786 710722 462022 710958
rect 458186 709202 458422 709438
rect 458186 708882 458422 709118
rect 454586 707362 454822 707598
rect 454586 707042 454822 707278
rect 443786 697018 444022 697254
rect 443786 696698 444022 696934
rect 443786 661018 444022 661254
rect 443786 660698 444022 660934
rect 443786 625018 444022 625254
rect 443786 624698 444022 624934
rect 443786 589018 444022 589254
rect 443786 588698 444022 588934
rect 450986 705522 451222 705758
rect 450986 705202 451222 705438
rect 450986 668218 451222 668454
rect 450986 667898 451222 668134
rect 450986 632218 451222 632454
rect 450986 631898 451222 632134
rect 450986 596218 451222 596454
rect 450986 595898 451222 596134
rect 443786 553018 444022 553254
rect 443786 552698 444022 552934
rect 443786 517018 444022 517254
rect 443786 516698 444022 516934
rect 443786 481018 444022 481254
rect 443786 480698 444022 480934
rect 443786 445018 444022 445254
rect 443786 444698 444022 444934
rect 443786 409018 444022 409254
rect 443786 408698 444022 408934
rect 443786 373018 444022 373254
rect 443786 372698 444022 372934
rect 443786 337018 444022 337254
rect 443786 336698 444022 336934
rect 443786 301018 444022 301254
rect 443786 300698 444022 300934
rect 443786 265018 444022 265254
rect 443786 264698 444022 264934
rect 443786 229018 444022 229254
rect 443786 228698 444022 228934
rect 443786 193018 444022 193254
rect 443786 192698 444022 192934
rect 443786 157018 444022 157254
rect 443786 156698 444022 156934
rect 443786 121018 444022 121254
rect 443786 120698 444022 120934
rect 443786 85018 444022 85254
rect 443786 84698 444022 84934
rect 443786 49018 444022 49254
rect 443786 48698 444022 48934
rect 443786 13018 444022 13254
rect 443786 12698 444022 12934
rect 425786 -7022 426022 -6786
rect 425786 -7342 426022 -7106
rect 450986 560218 451222 560454
rect 450986 559898 451222 560134
rect 450986 524218 451222 524454
rect 450986 523898 451222 524134
rect 450986 488218 451222 488454
rect 450986 487898 451222 488134
rect 450986 452218 451222 452454
rect 450986 451898 451222 452134
rect 450986 416218 451222 416454
rect 450986 415898 451222 416134
rect 450986 380218 451222 380454
rect 450986 379898 451222 380134
rect 450986 344218 451222 344454
rect 450986 343898 451222 344134
rect 450986 308218 451222 308454
rect 450986 307898 451222 308134
rect 450986 272218 451222 272454
rect 450986 271898 451222 272134
rect 450986 236218 451222 236454
rect 450986 235898 451222 236134
rect 450986 200218 451222 200454
rect 450986 199898 451222 200134
rect 450986 164218 451222 164454
rect 450986 163898 451222 164134
rect 454586 671818 454822 672054
rect 454586 671498 454822 671734
rect 454586 635818 454822 636054
rect 454586 635498 454822 635734
rect 454586 599818 454822 600054
rect 454586 599498 454822 599734
rect 454586 563818 454822 564054
rect 454586 563498 454822 563734
rect 454586 527818 454822 528054
rect 454586 527498 454822 527734
rect 454586 491818 454822 492054
rect 454586 491498 454822 491734
rect 454586 455818 454822 456054
rect 454586 455498 454822 455734
rect 454586 419818 454822 420054
rect 454586 419498 454822 419734
rect 454586 383818 454822 384054
rect 454586 383498 454822 383734
rect 454586 347818 454822 348054
rect 454586 347498 454822 347734
rect 454586 311818 454822 312054
rect 454586 311498 454822 311734
rect 454586 275818 454822 276054
rect 454586 275498 454822 275734
rect 454586 239818 454822 240054
rect 454586 239498 454822 239734
rect 454586 203818 454822 204054
rect 454586 203498 454822 203734
rect 454586 167818 454822 168054
rect 454586 167498 454822 167734
rect 450986 128218 451222 128454
rect 450986 127898 451222 128134
rect 450986 92218 451222 92454
rect 450986 91898 451222 92134
rect 454586 131818 454822 132054
rect 454586 131498 454822 131734
rect 454586 95818 454822 96054
rect 454586 95498 454822 95734
rect 450986 56218 451222 56454
rect 450986 55898 451222 56134
rect 454586 59818 454822 60054
rect 454586 59498 454822 59734
rect 450986 20218 451222 20454
rect 450986 19898 451222 20134
rect 450986 -1502 451222 -1266
rect 450986 -1822 451222 -1586
rect 454586 23818 454822 24054
rect 454586 23498 454822 23734
rect 454586 -3342 454822 -3106
rect 454586 -3662 454822 -3426
rect 458186 675418 458422 675654
rect 458186 675098 458422 675334
rect 458186 639418 458422 639654
rect 458186 639098 458422 639334
rect 458186 603418 458422 603654
rect 458186 603098 458422 603334
rect 458186 567418 458422 567654
rect 458186 567098 458422 567334
rect 458186 531418 458422 531654
rect 458186 531098 458422 531334
rect 458186 495418 458422 495654
rect 458186 495098 458422 495334
rect 458186 459418 458422 459654
rect 458186 459098 458422 459334
rect 458186 423418 458422 423654
rect 458186 423098 458422 423334
rect 458186 387418 458422 387654
rect 458186 387098 458422 387334
rect 458186 351418 458422 351654
rect 458186 351098 458422 351334
rect 458186 315418 458422 315654
rect 458186 315098 458422 315334
rect 458186 279418 458422 279654
rect 458186 279098 458422 279334
rect 458186 243418 458422 243654
rect 458186 243098 458422 243334
rect 458186 207418 458422 207654
rect 458186 207098 458422 207334
rect 458186 171418 458422 171654
rect 458186 171098 458422 171334
rect 458186 135418 458422 135654
rect 458186 135098 458422 135334
rect 458186 99418 458422 99654
rect 458186 99098 458422 99334
rect 458186 63418 458422 63654
rect 458186 63098 458422 63334
rect 458186 27418 458422 27654
rect 458186 27098 458422 27334
rect 458186 -5182 458422 -4946
rect 458186 -5502 458422 -5266
rect 479786 710122 480022 710358
rect 479786 709802 480022 710038
rect 476186 708282 476422 708518
rect 476186 707962 476422 708198
rect 472586 706442 472822 706678
rect 472586 706122 472822 706358
rect 461786 679018 462022 679254
rect 461786 678698 462022 678934
rect 461786 643018 462022 643254
rect 461786 642698 462022 642934
rect 461786 607018 462022 607254
rect 461786 606698 462022 606934
rect 461786 571018 462022 571254
rect 461786 570698 462022 570934
rect 461786 535018 462022 535254
rect 461786 534698 462022 534934
rect 461786 499018 462022 499254
rect 461786 498698 462022 498934
rect 461786 463018 462022 463254
rect 461786 462698 462022 462934
rect 461786 427018 462022 427254
rect 461786 426698 462022 426934
rect 461786 391018 462022 391254
rect 461786 390698 462022 390934
rect 461786 355018 462022 355254
rect 461786 354698 462022 354934
rect 461786 319018 462022 319254
rect 461786 318698 462022 318934
rect 461786 283018 462022 283254
rect 461786 282698 462022 282934
rect 461786 247018 462022 247254
rect 461786 246698 462022 246934
rect 461786 211018 462022 211254
rect 461786 210698 462022 210934
rect 461786 175018 462022 175254
rect 461786 174698 462022 174934
rect 461786 139018 462022 139254
rect 461786 138698 462022 138934
rect 461786 103018 462022 103254
rect 461786 102698 462022 102934
rect 461786 67018 462022 67254
rect 461786 66698 462022 66934
rect 461786 31018 462022 31254
rect 461786 30698 462022 30934
rect 443786 -6102 444022 -5866
rect 443786 -6422 444022 -6186
rect 468986 704602 469222 704838
rect 468986 704282 469222 704518
rect 468986 686218 469222 686454
rect 468986 685898 469222 686134
rect 468986 650218 469222 650454
rect 468986 649898 469222 650134
rect 468986 614218 469222 614454
rect 468986 613898 469222 614134
rect 468986 578218 469222 578454
rect 468986 577898 469222 578134
rect 468986 542218 469222 542454
rect 468986 541898 469222 542134
rect 468986 506218 469222 506454
rect 468986 505898 469222 506134
rect 468986 470218 469222 470454
rect 468986 469898 469222 470134
rect 468986 434218 469222 434454
rect 468986 433898 469222 434134
rect 468986 398218 469222 398454
rect 468986 397898 469222 398134
rect 468986 362218 469222 362454
rect 468986 361898 469222 362134
rect 468986 326218 469222 326454
rect 468986 325898 469222 326134
rect 468986 290218 469222 290454
rect 468986 289898 469222 290134
rect 468986 254218 469222 254454
rect 468986 253898 469222 254134
rect 468986 218218 469222 218454
rect 468986 217898 469222 218134
rect 468986 182218 469222 182454
rect 468986 181898 469222 182134
rect 468986 146218 469222 146454
rect 468986 145898 469222 146134
rect 468986 110218 469222 110454
rect 468986 109898 469222 110134
rect 468986 74218 469222 74454
rect 468986 73898 469222 74134
rect 468986 38218 469222 38454
rect 468986 37898 469222 38134
rect 468986 2218 469222 2454
rect 468986 1898 469222 2134
rect 468986 -582 469222 -346
rect 468986 -902 469222 -666
rect 472586 689818 472822 690054
rect 472586 689498 472822 689734
rect 472586 653818 472822 654054
rect 472586 653498 472822 653734
rect 472586 617818 472822 618054
rect 472586 617498 472822 617734
rect 472586 581818 472822 582054
rect 472586 581498 472822 581734
rect 472586 545818 472822 546054
rect 472586 545498 472822 545734
rect 472586 509818 472822 510054
rect 472586 509498 472822 509734
rect 472586 473818 472822 474054
rect 472586 473498 472822 473734
rect 472586 437818 472822 438054
rect 472586 437498 472822 437734
rect 472586 401818 472822 402054
rect 472586 401498 472822 401734
rect 472586 365818 472822 366054
rect 472586 365498 472822 365734
rect 472586 329818 472822 330054
rect 472586 329498 472822 329734
rect 472586 293818 472822 294054
rect 472586 293498 472822 293734
rect 472586 257818 472822 258054
rect 472586 257498 472822 257734
rect 472586 221818 472822 222054
rect 472586 221498 472822 221734
rect 472586 185818 472822 186054
rect 472586 185498 472822 185734
rect 472586 149818 472822 150054
rect 472586 149498 472822 149734
rect 472586 113818 472822 114054
rect 472586 113498 472822 113734
rect 476186 693418 476422 693654
rect 476186 693098 476422 693334
rect 476186 657418 476422 657654
rect 476186 657098 476422 657334
rect 476186 621418 476422 621654
rect 476186 621098 476422 621334
rect 476186 585418 476422 585654
rect 476186 585098 476422 585334
rect 476186 549418 476422 549654
rect 476186 549098 476422 549334
rect 476186 513418 476422 513654
rect 476186 513098 476422 513334
rect 476186 477418 476422 477654
rect 476186 477098 476422 477334
rect 476186 441418 476422 441654
rect 476186 441098 476422 441334
rect 476186 405418 476422 405654
rect 476186 405098 476422 405334
rect 476186 369418 476422 369654
rect 476186 369098 476422 369334
rect 476186 333418 476422 333654
rect 476186 333098 476422 333334
rect 476186 297418 476422 297654
rect 476186 297098 476422 297334
rect 476186 261418 476422 261654
rect 476186 261098 476422 261334
rect 476186 225418 476422 225654
rect 476186 225098 476422 225334
rect 476186 189418 476422 189654
rect 476186 189098 476422 189334
rect 476186 153418 476422 153654
rect 476186 153098 476422 153334
rect 476186 117418 476422 117654
rect 476186 117098 476422 117334
rect 472586 77818 472822 78054
rect 472586 77498 472822 77734
rect 472586 41818 472822 42054
rect 472586 41498 472822 41734
rect 472586 5818 472822 6054
rect 472586 5498 472822 5734
rect 472586 -2422 472822 -2186
rect 472586 -2742 472822 -2506
rect 476186 81418 476422 81654
rect 476186 81098 476422 81334
rect 476186 45418 476422 45654
rect 476186 45098 476422 45334
rect 476186 9418 476422 9654
rect 476186 9098 476422 9334
rect 476186 -4262 476422 -4026
rect 476186 -4582 476422 -4346
rect 497786 711042 498022 711278
rect 497786 710722 498022 710958
rect 494186 709202 494422 709438
rect 494186 708882 494422 709118
rect 490586 707362 490822 707598
rect 490586 707042 490822 707278
rect 479786 697018 480022 697254
rect 479786 696698 480022 696934
rect 479786 661018 480022 661254
rect 479786 660698 480022 660934
rect 479786 625018 480022 625254
rect 479786 624698 480022 624934
rect 479786 589018 480022 589254
rect 479786 588698 480022 588934
rect 479786 553018 480022 553254
rect 479786 552698 480022 552934
rect 479786 517018 480022 517254
rect 479786 516698 480022 516934
rect 479786 481018 480022 481254
rect 479786 480698 480022 480934
rect 479786 445018 480022 445254
rect 479786 444698 480022 444934
rect 479786 409018 480022 409254
rect 479786 408698 480022 408934
rect 479786 373018 480022 373254
rect 479786 372698 480022 372934
rect 479786 337018 480022 337254
rect 479786 336698 480022 336934
rect 479786 301018 480022 301254
rect 479786 300698 480022 300934
rect 479786 265018 480022 265254
rect 479786 264698 480022 264934
rect 479786 229018 480022 229254
rect 479786 228698 480022 228934
rect 479786 193018 480022 193254
rect 479786 192698 480022 192934
rect 479786 157018 480022 157254
rect 479786 156698 480022 156934
rect 479786 121018 480022 121254
rect 479786 120698 480022 120934
rect 479786 85018 480022 85254
rect 479786 84698 480022 84934
rect 479786 49018 480022 49254
rect 479786 48698 480022 48934
rect 479786 13018 480022 13254
rect 479786 12698 480022 12934
rect 461786 -7022 462022 -6786
rect 461786 -7342 462022 -7106
rect 486986 705522 487222 705758
rect 486986 705202 487222 705438
rect 486986 668218 487222 668454
rect 486986 667898 487222 668134
rect 486986 632218 487222 632454
rect 486986 631898 487222 632134
rect 486986 596218 487222 596454
rect 486986 595898 487222 596134
rect 486986 560218 487222 560454
rect 486986 559898 487222 560134
rect 486986 524218 487222 524454
rect 486986 523898 487222 524134
rect 486986 488218 487222 488454
rect 486986 487898 487222 488134
rect 486986 452218 487222 452454
rect 486986 451898 487222 452134
rect 486986 416218 487222 416454
rect 486986 415898 487222 416134
rect 486986 380218 487222 380454
rect 486986 379898 487222 380134
rect 486986 344218 487222 344454
rect 486986 343898 487222 344134
rect 486986 308218 487222 308454
rect 486986 307898 487222 308134
rect 486986 272218 487222 272454
rect 486986 271898 487222 272134
rect 486986 236218 487222 236454
rect 486986 235898 487222 236134
rect 486986 200218 487222 200454
rect 486986 199898 487222 200134
rect 486986 164218 487222 164454
rect 486986 163898 487222 164134
rect 486986 128218 487222 128454
rect 486986 127898 487222 128134
rect 486986 92218 487222 92454
rect 486986 91898 487222 92134
rect 486986 56218 487222 56454
rect 486986 55898 487222 56134
rect 486986 20218 487222 20454
rect 486986 19898 487222 20134
rect 486986 -1502 487222 -1266
rect 486986 -1822 487222 -1586
rect 490586 671818 490822 672054
rect 490586 671498 490822 671734
rect 490586 635818 490822 636054
rect 490586 635498 490822 635734
rect 490586 599818 490822 600054
rect 490586 599498 490822 599734
rect 490586 563818 490822 564054
rect 490586 563498 490822 563734
rect 490586 527818 490822 528054
rect 490586 527498 490822 527734
rect 490586 491818 490822 492054
rect 490586 491498 490822 491734
rect 490586 455818 490822 456054
rect 490586 455498 490822 455734
rect 490586 419818 490822 420054
rect 490586 419498 490822 419734
rect 490586 383818 490822 384054
rect 490586 383498 490822 383734
rect 490586 347818 490822 348054
rect 490586 347498 490822 347734
rect 490586 311818 490822 312054
rect 490586 311498 490822 311734
rect 490586 275818 490822 276054
rect 490586 275498 490822 275734
rect 490586 239818 490822 240054
rect 490586 239498 490822 239734
rect 490586 203818 490822 204054
rect 490586 203498 490822 203734
rect 490586 167818 490822 168054
rect 490586 167498 490822 167734
rect 490586 131818 490822 132054
rect 490586 131498 490822 131734
rect 490586 95818 490822 96054
rect 490586 95498 490822 95734
rect 490586 59818 490822 60054
rect 490586 59498 490822 59734
rect 490586 23818 490822 24054
rect 490586 23498 490822 23734
rect 490586 -3342 490822 -3106
rect 490586 -3662 490822 -3426
rect 494186 675418 494422 675654
rect 494186 675098 494422 675334
rect 494186 639418 494422 639654
rect 494186 639098 494422 639334
rect 494186 603418 494422 603654
rect 494186 603098 494422 603334
rect 494186 567418 494422 567654
rect 494186 567098 494422 567334
rect 494186 531418 494422 531654
rect 494186 531098 494422 531334
rect 494186 495418 494422 495654
rect 494186 495098 494422 495334
rect 494186 459418 494422 459654
rect 494186 459098 494422 459334
rect 494186 423418 494422 423654
rect 494186 423098 494422 423334
rect 494186 387418 494422 387654
rect 494186 387098 494422 387334
rect 494186 351418 494422 351654
rect 494186 351098 494422 351334
rect 494186 315418 494422 315654
rect 494186 315098 494422 315334
rect 494186 279418 494422 279654
rect 494186 279098 494422 279334
rect 494186 243418 494422 243654
rect 494186 243098 494422 243334
rect 494186 207418 494422 207654
rect 494186 207098 494422 207334
rect 494186 171418 494422 171654
rect 494186 171098 494422 171334
rect 494186 135418 494422 135654
rect 494186 135098 494422 135334
rect 494186 99418 494422 99654
rect 494186 99098 494422 99334
rect 494186 63418 494422 63654
rect 494186 63098 494422 63334
rect 494186 27418 494422 27654
rect 494186 27098 494422 27334
rect 494186 -5182 494422 -4946
rect 494186 -5502 494422 -5266
rect 515786 710122 516022 710358
rect 515786 709802 516022 710038
rect 512186 708282 512422 708518
rect 512186 707962 512422 708198
rect 508586 706442 508822 706678
rect 508586 706122 508822 706358
rect 497786 679018 498022 679254
rect 497786 678698 498022 678934
rect 497786 643018 498022 643254
rect 497786 642698 498022 642934
rect 497786 607018 498022 607254
rect 497786 606698 498022 606934
rect 497786 571018 498022 571254
rect 497786 570698 498022 570934
rect 497786 535018 498022 535254
rect 497786 534698 498022 534934
rect 497786 499018 498022 499254
rect 497786 498698 498022 498934
rect 497786 463018 498022 463254
rect 497786 462698 498022 462934
rect 497786 427018 498022 427254
rect 497786 426698 498022 426934
rect 497786 391018 498022 391254
rect 497786 390698 498022 390934
rect 497786 355018 498022 355254
rect 497786 354698 498022 354934
rect 497786 319018 498022 319254
rect 497786 318698 498022 318934
rect 497786 283018 498022 283254
rect 497786 282698 498022 282934
rect 497786 247018 498022 247254
rect 497786 246698 498022 246934
rect 497786 211018 498022 211254
rect 497786 210698 498022 210934
rect 497786 175018 498022 175254
rect 497786 174698 498022 174934
rect 497786 139018 498022 139254
rect 497786 138698 498022 138934
rect 497786 103018 498022 103254
rect 497786 102698 498022 102934
rect 497786 67018 498022 67254
rect 497786 66698 498022 66934
rect 497786 31018 498022 31254
rect 497786 30698 498022 30934
rect 479786 -6102 480022 -5866
rect 479786 -6422 480022 -6186
rect 504986 704602 505222 704838
rect 504986 704282 505222 704518
rect 504986 686218 505222 686454
rect 504986 685898 505222 686134
rect 504986 650218 505222 650454
rect 504986 649898 505222 650134
rect 504986 614218 505222 614454
rect 504986 613898 505222 614134
rect 504986 578218 505222 578454
rect 504986 577898 505222 578134
rect 504986 542218 505222 542454
rect 504986 541898 505222 542134
rect 504986 506218 505222 506454
rect 504986 505898 505222 506134
rect 504986 470218 505222 470454
rect 504986 469898 505222 470134
rect 504986 434218 505222 434454
rect 504986 433898 505222 434134
rect 504986 398218 505222 398454
rect 504986 397898 505222 398134
rect 504986 362218 505222 362454
rect 504986 361898 505222 362134
rect 504986 326218 505222 326454
rect 504986 325898 505222 326134
rect 504986 290218 505222 290454
rect 504986 289898 505222 290134
rect 504986 254218 505222 254454
rect 504986 253898 505222 254134
rect 504986 218218 505222 218454
rect 504986 217898 505222 218134
rect 504986 182218 505222 182454
rect 504986 181898 505222 182134
rect 504986 146218 505222 146454
rect 504986 145898 505222 146134
rect 504986 110218 505222 110454
rect 504986 109898 505222 110134
rect 504986 74218 505222 74454
rect 504986 73898 505222 74134
rect 504986 38218 505222 38454
rect 504986 37898 505222 38134
rect 504986 2218 505222 2454
rect 504986 1898 505222 2134
rect 504986 -582 505222 -346
rect 504986 -902 505222 -666
rect 508586 689818 508822 690054
rect 508586 689498 508822 689734
rect 508586 653818 508822 654054
rect 508586 653498 508822 653734
rect 508586 617818 508822 618054
rect 508586 617498 508822 617734
rect 508586 581818 508822 582054
rect 508586 581498 508822 581734
rect 508586 545818 508822 546054
rect 508586 545498 508822 545734
rect 508586 509818 508822 510054
rect 508586 509498 508822 509734
rect 508586 473818 508822 474054
rect 508586 473498 508822 473734
rect 508586 437818 508822 438054
rect 508586 437498 508822 437734
rect 508586 401818 508822 402054
rect 508586 401498 508822 401734
rect 508586 365818 508822 366054
rect 508586 365498 508822 365734
rect 508586 329818 508822 330054
rect 508586 329498 508822 329734
rect 508586 293818 508822 294054
rect 508586 293498 508822 293734
rect 508586 257818 508822 258054
rect 508586 257498 508822 257734
rect 508586 221818 508822 222054
rect 508586 221498 508822 221734
rect 508586 185818 508822 186054
rect 508586 185498 508822 185734
rect 508586 149818 508822 150054
rect 508586 149498 508822 149734
rect 508586 113818 508822 114054
rect 508586 113498 508822 113734
rect 508586 77818 508822 78054
rect 508586 77498 508822 77734
rect 508586 41818 508822 42054
rect 508586 41498 508822 41734
rect 508586 5818 508822 6054
rect 508586 5498 508822 5734
rect 508586 -2422 508822 -2186
rect 508586 -2742 508822 -2506
rect 512186 693418 512422 693654
rect 512186 693098 512422 693334
rect 512186 657418 512422 657654
rect 512186 657098 512422 657334
rect 512186 621418 512422 621654
rect 512186 621098 512422 621334
rect 512186 585418 512422 585654
rect 512186 585098 512422 585334
rect 512186 549418 512422 549654
rect 512186 549098 512422 549334
rect 512186 513418 512422 513654
rect 512186 513098 512422 513334
rect 512186 477418 512422 477654
rect 512186 477098 512422 477334
rect 512186 441418 512422 441654
rect 512186 441098 512422 441334
rect 512186 405418 512422 405654
rect 512186 405098 512422 405334
rect 512186 369418 512422 369654
rect 512186 369098 512422 369334
rect 512186 333418 512422 333654
rect 512186 333098 512422 333334
rect 512186 297418 512422 297654
rect 512186 297098 512422 297334
rect 512186 261418 512422 261654
rect 512186 261098 512422 261334
rect 512186 225418 512422 225654
rect 512186 225098 512422 225334
rect 512186 189418 512422 189654
rect 512186 189098 512422 189334
rect 512186 153418 512422 153654
rect 512186 153098 512422 153334
rect 512186 117418 512422 117654
rect 512186 117098 512422 117334
rect 512186 81418 512422 81654
rect 512186 81098 512422 81334
rect 512186 45418 512422 45654
rect 512186 45098 512422 45334
rect 512186 9418 512422 9654
rect 512186 9098 512422 9334
rect 512186 -4262 512422 -4026
rect 512186 -4582 512422 -4346
rect 533786 711042 534022 711278
rect 533786 710722 534022 710958
rect 530186 709202 530422 709438
rect 530186 708882 530422 709118
rect 526586 707362 526822 707598
rect 526586 707042 526822 707278
rect 515786 697018 516022 697254
rect 515786 696698 516022 696934
rect 515786 661018 516022 661254
rect 515786 660698 516022 660934
rect 515786 625018 516022 625254
rect 515786 624698 516022 624934
rect 515786 589018 516022 589254
rect 515786 588698 516022 588934
rect 515786 553018 516022 553254
rect 515786 552698 516022 552934
rect 515786 517018 516022 517254
rect 515786 516698 516022 516934
rect 515786 481018 516022 481254
rect 515786 480698 516022 480934
rect 515786 445018 516022 445254
rect 515786 444698 516022 444934
rect 515786 409018 516022 409254
rect 515786 408698 516022 408934
rect 515786 373018 516022 373254
rect 515786 372698 516022 372934
rect 515786 337018 516022 337254
rect 515786 336698 516022 336934
rect 515786 301018 516022 301254
rect 515786 300698 516022 300934
rect 515786 265018 516022 265254
rect 515786 264698 516022 264934
rect 515786 229018 516022 229254
rect 515786 228698 516022 228934
rect 515786 193018 516022 193254
rect 515786 192698 516022 192934
rect 515786 157018 516022 157254
rect 515786 156698 516022 156934
rect 515786 121018 516022 121254
rect 515786 120698 516022 120934
rect 515786 85018 516022 85254
rect 515786 84698 516022 84934
rect 515786 49018 516022 49254
rect 515786 48698 516022 48934
rect 515786 13018 516022 13254
rect 515786 12698 516022 12934
rect 497786 -7022 498022 -6786
rect 497786 -7342 498022 -7106
rect 522986 705522 523222 705758
rect 522986 705202 523222 705438
rect 522986 668218 523222 668454
rect 522986 667898 523222 668134
rect 522986 632218 523222 632454
rect 522986 631898 523222 632134
rect 522986 596218 523222 596454
rect 522986 595898 523222 596134
rect 522986 560218 523222 560454
rect 522986 559898 523222 560134
rect 522986 524218 523222 524454
rect 522986 523898 523222 524134
rect 522986 488218 523222 488454
rect 522986 487898 523222 488134
rect 522986 452218 523222 452454
rect 522986 451898 523222 452134
rect 522986 416218 523222 416454
rect 522986 415898 523222 416134
rect 522986 380218 523222 380454
rect 522986 379898 523222 380134
rect 522986 344218 523222 344454
rect 522986 343898 523222 344134
rect 522986 308218 523222 308454
rect 522986 307898 523222 308134
rect 522986 272218 523222 272454
rect 522986 271898 523222 272134
rect 522986 236218 523222 236454
rect 522986 235898 523222 236134
rect 522986 200218 523222 200454
rect 522986 199898 523222 200134
rect 522986 164218 523222 164454
rect 522986 163898 523222 164134
rect 522986 128218 523222 128454
rect 522986 127898 523222 128134
rect 522986 92218 523222 92454
rect 522986 91898 523222 92134
rect 522986 56218 523222 56454
rect 522986 55898 523222 56134
rect 522986 20218 523222 20454
rect 522986 19898 523222 20134
rect 522986 -1502 523222 -1266
rect 522986 -1822 523222 -1586
rect 526586 671818 526822 672054
rect 526586 671498 526822 671734
rect 526586 635818 526822 636054
rect 526586 635498 526822 635734
rect 526586 599818 526822 600054
rect 526586 599498 526822 599734
rect 526586 563818 526822 564054
rect 526586 563498 526822 563734
rect 526586 527818 526822 528054
rect 526586 527498 526822 527734
rect 526586 491818 526822 492054
rect 526586 491498 526822 491734
rect 526586 455818 526822 456054
rect 526586 455498 526822 455734
rect 526586 419818 526822 420054
rect 526586 419498 526822 419734
rect 526586 383818 526822 384054
rect 526586 383498 526822 383734
rect 526586 347818 526822 348054
rect 526586 347498 526822 347734
rect 526586 311818 526822 312054
rect 526586 311498 526822 311734
rect 526586 275818 526822 276054
rect 526586 275498 526822 275734
rect 526586 239818 526822 240054
rect 526586 239498 526822 239734
rect 526586 203818 526822 204054
rect 526586 203498 526822 203734
rect 526586 167818 526822 168054
rect 526586 167498 526822 167734
rect 526586 131818 526822 132054
rect 526586 131498 526822 131734
rect 526586 95818 526822 96054
rect 526586 95498 526822 95734
rect 526586 59818 526822 60054
rect 526586 59498 526822 59734
rect 526586 23818 526822 24054
rect 526586 23498 526822 23734
rect 526586 -3342 526822 -3106
rect 526586 -3662 526822 -3426
rect 530186 675418 530422 675654
rect 530186 675098 530422 675334
rect 530186 639418 530422 639654
rect 530186 639098 530422 639334
rect 530186 603418 530422 603654
rect 530186 603098 530422 603334
rect 530186 567418 530422 567654
rect 530186 567098 530422 567334
rect 530186 531418 530422 531654
rect 530186 531098 530422 531334
rect 530186 495418 530422 495654
rect 530186 495098 530422 495334
rect 530186 459418 530422 459654
rect 530186 459098 530422 459334
rect 530186 423418 530422 423654
rect 530186 423098 530422 423334
rect 530186 387418 530422 387654
rect 530186 387098 530422 387334
rect 530186 351418 530422 351654
rect 530186 351098 530422 351334
rect 530186 315418 530422 315654
rect 530186 315098 530422 315334
rect 530186 279418 530422 279654
rect 530186 279098 530422 279334
rect 530186 243418 530422 243654
rect 530186 243098 530422 243334
rect 530186 207418 530422 207654
rect 530186 207098 530422 207334
rect 530186 171418 530422 171654
rect 530186 171098 530422 171334
rect 530186 135418 530422 135654
rect 530186 135098 530422 135334
rect 530186 99418 530422 99654
rect 530186 99098 530422 99334
rect 530186 63418 530422 63654
rect 530186 63098 530422 63334
rect 530186 27418 530422 27654
rect 530186 27098 530422 27334
rect 530186 -5182 530422 -4946
rect 530186 -5502 530422 -5266
rect 551786 710122 552022 710358
rect 551786 709802 552022 710038
rect 548186 708282 548422 708518
rect 548186 707962 548422 708198
rect 544586 706442 544822 706678
rect 544586 706122 544822 706358
rect 533786 679018 534022 679254
rect 533786 678698 534022 678934
rect 533786 643018 534022 643254
rect 533786 642698 534022 642934
rect 533786 607018 534022 607254
rect 533786 606698 534022 606934
rect 533786 571018 534022 571254
rect 533786 570698 534022 570934
rect 533786 535018 534022 535254
rect 533786 534698 534022 534934
rect 533786 499018 534022 499254
rect 533786 498698 534022 498934
rect 533786 463018 534022 463254
rect 533786 462698 534022 462934
rect 533786 427018 534022 427254
rect 533786 426698 534022 426934
rect 533786 391018 534022 391254
rect 533786 390698 534022 390934
rect 533786 355018 534022 355254
rect 533786 354698 534022 354934
rect 533786 319018 534022 319254
rect 533786 318698 534022 318934
rect 533786 283018 534022 283254
rect 533786 282698 534022 282934
rect 533786 247018 534022 247254
rect 533786 246698 534022 246934
rect 533786 211018 534022 211254
rect 533786 210698 534022 210934
rect 533786 175018 534022 175254
rect 533786 174698 534022 174934
rect 533786 139018 534022 139254
rect 533786 138698 534022 138934
rect 533786 103018 534022 103254
rect 533786 102698 534022 102934
rect 533786 67018 534022 67254
rect 533786 66698 534022 66934
rect 533786 31018 534022 31254
rect 533786 30698 534022 30934
rect 515786 -6102 516022 -5866
rect 515786 -6422 516022 -6186
rect 540986 704602 541222 704838
rect 540986 704282 541222 704518
rect 540986 686218 541222 686454
rect 540986 685898 541222 686134
rect 540986 650218 541222 650454
rect 540986 649898 541222 650134
rect 540986 614218 541222 614454
rect 540986 613898 541222 614134
rect 540986 578218 541222 578454
rect 540986 577898 541222 578134
rect 540986 542218 541222 542454
rect 540986 541898 541222 542134
rect 540986 506218 541222 506454
rect 540986 505898 541222 506134
rect 540986 470218 541222 470454
rect 540986 469898 541222 470134
rect 540986 434218 541222 434454
rect 540986 433898 541222 434134
rect 540986 398218 541222 398454
rect 540986 397898 541222 398134
rect 540986 362218 541222 362454
rect 540986 361898 541222 362134
rect 540986 326218 541222 326454
rect 540986 325898 541222 326134
rect 540986 290218 541222 290454
rect 540986 289898 541222 290134
rect 540986 254218 541222 254454
rect 540986 253898 541222 254134
rect 540986 218218 541222 218454
rect 540986 217898 541222 218134
rect 540986 182218 541222 182454
rect 540986 181898 541222 182134
rect 540986 146218 541222 146454
rect 540986 145898 541222 146134
rect 540986 110218 541222 110454
rect 540986 109898 541222 110134
rect 540986 74218 541222 74454
rect 540986 73898 541222 74134
rect 540986 38218 541222 38454
rect 540986 37898 541222 38134
rect 540986 2218 541222 2454
rect 540986 1898 541222 2134
rect 540986 -582 541222 -346
rect 540986 -902 541222 -666
rect 544586 689818 544822 690054
rect 544586 689498 544822 689734
rect 544586 653818 544822 654054
rect 544586 653498 544822 653734
rect 544586 617818 544822 618054
rect 544586 617498 544822 617734
rect 544586 581818 544822 582054
rect 544586 581498 544822 581734
rect 544586 545818 544822 546054
rect 544586 545498 544822 545734
rect 544586 509818 544822 510054
rect 544586 509498 544822 509734
rect 544586 473818 544822 474054
rect 544586 473498 544822 473734
rect 544586 437818 544822 438054
rect 544586 437498 544822 437734
rect 544586 401818 544822 402054
rect 544586 401498 544822 401734
rect 544586 365818 544822 366054
rect 544586 365498 544822 365734
rect 544586 329818 544822 330054
rect 544586 329498 544822 329734
rect 544586 293818 544822 294054
rect 544586 293498 544822 293734
rect 544586 257818 544822 258054
rect 544586 257498 544822 257734
rect 544586 221818 544822 222054
rect 544586 221498 544822 221734
rect 544586 185818 544822 186054
rect 544586 185498 544822 185734
rect 544586 149818 544822 150054
rect 544586 149498 544822 149734
rect 544586 113818 544822 114054
rect 544586 113498 544822 113734
rect 544586 77818 544822 78054
rect 544586 77498 544822 77734
rect 544586 41818 544822 42054
rect 544586 41498 544822 41734
rect 544586 5818 544822 6054
rect 544586 5498 544822 5734
rect 544586 -2422 544822 -2186
rect 544586 -2742 544822 -2506
rect 548186 693418 548422 693654
rect 548186 693098 548422 693334
rect 548186 657418 548422 657654
rect 548186 657098 548422 657334
rect 548186 621418 548422 621654
rect 548186 621098 548422 621334
rect 548186 585418 548422 585654
rect 548186 585098 548422 585334
rect 548186 549418 548422 549654
rect 548186 549098 548422 549334
rect 548186 513418 548422 513654
rect 548186 513098 548422 513334
rect 548186 477418 548422 477654
rect 548186 477098 548422 477334
rect 548186 441418 548422 441654
rect 548186 441098 548422 441334
rect 548186 405418 548422 405654
rect 548186 405098 548422 405334
rect 548186 369418 548422 369654
rect 548186 369098 548422 369334
rect 548186 333418 548422 333654
rect 548186 333098 548422 333334
rect 548186 297418 548422 297654
rect 548186 297098 548422 297334
rect 548186 261418 548422 261654
rect 548186 261098 548422 261334
rect 548186 225418 548422 225654
rect 548186 225098 548422 225334
rect 548186 189418 548422 189654
rect 548186 189098 548422 189334
rect 548186 153418 548422 153654
rect 548186 153098 548422 153334
rect 548186 117418 548422 117654
rect 548186 117098 548422 117334
rect 548186 81418 548422 81654
rect 548186 81098 548422 81334
rect 548186 45418 548422 45654
rect 548186 45098 548422 45334
rect 548186 9418 548422 9654
rect 548186 9098 548422 9334
rect 548186 -4262 548422 -4026
rect 548186 -4582 548422 -4346
rect 569786 711042 570022 711278
rect 569786 710722 570022 710958
rect 566186 709202 566422 709438
rect 566186 708882 566422 709118
rect 562586 707362 562822 707598
rect 562586 707042 562822 707278
rect 551786 697018 552022 697254
rect 551786 696698 552022 696934
rect 551786 661018 552022 661254
rect 551786 660698 552022 660934
rect 551786 625018 552022 625254
rect 551786 624698 552022 624934
rect 551786 589018 552022 589254
rect 551786 588698 552022 588934
rect 551786 553018 552022 553254
rect 551786 552698 552022 552934
rect 551786 517018 552022 517254
rect 551786 516698 552022 516934
rect 551786 481018 552022 481254
rect 551786 480698 552022 480934
rect 551786 445018 552022 445254
rect 551786 444698 552022 444934
rect 551786 409018 552022 409254
rect 551786 408698 552022 408934
rect 551786 373018 552022 373254
rect 551786 372698 552022 372934
rect 551786 337018 552022 337254
rect 551786 336698 552022 336934
rect 551786 301018 552022 301254
rect 551786 300698 552022 300934
rect 551786 265018 552022 265254
rect 551786 264698 552022 264934
rect 551786 229018 552022 229254
rect 551786 228698 552022 228934
rect 551786 193018 552022 193254
rect 551786 192698 552022 192934
rect 551786 157018 552022 157254
rect 551786 156698 552022 156934
rect 551786 121018 552022 121254
rect 551786 120698 552022 120934
rect 551786 85018 552022 85254
rect 551786 84698 552022 84934
rect 551786 49018 552022 49254
rect 551786 48698 552022 48934
rect 551786 13018 552022 13254
rect 551786 12698 552022 12934
rect 533786 -7022 534022 -6786
rect 533786 -7342 534022 -7106
rect 558986 705522 559222 705758
rect 558986 705202 559222 705438
rect 558986 668218 559222 668454
rect 558986 667898 559222 668134
rect 558986 632218 559222 632454
rect 558986 631898 559222 632134
rect 558986 596218 559222 596454
rect 558986 595898 559222 596134
rect 558986 560218 559222 560454
rect 558986 559898 559222 560134
rect 558986 524218 559222 524454
rect 558986 523898 559222 524134
rect 558986 488218 559222 488454
rect 558986 487898 559222 488134
rect 558986 452218 559222 452454
rect 558986 451898 559222 452134
rect 558986 416218 559222 416454
rect 558986 415898 559222 416134
rect 558986 380218 559222 380454
rect 558986 379898 559222 380134
rect 558986 344218 559222 344454
rect 558986 343898 559222 344134
rect 558986 308218 559222 308454
rect 558986 307898 559222 308134
rect 558986 272218 559222 272454
rect 558986 271898 559222 272134
rect 558986 236218 559222 236454
rect 558986 235898 559222 236134
rect 558986 200218 559222 200454
rect 558986 199898 559222 200134
rect 558986 164218 559222 164454
rect 558986 163898 559222 164134
rect 558986 128218 559222 128454
rect 558986 127898 559222 128134
rect 558986 92218 559222 92454
rect 558986 91898 559222 92134
rect 558986 56218 559222 56454
rect 558986 55898 559222 56134
rect 558986 20218 559222 20454
rect 558986 19898 559222 20134
rect 558986 -1502 559222 -1266
rect 558986 -1822 559222 -1586
rect 562586 671818 562822 672054
rect 562586 671498 562822 671734
rect 562586 635818 562822 636054
rect 562586 635498 562822 635734
rect 562586 599818 562822 600054
rect 562586 599498 562822 599734
rect 562586 563818 562822 564054
rect 562586 563498 562822 563734
rect 562586 527818 562822 528054
rect 562586 527498 562822 527734
rect 562586 491818 562822 492054
rect 562586 491498 562822 491734
rect 562586 455818 562822 456054
rect 562586 455498 562822 455734
rect 562586 419818 562822 420054
rect 562586 419498 562822 419734
rect 562586 383818 562822 384054
rect 562586 383498 562822 383734
rect 562586 347818 562822 348054
rect 562586 347498 562822 347734
rect 562586 311818 562822 312054
rect 562586 311498 562822 311734
rect 562586 275818 562822 276054
rect 562586 275498 562822 275734
rect 562586 239818 562822 240054
rect 562586 239498 562822 239734
rect 562586 203818 562822 204054
rect 562586 203498 562822 203734
rect 562586 167818 562822 168054
rect 562586 167498 562822 167734
rect 562586 131818 562822 132054
rect 562586 131498 562822 131734
rect 562586 95818 562822 96054
rect 562586 95498 562822 95734
rect 562586 59818 562822 60054
rect 562586 59498 562822 59734
rect 562586 23818 562822 24054
rect 562586 23498 562822 23734
rect 562586 -3342 562822 -3106
rect 562586 -3662 562822 -3426
rect 566186 675418 566422 675654
rect 566186 675098 566422 675334
rect 566186 639418 566422 639654
rect 566186 639098 566422 639334
rect 566186 603418 566422 603654
rect 566186 603098 566422 603334
rect 566186 567418 566422 567654
rect 566186 567098 566422 567334
rect 566186 531418 566422 531654
rect 566186 531098 566422 531334
rect 566186 495418 566422 495654
rect 566186 495098 566422 495334
rect 566186 459418 566422 459654
rect 566186 459098 566422 459334
rect 566186 423418 566422 423654
rect 566186 423098 566422 423334
rect 566186 387418 566422 387654
rect 566186 387098 566422 387334
rect 566186 351418 566422 351654
rect 566186 351098 566422 351334
rect 566186 315418 566422 315654
rect 566186 315098 566422 315334
rect 566186 279418 566422 279654
rect 566186 279098 566422 279334
rect 566186 243418 566422 243654
rect 566186 243098 566422 243334
rect 566186 207418 566422 207654
rect 566186 207098 566422 207334
rect 566186 171418 566422 171654
rect 566186 171098 566422 171334
rect 566186 135418 566422 135654
rect 566186 135098 566422 135334
rect 566186 99418 566422 99654
rect 566186 99098 566422 99334
rect 566186 63418 566422 63654
rect 566186 63098 566422 63334
rect 566186 27418 566422 27654
rect 566186 27098 566422 27334
rect 566186 -5182 566422 -4946
rect 566186 -5502 566422 -5266
rect 591942 711042 592178 711278
rect 591942 710722 592178 710958
rect 591022 710122 591258 710358
rect 591022 709802 591258 710038
rect 590102 709202 590338 709438
rect 590102 708882 590338 709118
rect 589182 708282 589418 708518
rect 589182 707962 589418 708198
rect 588262 707362 588498 707598
rect 588262 707042 588498 707278
rect 580586 706442 580822 706678
rect 580586 706122 580822 706358
rect 569786 679018 570022 679254
rect 569786 678698 570022 678934
rect 569786 643018 570022 643254
rect 569786 642698 570022 642934
rect 569786 607018 570022 607254
rect 569786 606698 570022 606934
rect 569786 571018 570022 571254
rect 569786 570698 570022 570934
rect 569786 535018 570022 535254
rect 569786 534698 570022 534934
rect 569786 499018 570022 499254
rect 569786 498698 570022 498934
rect 569786 463018 570022 463254
rect 569786 462698 570022 462934
rect 569786 427018 570022 427254
rect 569786 426698 570022 426934
rect 569786 391018 570022 391254
rect 569786 390698 570022 390934
rect 569786 355018 570022 355254
rect 569786 354698 570022 354934
rect 569786 319018 570022 319254
rect 569786 318698 570022 318934
rect 569786 283018 570022 283254
rect 569786 282698 570022 282934
rect 569786 247018 570022 247254
rect 569786 246698 570022 246934
rect 569786 211018 570022 211254
rect 569786 210698 570022 210934
rect 569786 175018 570022 175254
rect 569786 174698 570022 174934
rect 569786 139018 570022 139254
rect 569786 138698 570022 138934
rect 569786 103018 570022 103254
rect 569786 102698 570022 102934
rect 569786 67018 570022 67254
rect 569786 66698 570022 66934
rect 569786 31018 570022 31254
rect 569786 30698 570022 30934
rect 551786 -6102 552022 -5866
rect 551786 -6422 552022 -6186
rect 576986 704602 577222 704838
rect 576986 704282 577222 704518
rect 576986 686218 577222 686454
rect 576986 685898 577222 686134
rect 576986 650218 577222 650454
rect 576986 649898 577222 650134
rect 576986 614218 577222 614454
rect 576986 613898 577222 614134
rect 576986 578218 577222 578454
rect 576986 577898 577222 578134
rect 576986 542218 577222 542454
rect 576986 541898 577222 542134
rect 576986 506218 577222 506454
rect 576986 505898 577222 506134
rect 576986 470218 577222 470454
rect 576986 469898 577222 470134
rect 576986 434218 577222 434454
rect 576986 433898 577222 434134
rect 576986 398218 577222 398454
rect 576986 397898 577222 398134
rect 576986 362218 577222 362454
rect 576986 361898 577222 362134
rect 576986 326218 577222 326454
rect 576986 325898 577222 326134
rect 576986 290218 577222 290454
rect 576986 289898 577222 290134
rect 576986 254218 577222 254454
rect 576986 253898 577222 254134
rect 576986 218218 577222 218454
rect 576986 217898 577222 218134
rect 576986 182218 577222 182454
rect 576986 181898 577222 182134
rect 576986 146218 577222 146454
rect 576986 145898 577222 146134
rect 576986 110218 577222 110454
rect 576986 109898 577222 110134
rect 576986 74218 577222 74454
rect 576986 73898 577222 74134
rect 576986 38218 577222 38454
rect 576986 37898 577222 38134
rect 576986 2218 577222 2454
rect 576986 1898 577222 2134
rect 576986 -582 577222 -346
rect 576986 -902 577222 -666
rect 587342 706442 587578 706678
rect 587342 706122 587578 706358
rect 586422 705522 586658 705758
rect 586422 705202 586658 705438
rect 580586 689818 580822 690054
rect 580586 689498 580822 689734
rect 580586 653818 580822 654054
rect 580586 653498 580822 653734
rect 580586 617818 580822 618054
rect 580586 617498 580822 617734
rect 580586 581818 580822 582054
rect 580586 581498 580822 581734
rect 580586 545818 580822 546054
rect 580586 545498 580822 545734
rect 580586 509818 580822 510054
rect 580586 509498 580822 509734
rect 580586 473818 580822 474054
rect 580586 473498 580822 473734
rect 580586 437818 580822 438054
rect 580586 437498 580822 437734
rect 580586 401818 580822 402054
rect 580586 401498 580822 401734
rect 580586 365818 580822 366054
rect 580586 365498 580822 365734
rect 580586 329818 580822 330054
rect 580586 329498 580822 329734
rect 580586 293818 580822 294054
rect 580586 293498 580822 293734
rect 580586 257818 580822 258054
rect 580586 257498 580822 257734
rect 580586 221818 580822 222054
rect 580586 221498 580822 221734
rect 580586 185818 580822 186054
rect 580586 185498 580822 185734
rect 580586 149818 580822 150054
rect 580586 149498 580822 149734
rect 580586 113818 580822 114054
rect 580586 113498 580822 113734
rect 580586 77818 580822 78054
rect 580586 77498 580822 77734
rect 580586 41818 580822 42054
rect 580586 41498 580822 41734
rect 580586 5818 580822 6054
rect 580586 5498 580822 5734
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 686218 585738 686454
rect 585502 685898 585738 686134
rect 585502 650218 585738 650454
rect 585502 649898 585738 650134
rect 585502 614218 585738 614454
rect 585502 613898 585738 614134
rect 585502 578218 585738 578454
rect 585502 577898 585738 578134
rect 585502 542218 585738 542454
rect 585502 541898 585738 542134
rect 585502 506218 585738 506454
rect 585502 505898 585738 506134
rect 585502 470218 585738 470454
rect 585502 469898 585738 470134
rect 585502 434218 585738 434454
rect 585502 433898 585738 434134
rect 585502 398218 585738 398454
rect 585502 397898 585738 398134
rect 585502 362218 585738 362454
rect 585502 361898 585738 362134
rect 585502 326218 585738 326454
rect 585502 325898 585738 326134
rect 585502 290218 585738 290454
rect 585502 289898 585738 290134
rect 585502 254218 585738 254454
rect 585502 253898 585738 254134
rect 585502 218218 585738 218454
rect 585502 217898 585738 218134
rect 585502 182218 585738 182454
rect 585502 181898 585738 182134
rect 585502 146218 585738 146454
rect 585502 145898 585738 146134
rect 585502 110218 585738 110454
rect 585502 109898 585738 110134
rect 585502 74218 585738 74454
rect 585502 73898 585738 74134
rect 585502 38218 585738 38454
rect 585502 37898 585738 38134
rect 585502 2218 585738 2454
rect 585502 1898 585738 2134
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586422 668218 586658 668454
rect 586422 667898 586658 668134
rect 586422 632218 586658 632454
rect 586422 631898 586658 632134
rect 586422 596218 586658 596454
rect 586422 595898 586658 596134
rect 586422 560218 586658 560454
rect 586422 559898 586658 560134
rect 586422 524218 586658 524454
rect 586422 523898 586658 524134
rect 586422 488218 586658 488454
rect 586422 487898 586658 488134
rect 586422 452218 586658 452454
rect 586422 451898 586658 452134
rect 586422 416218 586658 416454
rect 586422 415898 586658 416134
rect 586422 380218 586658 380454
rect 586422 379898 586658 380134
rect 586422 344218 586658 344454
rect 586422 343898 586658 344134
rect 586422 308218 586658 308454
rect 586422 307898 586658 308134
rect 586422 272218 586658 272454
rect 586422 271898 586658 272134
rect 586422 236218 586658 236454
rect 586422 235898 586658 236134
rect 586422 200218 586658 200454
rect 586422 199898 586658 200134
rect 586422 164218 586658 164454
rect 586422 163898 586658 164134
rect 586422 128218 586658 128454
rect 586422 127898 586658 128134
rect 586422 92218 586658 92454
rect 586422 91898 586658 92134
rect 586422 56218 586658 56454
rect 586422 55898 586658 56134
rect 586422 20218 586658 20454
rect 586422 19898 586658 20134
rect 586422 -1502 586658 -1266
rect 586422 -1822 586658 -1586
rect 587342 689818 587578 690054
rect 587342 689498 587578 689734
rect 587342 653818 587578 654054
rect 587342 653498 587578 653734
rect 587342 617818 587578 618054
rect 587342 617498 587578 617734
rect 587342 581818 587578 582054
rect 587342 581498 587578 581734
rect 587342 545818 587578 546054
rect 587342 545498 587578 545734
rect 587342 509818 587578 510054
rect 587342 509498 587578 509734
rect 587342 473818 587578 474054
rect 587342 473498 587578 473734
rect 587342 437818 587578 438054
rect 587342 437498 587578 437734
rect 587342 401818 587578 402054
rect 587342 401498 587578 401734
rect 587342 365818 587578 366054
rect 587342 365498 587578 365734
rect 587342 329818 587578 330054
rect 587342 329498 587578 329734
rect 587342 293818 587578 294054
rect 587342 293498 587578 293734
rect 587342 257818 587578 258054
rect 587342 257498 587578 257734
rect 587342 221818 587578 222054
rect 587342 221498 587578 221734
rect 587342 185818 587578 186054
rect 587342 185498 587578 185734
rect 587342 149818 587578 150054
rect 587342 149498 587578 149734
rect 587342 113818 587578 114054
rect 587342 113498 587578 113734
rect 587342 77818 587578 78054
rect 587342 77498 587578 77734
rect 587342 41818 587578 42054
rect 587342 41498 587578 41734
rect 587342 5818 587578 6054
rect 587342 5498 587578 5734
rect 580586 -2422 580822 -2186
rect 580586 -2742 580822 -2506
rect 587342 -2422 587578 -2186
rect 587342 -2742 587578 -2506
rect 588262 671818 588498 672054
rect 588262 671498 588498 671734
rect 588262 635818 588498 636054
rect 588262 635498 588498 635734
rect 588262 599818 588498 600054
rect 588262 599498 588498 599734
rect 588262 563818 588498 564054
rect 588262 563498 588498 563734
rect 588262 527818 588498 528054
rect 588262 527498 588498 527734
rect 588262 491818 588498 492054
rect 588262 491498 588498 491734
rect 588262 455818 588498 456054
rect 588262 455498 588498 455734
rect 588262 419818 588498 420054
rect 588262 419498 588498 419734
rect 588262 383818 588498 384054
rect 588262 383498 588498 383734
rect 588262 347818 588498 348054
rect 588262 347498 588498 347734
rect 588262 311818 588498 312054
rect 588262 311498 588498 311734
rect 588262 275818 588498 276054
rect 588262 275498 588498 275734
rect 588262 239818 588498 240054
rect 588262 239498 588498 239734
rect 588262 203818 588498 204054
rect 588262 203498 588498 203734
rect 588262 167818 588498 168054
rect 588262 167498 588498 167734
rect 588262 131818 588498 132054
rect 588262 131498 588498 131734
rect 588262 95818 588498 96054
rect 588262 95498 588498 95734
rect 588262 59818 588498 60054
rect 588262 59498 588498 59734
rect 588262 23818 588498 24054
rect 588262 23498 588498 23734
rect 588262 -3342 588498 -3106
rect 588262 -3662 588498 -3426
rect 589182 693418 589418 693654
rect 589182 693098 589418 693334
rect 589182 657418 589418 657654
rect 589182 657098 589418 657334
rect 589182 621418 589418 621654
rect 589182 621098 589418 621334
rect 589182 585418 589418 585654
rect 589182 585098 589418 585334
rect 589182 549418 589418 549654
rect 589182 549098 589418 549334
rect 589182 513418 589418 513654
rect 589182 513098 589418 513334
rect 589182 477418 589418 477654
rect 589182 477098 589418 477334
rect 589182 441418 589418 441654
rect 589182 441098 589418 441334
rect 589182 405418 589418 405654
rect 589182 405098 589418 405334
rect 589182 369418 589418 369654
rect 589182 369098 589418 369334
rect 589182 333418 589418 333654
rect 589182 333098 589418 333334
rect 589182 297418 589418 297654
rect 589182 297098 589418 297334
rect 589182 261418 589418 261654
rect 589182 261098 589418 261334
rect 589182 225418 589418 225654
rect 589182 225098 589418 225334
rect 589182 189418 589418 189654
rect 589182 189098 589418 189334
rect 589182 153418 589418 153654
rect 589182 153098 589418 153334
rect 589182 117418 589418 117654
rect 589182 117098 589418 117334
rect 589182 81418 589418 81654
rect 589182 81098 589418 81334
rect 589182 45418 589418 45654
rect 589182 45098 589418 45334
rect 589182 9418 589418 9654
rect 589182 9098 589418 9334
rect 589182 -4262 589418 -4026
rect 589182 -4582 589418 -4346
rect 590102 675418 590338 675654
rect 590102 675098 590338 675334
rect 590102 639418 590338 639654
rect 590102 639098 590338 639334
rect 590102 603418 590338 603654
rect 590102 603098 590338 603334
rect 590102 567418 590338 567654
rect 590102 567098 590338 567334
rect 590102 531418 590338 531654
rect 590102 531098 590338 531334
rect 590102 495418 590338 495654
rect 590102 495098 590338 495334
rect 590102 459418 590338 459654
rect 590102 459098 590338 459334
rect 590102 423418 590338 423654
rect 590102 423098 590338 423334
rect 590102 387418 590338 387654
rect 590102 387098 590338 387334
rect 590102 351418 590338 351654
rect 590102 351098 590338 351334
rect 590102 315418 590338 315654
rect 590102 315098 590338 315334
rect 590102 279418 590338 279654
rect 590102 279098 590338 279334
rect 590102 243418 590338 243654
rect 590102 243098 590338 243334
rect 590102 207418 590338 207654
rect 590102 207098 590338 207334
rect 590102 171418 590338 171654
rect 590102 171098 590338 171334
rect 590102 135418 590338 135654
rect 590102 135098 590338 135334
rect 590102 99418 590338 99654
rect 590102 99098 590338 99334
rect 590102 63418 590338 63654
rect 590102 63098 590338 63334
rect 590102 27418 590338 27654
rect 590102 27098 590338 27334
rect 590102 -5182 590338 -4946
rect 590102 -5502 590338 -5266
rect 591022 697018 591258 697254
rect 591022 696698 591258 696934
rect 591022 661018 591258 661254
rect 591022 660698 591258 660934
rect 591022 625018 591258 625254
rect 591022 624698 591258 624934
rect 591022 589018 591258 589254
rect 591022 588698 591258 588934
rect 591022 553018 591258 553254
rect 591022 552698 591258 552934
rect 591022 517018 591258 517254
rect 591022 516698 591258 516934
rect 591022 481018 591258 481254
rect 591022 480698 591258 480934
rect 591022 445018 591258 445254
rect 591022 444698 591258 444934
rect 591022 409018 591258 409254
rect 591022 408698 591258 408934
rect 591022 373018 591258 373254
rect 591022 372698 591258 372934
rect 591022 337018 591258 337254
rect 591022 336698 591258 336934
rect 591022 301018 591258 301254
rect 591022 300698 591258 300934
rect 591022 265018 591258 265254
rect 591022 264698 591258 264934
rect 591022 229018 591258 229254
rect 591022 228698 591258 228934
rect 591022 193018 591258 193254
rect 591022 192698 591258 192934
rect 591022 157018 591258 157254
rect 591022 156698 591258 156934
rect 591022 121018 591258 121254
rect 591022 120698 591258 120934
rect 591022 85018 591258 85254
rect 591022 84698 591258 84934
rect 591022 49018 591258 49254
rect 591022 48698 591258 48934
rect 591022 13018 591258 13254
rect 591022 12698 591258 12934
rect 591022 -6102 591258 -5866
rect 591022 -6422 591258 -6186
rect 591942 679018 592178 679254
rect 591942 678698 592178 678934
rect 591942 643018 592178 643254
rect 591942 642698 592178 642934
rect 591942 607018 592178 607254
rect 591942 606698 592178 606934
rect 591942 571018 592178 571254
rect 591942 570698 592178 570934
rect 591942 535018 592178 535254
rect 591942 534698 592178 534934
rect 591942 499018 592178 499254
rect 591942 498698 592178 498934
rect 591942 463018 592178 463254
rect 591942 462698 592178 462934
rect 591942 427018 592178 427254
rect 591942 426698 592178 426934
rect 591942 391018 592178 391254
rect 591942 390698 592178 390934
rect 591942 355018 592178 355254
rect 591942 354698 592178 354934
rect 591942 319018 592178 319254
rect 591942 318698 592178 318934
rect 591942 283018 592178 283254
rect 591942 282698 592178 282934
rect 591942 247018 592178 247254
rect 591942 246698 592178 246934
rect 591942 211018 592178 211254
rect 591942 210698 592178 210934
rect 591942 175018 592178 175254
rect 591942 174698 592178 174934
rect 591942 139018 592178 139254
rect 591942 138698 592178 138934
rect 591942 103018 592178 103254
rect 591942 102698 592178 102934
rect 591942 67018 592178 67254
rect 591942 66698 592178 66934
rect 591942 31018 592178 31254
rect 591942 30698 592178 30934
rect 569786 -7022 570022 -6786
rect 569786 -7342 570022 -7106
rect 591942 -7022 592178 -6786
rect 591942 -7342 592178 -7106
<< metal5 >>
rect -8436 711300 -7836 711302
rect 29604 711300 30204 711302
rect 65604 711300 66204 711302
rect 101604 711300 102204 711302
rect 137604 711300 138204 711302
rect 173604 711300 174204 711302
rect 209604 711300 210204 711302
rect 245604 711300 246204 711302
rect 281604 711300 282204 711302
rect 317604 711300 318204 711302
rect 353604 711300 354204 711302
rect 389604 711300 390204 711302
rect 425604 711300 426204 711302
rect 461604 711300 462204 711302
rect 497604 711300 498204 711302
rect 533604 711300 534204 711302
rect 569604 711300 570204 711302
rect 591760 711300 592360 711302
rect -8436 711278 592360 711300
rect -8436 711042 -8254 711278
rect -8018 711042 29786 711278
rect 30022 711042 65786 711278
rect 66022 711042 101786 711278
rect 102022 711042 137786 711278
rect 138022 711042 173786 711278
rect 174022 711042 209786 711278
rect 210022 711042 245786 711278
rect 246022 711042 281786 711278
rect 282022 711042 317786 711278
rect 318022 711042 353786 711278
rect 354022 711042 389786 711278
rect 390022 711042 425786 711278
rect 426022 711042 461786 711278
rect 462022 711042 497786 711278
rect 498022 711042 533786 711278
rect 534022 711042 569786 711278
rect 570022 711042 591942 711278
rect 592178 711042 592360 711278
rect -8436 710958 592360 711042
rect -8436 710722 -8254 710958
rect -8018 710722 29786 710958
rect 30022 710722 65786 710958
rect 66022 710722 101786 710958
rect 102022 710722 137786 710958
rect 138022 710722 173786 710958
rect 174022 710722 209786 710958
rect 210022 710722 245786 710958
rect 246022 710722 281786 710958
rect 282022 710722 317786 710958
rect 318022 710722 353786 710958
rect 354022 710722 389786 710958
rect 390022 710722 425786 710958
rect 426022 710722 461786 710958
rect 462022 710722 497786 710958
rect 498022 710722 533786 710958
rect 534022 710722 569786 710958
rect 570022 710722 591942 710958
rect 592178 710722 592360 710958
rect -8436 710700 592360 710722
rect -8436 710698 -7836 710700
rect 29604 710698 30204 710700
rect 65604 710698 66204 710700
rect 101604 710698 102204 710700
rect 137604 710698 138204 710700
rect 173604 710698 174204 710700
rect 209604 710698 210204 710700
rect 245604 710698 246204 710700
rect 281604 710698 282204 710700
rect 317604 710698 318204 710700
rect 353604 710698 354204 710700
rect 389604 710698 390204 710700
rect 425604 710698 426204 710700
rect 461604 710698 462204 710700
rect 497604 710698 498204 710700
rect 533604 710698 534204 710700
rect 569604 710698 570204 710700
rect 591760 710698 592360 710700
rect -7516 710380 -6916 710382
rect 11604 710380 12204 710382
rect 47604 710380 48204 710382
rect 83604 710380 84204 710382
rect 119604 710380 120204 710382
rect 155604 710380 156204 710382
rect 191604 710380 192204 710382
rect 227604 710380 228204 710382
rect 263604 710380 264204 710382
rect 299604 710380 300204 710382
rect 335604 710380 336204 710382
rect 371604 710380 372204 710382
rect 407604 710380 408204 710382
rect 443604 710380 444204 710382
rect 479604 710380 480204 710382
rect 515604 710380 516204 710382
rect 551604 710380 552204 710382
rect 590840 710380 591440 710382
rect -7516 710358 591440 710380
rect -7516 710122 -7334 710358
rect -7098 710122 11786 710358
rect 12022 710122 47786 710358
rect 48022 710122 83786 710358
rect 84022 710122 119786 710358
rect 120022 710122 155786 710358
rect 156022 710122 191786 710358
rect 192022 710122 227786 710358
rect 228022 710122 263786 710358
rect 264022 710122 299786 710358
rect 300022 710122 335786 710358
rect 336022 710122 371786 710358
rect 372022 710122 407786 710358
rect 408022 710122 443786 710358
rect 444022 710122 479786 710358
rect 480022 710122 515786 710358
rect 516022 710122 551786 710358
rect 552022 710122 591022 710358
rect 591258 710122 591440 710358
rect -7516 710038 591440 710122
rect -7516 709802 -7334 710038
rect -7098 709802 11786 710038
rect 12022 709802 47786 710038
rect 48022 709802 83786 710038
rect 84022 709802 119786 710038
rect 120022 709802 155786 710038
rect 156022 709802 191786 710038
rect 192022 709802 227786 710038
rect 228022 709802 263786 710038
rect 264022 709802 299786 710038
rect 300022 709802 335786 710038
rect 336022 709802 371786 710038
rect 372022 709802 407786 710038
rect 408022 709802 443786 710038
rect 444022 709802 479786 710038
rect 480022 709802 515786 710038
rect 516022 709802 551786 710038
rect 552022 709802 591022 710038
rect 591258 709802 591440 710038
rect -7516 709780 591440 709802
rect -7516 709778 -6916 709780
rect 11604 709778 12204 709780
rect 47604 709778 48204 709780
rect 83604 709778 84204 709780
rect 119604 709778 120204 709780
rect 155604 709778 156204 709780
rect 191604 709778 192204 709780
rect 227604 709778 228204 709780
rect 263604 709778 264204 709780
rect 299604 709778 300204 709780
rect 335604 709778 336204 709780
rect 371604 709778 372204 709780
rect 407604 709778 408204 709780
rect 443604 709778 444204 709780
rect 479604 709778 480204 709780
rect 515604 709778 516204 709780
rect 551604 709778 552204 709780
rect 590840 709778 591440 709780
rect -6596 709460 -5996 709462
rect 26004 709460 26604 709462
rect 62004 709460 62604 709462
rect 98004 709460 98604 709462
rect 134004 709460 134604 709462
rect 170004 709460 170604 709462
rect 206004 709460 206604 709462
rect 242004 709460 242604 709462
rect 278004 709460 278604 709462
rect 314004 709460 314604 709462
rect 350004 709460 350604 709462
rect 386004 709460 386604 709462
rect 422004 709460 422604 709462
rect 458004 709460 458604 709462
rect 494004 709460 494604 709462
rect 530004 709460 530604 709462
rect 566004 709460 566604 709462
rect 589920 709460 590520 709462
rect -6596 709438 590520 709460
rect -6596 709202 -6414 709438
rect -6178 709202 26186 709438
rect 26422 709202 62186 709438
rect 62422 709202 98186 709438
rect 98422 709202 134186 709438
rect 134422 709202 170186 709438
rect 170422 709202 206186 709438
rect 206422 709202 242186 709438
rect 242422 709202 278186 709438
rect 278422 709202 314186 709438
rect 314422 709202 350186 709438
rect 350422 709202 386186 709438
rect 386422 709202 422186 709438
rect 422422 709202 458186 709438
rect 458422 709202 494186 709438
rect 494422 709202 530186 709438
rect 530422 709202 566186 709438
rect 566422 709202 590102 709438
rect 590338 709202 590520 709438
rect -6596 709118 590520 709202
rect -6596 708882 -6414 709118
rect -6178 708882 26186 709118
rect 26422 708882 62186 709118
rect 62422 708882 98186 709118
rect 98422 708882 134186 709118
rect 134422 708882 170186 709118
rect 170422 708882 206186 709118
rect 206422 708882 242186 709118
rect 242422 708882 278186 709118
rect 278422 708882 314186 709118
rect 314422 708882 350186 709118
rect 350422 708882 386186 709118
rect 386422 708882 422186 709118
rect 422422 708882 458186 709118
rect 458422 708882 494186 709118
rect 494422 708882 530186 709118
rect 530422 708882 566186 709118
rect 566422 708882 590102 709118
rect 590338 708882 590520 709118
rect -6596 708860 590520 708882
rect -6596 708858 -5996 708860
rect 26004 708858 26604 708860
rect 62004 708858 62604 708860
rect 98004 708858 98604 708860
rect 134004 708858 134604 708860
rect 170004 708858 170604 708860
rect 206004 708858 206604 708860
rect 242004 708858 242604 708860
rect 278004 708858 278604 708860
rect 314004 708858 314604 708860
rect 350004 708858 350604 708860
rect 386004 708858 386604 708860
rect 422004 708858 422604 708860
rect 458004 708858 458604 708860
rect 494004 708858 494604 708860
rect 530004 708858 530604 708860
rect 566004 708858 566604 708860
rect 589920 708858 590520 708860
rect -5676 708540 -5076 708542
rect 8004 708540 8604 708542
rect 44004 708540 44604 708542
rect 80004 708540 80604 708542
rect 116004 708540 116604 708542
rect 152004 708540 152604 708542
rect 188004 708540 188604 708542
rect 224004 708540 224604 708542
rect 260004 708540 260604 708542
rect 296004 708540 296604 708542
rect 332004 708540 332604 708542
rect 368004 708540 368604 708542
rect 404004 708540 404604 708542
rect 440004 708540 440604 708542
rect 476004 708540 476604 708542
rect 512004 708540 512604 708542
rect 548004 708540 548604 708542
rect 589000 708540 589600 708542
rect -5676 708518 589600 708540
rect -5676 708282 -5494 708518
rect -5258 708282 8186 708518
rect 8422 708282 44186 708518
rect 44422 708282 80186 708518
rect 80422 708282 116186 708518
rect 116422 708282 152186 708518
rect 152422 708282 188186 708518
rect 188422 708282 224186 708518
rect 224422 708282 260186 708518
rect 260422 708282 296186 708518
rect 296422 708282 332186 708518
rect 332422 708282 368186 708518
rect 368422 708282 404186 708518
rect 404422 708282 440186 708518
rect 440422 708282 476186 708518
rect 476422 708282 512186 708518
rect 512422 708282 548186 708518
rect 548422 708282 589182 708518
rect 589418 708282 589600 708518
rect -5676 708198 589600 708282
rect -5676 707962 -5494 708198
rect -5258 707962 8186 708198
rect 8422 707962 44186 708198
rect 44422 707962 80186 708198
rect 80422 707962 116186 708198
rect 116422 707962 152186 708198
rect 152422 707962 188186 708198
rect 188422 707962 224186 708198
rect 224422 707962 260186 708198
rect 260422 707962 296186 708198
rect 296422 707962 332186 708198
rect 332422 707962 368186 708198
rect 368422 707962 404186 708198
rect 404422 707962 440186 708198
rect 440422 707962 476186 708198
rect 476422 707962 512186 708198
rect 512422 707962 548186 708198
rect 548422 707962 589182 708198
rect 589418 707962 589600 708198
rect -5676 707940 589600 707962
rect -5676 707938 -5076 707940
rect 8004 707938 8604 707940
rect 44004 707938 44604 707940
rect 80004 707938 80604 707940
rect 116004 707938 116604 707940
rect 152004 707938 152604 707940
rect 188004 707938 188604 707940
rect 224004 707938 224604 707940
rect 260004 707938 260604 707940
rect 296004 707938 296604 707940
rect 332004 707938 332604 707940
rect 368004 707938 368604 707940
rect 404004 707938 404604 707940
rect 440004 707938 440604 707940
rect 476004 707938 476604 707940
rect 512004 707938 512604 707940
rect 548004 707938 548604 707940
rect 589000 707938 589600 707940
rect -4756 707620 -4156 707622
rect 22404 707620 23004 707622
rect 58404 707620 59004 707622
rect 94404 707620 95004 707622
rect 130404 707620 131004 707622
rect 166404 707620 167004 707622
rect 202404 707620 203004 707622
rect 238404 707620 239004 707622
rect 274404 707620 275004 707622
rect 310404 707620 311004 707622
rect 346404 707620 347004 707622
rect 382404 707620 383004 707622
rect 418404 707620 419004 707622
rect 454404 707620 455004 707622
rect 490404 707620 491004 707622
rect 526404 707620 527004 707622
rect 562404 707620 563004 707622
rect 588080 707620 588680 707622
rect -4756 707598 588680 707620
rect -4756 707362 -4574 707598
rect -4338 707362 22586 707598
rect 22822 707362 58586 707598
rect 58822 707362 94586 707598
rect 94822 707362 130586 707598
rect 130822 707362 166586 707598
rect 166822 707362 202586 707598
rect 202822 707362 238586 707598
rect 238822 707362 274586 707598
rect 274822 707362 310586 707598
rect 310822 707362 346586 707598
rect 346822 707362 382586 707598
rect 382822 707362 418586 707598
rect 418822 707362 454586 707598
rect 454822 707362 490586 707598
rect 490822 707362 526586 707598
rect 526822 707362 562586 707598
rect 562822 707362 588262 707598
rect 588498 707362 588680 707598
rect -4756 707278 588680 707362
rect -4756 707042 -4574 707278
rect -4338 707042 22586 707278
rect 22822 707042 58586 707278
rect 58822 707042 94586 707278
rect 94822 707042 130586 707278
rect 130822 707042 166586 707278
rect 166822 707042 202586 707278
rect 202822 707042 238586 707278
rect 238822 707042 274586 707278
rect 274822 707042 310586 707278
rect 310822 707042 346586 707278
rect 346822 707042 382586 707278
rect 382822 707042 418586 707278
rect 418822 707042 454586 707278
rect 454822 707042 490586 707278
rect 490822 707042 526586 707278
rect 526822 707042 562586 707278
rect 562822 707042 588262 707278
rect 588498 707042 588680 707278
rect -4756 707020 588680 707042
rect -4756 707018 -4156 707020
rect 22404 707018 23004 707020
rect 58404 707018 59004 707020
rect 94404 707018 95004 707020
rect 130404 707018 131004 707020
rect 166404 707018 167004 707020
rect 202404 707018 203004 707020
rect 238404 707018 239004 707020
rect 274404 707018 275004 707020
rect 310404 707018 311004 707020
rect 346404 707018 347004 707020
rect 382404 707018 383004 707020
rect 418404 707018 419004 707020
rect 454404 707018 455004 707020
rect 490404 707018 491004 707020
rect 526404 707018 527004 707020
rect 562404 707018 563004 707020
rect 588080 707018 588680 707020
rect -3836 706700 -3236 706702
rect 4404 706700 5004 706702
rect 40404 706700 41004 706702
rect 76404 706700 77004 706702
rect 112404 706700 113004 706702
rect 148404 706700 149004 706702
rect 184404 706700 185004 706702
rect 220404 706700 221004 706702
rect 256404 706700 257004 706702
rect 292404 706700 293004 706702
rect 328404 706700 329004 706702
rect 364404 706700 365004 706702
rect 400404 706700 401004 706702
rect 436404 706700 437004 706702
rect 472404 706700 473004 706702
rect 508404 706700 509004 706702
rect 544404 706700 545004 706702
rect 580404 706700 581004 706702
rect 587160 706700 587760 706702
rect -3836 706678 587760 706700
rect -3836 706442 -3654 706678
rect -3418 706442 4586 706678
rect 4822 706442 40586 706678
rect 40822 706442 76586 706678
rect 76822 706442 112586 706678
rect 112822 706442 148586 706678
rect 148822 706442 184586 706678
rect 184822 706442 220586 706678
rect 220822 706442 256586 706678
rect 256822 706442 292586 706678
rect 292822 706442 328586 706678
rect 328822 706442 364586 706678
rect 364822 706442 400586 706678
rect 400822 706442 436586 706678
rect 436822 706442 472586 706678
rect 472822 706442 508586 706678
rect 508822 706442 544586 706678
rect 544822 706442 580586 706678
rect 580822 706442 587342 706678
rect 587578 706442 587760 706678
rect -3836 706358 587760 706442
rect -3836 706122 -3654 706358
rect -3418 706122 4586 706358
rect 4822 706122 40586 706358
rect 40822 706122 76586 706358
rect 76822 706122 112586 706358
rect 112822 706122 148586 706358
rect 148822 706122 184586 706358
rect 184822 706122 220586 706358
rect 220822 706122 256586 706358
rect 256822 706122 292586 706358
rect 292822 706122 328586 706358
rect 328822 706122 364586 706358
rect 364822 706122 400586 706358
rect 400822 706122 436586 706358
rect 436822 706122 472586 706358
rect 472822 706122 508586 706358
rect 508822 706122 544586 706358
rect 544822 706122 580586 706358
rect 580822 706122 587342 706358
rect 587578 706122 587760 706358
rect -3836 706100 587760 706122
rect -3836 706098 -3236 706100
rect 4404 706098 5004 706100
rect 40404 706098 41004 706100
rect 76404 706098 77004 706100
rect 112404 706098 113004 706100
rect 148404 706098 149004 706100
rect 184404 706098 185004 706100
rect 220404 706098 221004 706100
rect 256404 706098 257004 706100
rect 292404 706098 293004 706100
rect 328404 706098 329004 706100
rect 364404 706098 365004 706100
rect 400404 706098 401004 706100
rect 436404 706098 437004 706100
rect 472404 706098 473004 706100
rect 508404 706098 509004 706100
rect 544404 706098 545004 706100
rect 580404 706098 581004 706100
rect 587160 706098 587760 706100
rect -2916 705780 -2316 705782
rect 18804 705780 19404 705782
rect 54804 705780 55404 705782
rect 90804 705780 91404 705782
rect 126804 705780 127404 705782
rect 162804 705780 163404 705782
rect 198804 705780 199404 705782
rect 234804 705780 235404 705782
rect 270804 705780 271404 705782
rect 306804 705780 307404 705782
rect 342804 705780 343404 705782
rect 378804 705780 379404 705782
rect 414804 705780 415404 705782
rect 450804 705780 451404 705782
rect 486804 705780 487404 705782
rect 522804 705780 523404 705782
rect 558804 705780 559404 705782
rect 586240 705780 586840 705782
rect -2916 705758 586840 705780
rect -2916 705522 -2734 705758
rect -2498 705522 18986 705758
rect 19222 705522 54986 705758
rect 55222 705522 90986 705758
rect 91222 705522 126986 705758
rect 127222 705522 162986 705758
rect 163222 705522 198986 705758
rect 199222 705522 234986 705758
rect 235222 705522 270986 705758
rect 271222 705522 306986 705758
rect 307222 705522 342986 705758
rect 343222 705522 378986 705758
rect 379222 705522 414986 705758
rect 415222 705522 450986 705758
rect 451222 705522 486986 705758
rect 487222 705522 522986 705758
rect 523222 705522 558986 705758
rect 559222 705522 586422 705758
rect 586658 705522 586840 705758
rect -2916 705438 586840 705522
rect -2916 705202 -2734 705438
rect -2498 705202 18986 705438
rect 19222 705202 54986 705438
rect 55222 705202 90986 705438
rect 91222 705202 126986 705438
rect 127222 705202 162986 705438
rect 163222 705202 198986 705438
rect 199222 705202 234986 705438
rect 235222 705202 270986 705438
rect 271222 705202 306986 705438
rect 307222 705202 342986 705438
rect 343222 705202 378986 705438
rect 379222 705202 414986 705438
rect 415222 705202 450986 705438
rect 451222 705202 486986 705438
rect 487222 705202 522986 705438
rect 523222 705202 558986 705438
rect 559222 705202 586422 705438
rect 586658 705202 586840 705438
rect -2916 705180 586840 705202
rect -2916 705178 -2316 705180
rect 18804 705178 19404 705180
rect 54804 705178 55404 705180
rect 90804 705178 91404 705180
rect 126804 705178 127404 705180
rect 162804 705178 163404 705180
rect 198804 705178 199404 705180
rect 234804 705178 235404 705180
rect 270804 705178 271404 705180
rect 306804 705178 307404 705180
rect 342804 705178 343404 705180
rect 378804 705178 379404 705180
rect 414804 705178 415404 705180
rect 450804 705178 451404 705180
rect 486804 705178 487404 705180
rect 522804 705178 523404 705180
rect 558804 705178 559404 705180
rect 586240 705178 586840 705180
rect -1996 704860 -1396 704862
rect 804 704860 1404 704862
rect 36804 704860 37404 704862
rect 72804 704860 73404 704862
rect 108804 704860 109404 704862
rect 144804 704860 145404 704862
rect 180804 704860 181404 704862
rect 216804 704860 217404 704862
rect 252804 704860 253404 704862
rect 288804 704860 289404 704862
rect 324804 704860 325404 704862
rect 360804 704860 361404 704862
rect 396804 704860 397404 704862
rect 432804 704860 433404 704862
rect 468804 704860 469404 704862
rect 504804 704860 505404 704862
rect 540804 704860 541404 704862
rect 576804 704860 577404 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 986 704838
rect 1222 704602 36986 704838
rect 37222 704602 72986 704838
rect 73222 704602 108986 704838
rect 109222 704602 144986 704838
rect 145222 704602 180986 704838
rect 181222 704602 216986 704838
rect 217222 704602 252986 704838
rect 253222 704602 288986 704838
rect 289222 704602 324986 704838
rect 325222 704602 360986 704838
rect 361222 704602 396986 704838
rect 397222 704602 432986 704838
rect 433222 704602 468986 704838
rect 469222 704602 504986 704838
rect 505222 704602 540986 704838
rect 541222 704602 576986 704838
rect 577222 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 986 704518
rect 1222 704282 36986 704518
rect 37222 704282 72986 704518
rect 73222 704282 108986 704518
rect 109222 704282 144986 704518
rect 145222 704282 180986 704518
rect 181222 704282 216986 704518
rect 217222 704282 252986 704518
rect 253222 704282 288986 704518
rect 289222 704282 324986 704518
rect 325222 704282 360986 704518
rect 361222 704282 396986 704518
rect 397222 704282 432986 704518
rect 433222 704282 468986 704518
rect 469222 704282 504986 704518
rect 505222 704282 540986 704518
rect 541222 704282 576986 704518
rect 577222 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 804 704258 1404 704260
rect 36804 704258 37404 704260
rect 72804 704258 73404 704260
rect 108804 704258 109404 704260
rect 144804 704258 145404 704260
rect 180804 704258 181404 704260
rect 216804 704258 217404 704260
rect 252804 704258 253404 704260
rect 288804 704258 289404 704260
rect 324804 704258 325404 704260
rect 360804 704258 361404 704260
rect 396804 704258 397404 704260
rect 432804 704258 433404 704260
rect 468804 704258 469404 704260
rect 504804 704258 505404 704260
rect 540804 704258 541404 704260
rect 576804 704258 577404 704260
rect 585320 704258 585920 704260
rect -7516 697276 -6916 697278
rect 11604 697276 12204 697278
rect 47604 697276 48204 697278
rect 83604 697276 84204 697278
rect 119604 697276 120204 697278
rect 155604 697276 156204 697278
rect 191604 697276 192204 697278
rect 227604 697276 228204 697278
rect 263604 697276 264204 697278
rect 299604 697276 300204 697278
rect 335604 697276 336204 697278
rect 371604 697276 372204 697278
rect 407604 697276 408204 697278
rect 443604 697276 444204 697278
rect 479604 697276 480204 697278
rect 515604 697276 516204 697278
rect 551604 697276 552204 697278
rect 590840 697276 591440 697278
rect -8436 697254 592360 697276
rect -8436 697018 -7334 697254
rect -7098 697018 11786 697254
rect 12022 697018 47786 697254
rect 48022 697018 83786 697254
rect 84022 697018 119786 697254
rect 120022 697018 155786 697254
rect 156022 697018 191786 697254
rect 192022 697018 227786 697254
rect 228022 697018 263786 697254
rect 264022 697018 299786 697254
rect 300022 697018 335786 697254
rect 336022 697018 371786 697254
rect 372022 697018 407786 697254
rect 408022 697018 443786 697254
rect 444022 697018 479786 697254
rect 480022 697018 515786 697254
rect 516022 697018 551786 697254
rect 552022 697018 591022 697254
rect 591258 697018 592360 697254
rect -8436 696934 592360 697018
rect -8436 696698 -7334 696934
rect -7098 696698 11786 696934
rect 12022 696698 47786 696934
rect 48022 696698 83786 696934
rect 84022 696698 119786 696934
rect 120022 696698 155786 696934
rect 156022 696698 191786 696934
rect 192022 696698 227786 696934
rect 228022 696698 263786 696934
rect 264022 696698 299786 696934
rect 300022 696698 335786 696934
rect 336022 696698 371786 696934
rect 372022 696698 407786 696934
rect 408022 696698 443786 696934
rect 444022 696698 479786 696934
rect 480022 696698 515786 696934
rect 516022 696698 551786 696934
rect 552022 696698 591022 696934
rect 591258 696698 592360 696934
rect -8436 696676 592360 696698
rect -7516 696674 -6916 696676
rect 11604 696674 12204 696676
rect 47604 696674 48204 696676
rect 83604 696674 84204 696676
rect 119604 696674 120204 696676
rect 155604 696674 156204 696676
rect 191604 696674 192204 696676
rect 227604 696674 228204 696676
rect 263604 696674 264204 696676
rect 299604 696674 300204 696676
rect 335604 696674 336204 696676
rect 371604 696674 372204 696676
rect 407604 696674 408204 696676
rect 443604 696674 444204 696676
rect 479604 696674 480204 696676
rect 515604 696674 516204 696676
rect 551604 696674 552204 696676
rect 590840 696674 591440 696676
rect -5676 693676 -5076 693678
rect 8004 693676 8604 693678
rect 44004 693676 44604 693678
rect 80004 693676 80604 693678
rect 116004 693676 116604 693678
rect 152004 693676 152604 693678
rect 188004 693676 188604 693678
rect 224004 693676 224604 693678
rect 260004 693676 260604 693678
rect 296004 693676 296604 693678
rect 332004 693676 332604 693678
rect 368004 693676 368604 693678
rect 404004 693676 404604 693678
rect 440004 693676 440604 693678
rect 476004 693676 476604 693678
rect 512004 693676 512604 693678
rect 548004 693676 548604 693678
rect 589000 693676 589600 693678
rect -6596 693654 590520 693676
rect -6596 693418 -5494 693654
rect -5258 693418 8186 693654
rect 8422 693418 44186 693654
rect 44422 693418 80186 693654
rect 80422 693418 116186 693654
rect 116422 693418 152186 693654
rect 152422 693418 188186 693654
rect 188422 693418 224186 693654
rect 224422 693418 260186 693654
rect 260422 693418 296186 693654
rect 296422 693418 332186 693654
rect 332422 693418 368186 693654
rect 368422 693418 404186 693654
rect 404422 693418 440186 693654
rect 440422 693418 476186 693654
rect 476422 693418 512186 693654
rect 512422 693418 548186 693654
rect 548422 693418 589182 693654
rect 589418 693418 590520 693654
rect -6596 693334 590520 693418
rect -6596 693098 -5494 693334
rect -5258 693098 8186 693334
rect 8422 693098 44186 693334
rect 44422 693098 80186 693334
rect 80422 693098 116186 693334
rect 116422 693098 152186 693334
rect 152422 693098 188186 693334
rect 188422 693098 224186 693334
rect 224422 693098 260186 693334
rect 260422 693098 296186 693334
rect 296422 693098 332186 693334
rect 332422 693098 368186 693334
rect 368422 693098 404186 693334
rect 404422 693098 440186 693334
rect 440422 693098 476186 693334
rect 476422 693098 512186 693334
rect 512422 693098 548186 693334
rect 548422 693098 589182 693334
rect 589418 693098 590520 693334
rect -6596 693076 590520 693098
rect -5676 693074 -5076 693076
rect 8004 693074 8604 693076
rect 44004 693074 44604 693076
rect 80004 693074 80604 693076
rect 116004 693074 116604 693076
rect 152004 693074 152604 693076
rect 188004 693074 188604 693076
rect 224004 693074 224604 693076
rect 260004 693074 260604 693076
rect 296004 693074 296604 693076
rect 332004 693074 332604 693076
rect 368004 693074 368604 693076
rect 404004 693074 404604 693076
rect 440004 693074 440604 693076
rect 476004 693074 476604 693076
rect 512004 693074 512604 693076
rect 548004 693074 548604 693076
rect 589000 693074 589600 693076
rect -3836 690076 -3236 690078
rect 4404 690076 5004 690078
rect 40404 690076 41004 690078
rect 76404 690076 77004 690078
rect 112404 690076 113004 690078
rect 148404 690076 149004 690078
rect 184404 690076 185004 690078
rect 220404 690076 221004 690078
rect 256404 690076 257004 690078
rect 292404 690076 293004 690078
rect 328404 690076 329004 690078
rect 364404 690076 365004 690078
rect 400404 690076 401004 690078
rect 436404 690076 437004 690078
rect 472404 690076 473004 690078
rect 508404 690076 509004 690078
rect 544404 690076 545004 690078
rect 580404 690076 581004 690078
rect 587160 690076 587760 690078
rect -4756 690054 588680 690076
rect -4756 689818 -3654 690054
rect -3418 689818 4586 690054
rect 4822 689818 40586 690054
rect 40822 689818 76586 690054
rect 76822 689818 112586 690054
rect 112822 689818 148586 690054
rect 148822 689818 184586 690054
rect 184822 689818 220586 690054
rect 220822 689818 256586 690054
rect 256822 689818 292586 690054
rect 292822 689818 328586 690054
rect 328822 689818 364586 690054
rect 364822 689818 400586 690054
rect 400822 689818 436586 690054
rect 436822 689818 472586 690054
rect 472822 689818 508586 690054
rect 508822 689818 544586 690054
rect 544822 689818 580586 690054
rect 580822 689818 587342 690054
rect 587578 689818 588680 690054
rect -4756 689734 588680 689818
rect -4756 689498 -3654 689734
rect -3418 689498 4586 689734
rect 4822 689498 40586 689734
rect 40822 689498 76586 689734
rect 76822 689498 112586 689734
rect 112822 689498 148586 689734
rect 148822 689498 184586 689734
rect 184822 689498 220586 689734
rect 220822 689498 256586 689734
rect 256822 689498 292586 689734
rect 292822 689498 328586 689734
rect 328822 689498 364586 689734
rect 364822 689498 400586 689734
rect 400822 689498 436586 689734
rect 436822 689498 472586 689734
rect 472822 689498 508586 689734
rect 508822 689498 544586 689734
rect 544822 689498 580586 689734
rect 580822 689498 587342 689734
rect 587578 689498 588680 689734
rect -4756 689476 588680 689498
rect -3836 689474 -3236 689476
rect 4404 689474 5004 689476
rect 40404 689474 41004 689476
rect 76404 689474 77004 689476
rect 112404 689474 113004 689476
rect 148404 689474 149004 689476
rect 184404 689474 185004 689476
rect 220404 689474 221004 689476
rect 256404 689474 257004 689476
rect 292404 689474 293004 689476
rect 328404 689474 329004 689476
rect 364404 689474 365004 689476
rect 400404 689474 401004 689476
rect 436404 689474 437004 689476
rect 472404 689474 473004 689476
rect 508404 689474 509004 689476
rect 544404 689474 545004 689476
rect 580404 689474 581004 689476
rect 587160 689474 587760 689476
rect -1996 686476 -1396 686478
rect 804 686476 1404 686478
rect 36804 686476 37404 686478
rect 72804 686476 73404 686478
rect 108804 686476 109404 686478
rect 144804 686476 145404 686478
rect 180804 686476 181404 686478
rect 216804 686476 217404 686478
rect 252804 686476 253404 686478
rect 288804 686476 289404 686478
rect 324804 686476 325404 686478
rect 360804 686476 361404 686478
rect 396804 686476 397404 686478
rect 432804 686476 433404 686478
rect 468804 686476 469404 686478
rect 504804 686476 505404 686478
rect 540804 686476 541404 686478
rect 576804 686476 577404 686478
rect 585320 686476 585920 686478
rect -2916 686454 586840 686476
rect -2916 686218 -1814 686454
rect -1578 686218 986 686454
rect 1222 686218 36986 686454
rect 37222 686218 72986 686454
rect 73222 686218 108986 686454
rect 109222 686218 144986 686454
rect 145222 686218 180986 686454
rect 181222 686218 216986 686454
rect 217222 686218 252986 686454
rect 253222 686218 288986 686454
rect 289222 686218 324986 686454
rect 325222 686218 360986 686454
rect 361222 686218 396986 686454
rect 397222 686218 432986 686454
rect 433222 686218 468986 686454
rect 469222 686218 504986 686454
rect 505222 686218 540986 686454
rect 541222 686218 576986 686454
rect 577222 686218 585502 686454
rect 585738 686218 586840 686454
rect -2916 686134 586840 686218
rect -2916 685898 -1814 686134
rect -1578 685898 986 686134
rect 1222 685898 36986 686134
rect 37222 685898 72986 686134
rect 73222 685898 108986 686134
rect 109222 685898 144986 686134
rect 145222 685898 180986 686134
rect 181222 685898 216986 686134
rect 217222 685898 252986 686134
rect 253222 685898 288986 686134
rect 289222 685898 324986 686134
rect 325222 685898 360986 686134
rect 361222 685898 396986 686134
rect 397222 685898 432986 686134
rect 433222 685898 468986 686134
rect 469222 685898 504986 686134
rect 505222 685898 540986 686134
rect 541222 685898 576986 686134
rect 577222 685898 585502 686134
rect 585738 685898 586840 686134
rect -2916 685876 586840 685898
rect -1996 685874 -1396 685876
rect 804 685874 1404 685876
rect 36804 685874 37404 685876
rect 72804 685874 73404 685876
rect 108804 685874 109404 685876
rect 144804 685874 145404 685876
rect 180804 685874 181404 685876
rect 216804 685874 217404 685876
rect 252804 685874 253404 685876
rect 288804 685874 289404 685876
rect 324804 685874 325404 685876
rect 360804 685874 361404 685876
rect 396804 685874 397404 685876
rect 432804 685874 433404 685876
rect 468804 685874 469404 685876
rect 504804 685874 505404 685876
rect 540804 685874 541404 685876
rect 576804 685874 577404 685876
rect 585320 685874 585920 685876
rect -8436 679276 -7836 679278
rect 29604 679276 30204 679278
rect 65604 679276 66204 679278
rect 101604 679276 102204 679278
rect 137604 679276 138204 679278
rect 173604 679276 174204 679278
rect 209604 679276 210204 679278
rect 245604 679276 246204 679278
rect 281604 679276 282204 679278
rect 317604 679276 318204 679278
rect 353604 679276 354204 679278
rect 389604 679276 390204 679278
rect 425604 679276 426204 679278
rect 461604 679276 462204 679278
rect 497604 679276 498204 679278
rect 533604 679276 534204 679278
rect 569604 679276 570204 679278
rect 591760 679276 592360 679278
rect -8436 679254 592360 679276
rect -8436 679018 -8254 679254
rect -8018 679018 29786 679254
rect 30022 679018 65786 679254
rect 66022 679018 101786 679254
rect 102022 679018 137786 679254
rect 138022 679018 173786 679254
rect 174022 679018 209786 679254
rect 210022 679018 245786 679254
rect 246022 679018 281786 679254
rect 282022 679018 317786 679254
rect 318022 679018 353786 679254
rect 354022 679018 389786 679254
rect 390022 679018 425786 679254
rect 426022 679018 461786 679254
rect 462022 679018 497786 679254
rect 498022 679018 533786 679254
rect 534022 679018 569786 679254
rect 570022 679018 591942 679254
rect 592178 679018 592360 679254
rect -8436 678934 592360 679018
rect -8436 678698 -8254 678934
rect -8018 678698 29786 678934
rect 30022 678698 65786 678934
rect 66022 678698 101786 678934
rect 102022 678698 137786 678934
rect 138022 678698 173786 678934
rect 174022 678698 209786 678934
rect 210022 678698 245786 678934
rect 246022 678698 281786 678934
rect 282022 678698 317786 678934
rect 318022 678698 353786 678934
rect 354022 678698 389786 678934
rect 390022 678698 425786 678934
rect 426022 678698 461786 678934
rect 462022 678698 497786 678934
rect 498022 678698 533786 678934
rect 534022 678698 569786 678934
rect 570022 678698 591942 678934
rect 592178 678698 592360 678934
rect -8436 678676 592360 678698
rect -8436 678674 -7836 678676
rect 29604 678674 30204 678676
rect 65604 678674 66204 678676
rect 101604 678674 102204 678676
rect 137604 678674 138204 678676
rect 173604 678674 174204 678676
rect 209604 678674 210204 678676
rect 245604 678674 246204 678676
rect 281604 678674 282204 678676
rect 317604 678674 318204 678676
rect 353604 678674 354204 678676
rect 389604 678674 390204 678676
rect 425604 678674 426204 678676
rect 461604 678674 462204 678676
rect 497604 678674 498204 678676
rect 533604 678674 534204 678676
rect 569604 678674 570204 678676
rect 591760 678674 592360 678676
rect -6596 675676 -5996 675678
rect 26004 675676 26604 675678
rect 62004 675676 62604 675678
rect 98004 675676 98604 675678
rect 134004 675676 134604 675678
rect 170004 675676 170604 675678
rect 206004 675676 206604 675678
rect 242004 675676 242604 675678
rect 278004 675676 278604 675678
rect 314004 675676 314604 675678
rect 350004 675676 350604 675678
rect 386004 675676 386604 675678
rect 422004 675676 422604 675678
rect 458004 675676 458604 675678
rect 494004 675676 494604 675678
rect 530004 675676 530604 675678
rect 566004 675676 566604 675678
rect 589920 675676 590520 675678
rect -6596 675654 590520 675676
rect -6596 675418 -6414 675654
rect -6178 675418 26186 675654
rect 26422 675418 62186 675654
rect 62422 675418 98186 675654
rect 98422 675418 134186 675654
rect 134422 675418 170186 675654
rect 170422 675418 206186 675654
rect 206422 675418 242186 675654
rect 242422 675418 278186 675654
rect 278422 675418 314186 675654
rect 314422 675418 350186 675654
rect 350422 675418 386186 675654
rect 386422 675418 422186 675654
rect 422422 675418 458186 675654
rect 458422 675418 494186 675654
rect 494422 675418 530186 675654
rect 530422 675418 566186 675654
rect 566422 675418 590102 675654
rect 590338 675418 590520 675654
rect -6596 675334 590520 675418
rect -6596 675098 -6414 675334
rect -6178 675098 26186 675334
rect 26422 675098 62186 675334
rect 62422 675098 98186 675334
rect 98422 675098 134186 675334
rect 134422 675098 170186 675334
rect 170422 675098 206186 675334
rect 206422 675098 242186 675334
rect 242422 675098 278186 675334
rect 278422 675098 314186 675334
rect 314422 675098 350186 675334
rect 350422 675098 386186 675334
rect 386422 675098 422186 675334
rect 422422 675098 458186 675334
rect 458422 675098 494186 675334
rect 494422 675098 530186 675334
rect 530422 675098 566186 675334
rect 566422 675098 590102 675334
rect 590338 675098 590520 675334
rect -6596 675076 590520 675098
rect -6596 675074 -5996 675076
rect 26004 675074 26604 675076
rect 62004 675074 62604 675076
rect 98004 675074 98604 675076
rect 134004 675074 134604 675076
rect 170004 675074 170604 675076
rect 206004 675074 206604 675076
rect 242004 675074 242604 675076
rect 278004 675074 278604 675076
rect 314004 675074 314604 675076
rect 350004 675074 350604 675076
rect 386004 675074 386604 675076
rect 422004 675074 422604 675076
rect 458004 675074 458604 675076
rect 494004 675074 494604 675076
rect 530004 675074 530604 675076
rect 566004 675074 566604 675076
rect 589920 675074 590520 675076
rect -4756 672076 -4156 672078
rect 22404 672076 23004 672078
rect 58404 672076 59004 672078
rect 94404 672076 95004 672078
rect 130404 672076 131004 672078
rect 166404 672076 167004 672078
rect 202404 672076 203004 672078
rect 238404 672076 239004 672078
rect 274404 672076 275004 672078
rect 310404 672076 311004 672078
rect 346404 672076 347004 672078
rect 382404 672076 383004 672078
rect 418404 672076 419004 672078
rect 454404 672076 455004 672078
rect 490404 672076 491004 672078
rect 526404 672076 527004 672078
rect 562404 672076 563004 672078
rect 588080 672076 588680 672078
rect -4756 672054 588680 672076
rect -4756 671818 -4574 672054
rect -4338 671818 22586 672054
rect 22822 671818 58586 672054
rect 58822 671818 94586 672054
rect 94822 671818 130586 672054
rect 130822 671818 166586 672054
rect 166822 671818 202586 672054
rect 202822 671818 238586 672054
rect 238822 671818 274586 672054
rect 274822 671818 310586 672054
rect 310822 671818 346586 672054
rect 346822 671818 382586 672054
rect 382822 671818 418586 672054
rect 418822 671818 454586 672054
rect 454822 671818 490586 672054
rect 490822 671818 526586 672054
rect 526822 671818 562586 672054
rect 562822 671818 588262 672054
rect 588498 671818 588680 672054
rect -4756 671734 588680 671818
rect -4756 671498 -4574 671734
rect -4338 671498 22586 671734
rect 22822 671498 58586 671734
rect 58822 671498 94586 671734
rect 94822 671498 130586 671734
rect 130822 671498 166586 671734
rect 166822 671498 202586 671734
rect 202822 671498 238586 671734
rect 238822 671498 274586 671734
rect 274822 671498 310586 671734
rect 310822 671498 346586 671734
rect 346822 671498 382586 671734
rect 382822 671498 418586 671734
rect 418822 671498 454586 671734
rect 454822 671498 490586 671734
rect 490822 671498 526586 671734
rect 526822 671498 562586 671734
rect 562822 671498 588262 671734
rect 588498 671498 588680 671734
rect -4756 671476 588680 671498
rect -4756 671474 -4156 671476
rect 22404 671474 23004 671476
rect 58404 671474 59004 671476
rect 94404 671474 95004 671476
rect 130404 671474 131004 671476
rect 166404 671474 167004 671476
rect 202404 671474 203004 671476
rect 238404 671474 239004 671476
rect 274404 671474 275004 671476
rect 310404 671474 311004 671476
rect 346404 671474 347004 671476
rect 382404 671474 383004 671476
rect 418404 671474 419004 671476
rect 454404 671474 455004 671476
rect 490404 671474 491004 671476
rect 526404 671474 527004 671476
rect 562404 671474 563004 671476
rect 588080 671474 588680 671476
rect -2916 668476 -2316 668478
rect 18804 668476 19404 668478
rect 54804 668476 55404 668478
rect 90804 668476 91404 668478
rect 126804 668476 127404 668478
rect 162804 668476 163404 668478
rect 198804 668476 199404 668478
rect 234804 668476 235404 668478
rect 270804 668476 271404 668478
rect 306804 668476 307404 668478
rect 342804 668476 343404 668478
rect 378804 668476 379404 668478
rect 414804 668476 415404 668478
rect 450804 668476 451404 668478
rect 486804 668476 487404 668478
rect 522804 668476 523404 668478
rect 558804 668476 559404 668478
rect 586240 668476 586840 668478
rect -2916 668454 586840 668476
rect -2916 668218 -2734 668454
rect -2498 668218 18986 668454
rect 19222 668218 54986 668454
rect 55222 668218 90986 668454
rect 91222 668218 126986 668454
rect 127222 668218 162986 668454
rect 163222 668218 198986 668454
rect 199222 668218 234986 668454
rect 235222 668218 270986 668454
rect 271222 668218 306986 668454
rect 307222 668218 342986 668454
rect 343222 668218 378986 668454
rect 379222 668218 414986 668454
rect 415222 668218 450986 668454
rect 451222 668218 486986 668454
rect 487222 668218 522986 668454
rect 523222 668218 558986 668454
rect 559222 668218 586422 668454
rect 586658 668218 586840 668454
rect -2916 668134 586840 668218
rect -2916 667898 -2734 668134
rect -2498 667898 18986 668134
rect 19222 667898 54986 668134
rect 55222 667898 90986 668134
rect 91222 667898 126986 668134
rect 127222 667898 162986 668134
rect 163222 667898 198986 668134
rect 199222 667898 234986 668134
rect 235222 667898 270986 668134
rect 271222 667898 306986 668134
rect 307222 667898 342986 668134
rect 343222 667898 378986 668134
rect 379222 667898 414986 668134
rect 415222 667898 450986 668134
rect 451222 667898 486986 668134
rect 487222 667898 522986 668134
rect 523222 667898 558986 668134
rect 559222 667898 586422 668134
rect 586658 667898 586840 668134
rect -2916 667876 586840 667898
rect -2916 667874 -2316 667876
rect 18804 667874 19404 667876
rect 54804 667874 55404 667876
rect 90804 667874 91404 667876
rect 126804 667874 127404 667876
rect 162804 667874 163404 667876
rect 198804 667874 199404 667876
rect 234804 667874 235404 667876
rect 270804 667874 271404 667876
rect 306804 667874 307404 667876
rect 342804 667874 343404 667876
rect 378804 667874 379404 667876
rect 414804 667874 415404 667876
rect 450804 667874 451404 667876
rect 486804 667874 487404 667876
rect 522804 667874 523404 667876
rect 558804 667874 559404 667876
rect 586240 667874 586840 667876
rect -7516 661276 -6916 661278
rect 11604 661276 12204 661278
rect 47604 661276 48204 661278
rect 83604 661276 84204 661278
rect 119604 661276 120204 661278
rect 155604 661276 156204 661278
rect 191604 661276 192204 661278
rect 227604 661276 228204 661278
rect 263604 661276 264204 661278
rect 299604 661276 300204 661278
rect 335604 661276 336204 661278
rect 371604 661276 372204 661278
rect 407604 661276 408204 661278
rect 443604 661276 444204 661278
rect 479604 661276 480204 661278
rect 515604 661276 516204 661278
rect 551604 661276 552204 661278
rect 590840 661276 591440 661278
rect -8436 661254 592360 661276
rect -8436 661018 -7334 661254
rect -7098 661018 11786 661254
rect 12022 661018 47786 661254
rect 48022 661018 83786 661254
rect 84022 661018 119786 661254
rect 120022 661018 155786 661254
rect 156022 661018 191786 661254
rect 192022 661018 227786 661254
rect 228022 661018 263786 661254
rect 264022 661018 299786 661254
rect 300022 661018 335786 661254
rect 336022 661018 371786 661254
rect 372022 661018 407786 661254
rect 408022 661018 443786 661254
rect 444022 661018 479786 661254
rect 480022 661018 515786 661254
rect 516022 661018 551786 661254
rect 552022 661018 591022 661254
rect 591258 661018 592360 661254
rect -8436 660934 592360 661018
rect -8436 660698 -7334 660934
rect -7098 660698 11786 660934
rect 12022 660698 47786 660934
rect 48022 660698 83786 660934
rect 84022 660698 119786 660934
rect 120022 660698 155786 660934
rect 156022 660698 191786 660934
rect 192022 660698 227786 660934
rect 228022 660698 263786 660934
rect 264022 660698 299786 660934
rect 300022 660698 335786 660934
rect 336022 660698 371786 660934
rect 372022 660698 407786 660934
rect 408022 660698 443786 660934
rect 444022 660698 479786 660934
rect 480022 660698 515786 660934
rect 516022 660698 551786 660934
rect 552022 660698 591022 660934
rect 591258 660698 592360 660934
rect -8436 660676 592360 660698
rect -7516 660674 -6916 660676
rect 11604 660674 12204 660676
rect 47604 660674 48204 660676
rect 83604 660674 84204 660676
rect 119604 660674 120204 660676
rect 155604 660674 156204 660676
rect 191604 660674 192204 660676
rect 227604 660674 228204 660676
rect 263604 660674 264204 660676
rect 299604 660674 300204 660676
rect 335604 660674 336204 660676
rect 371604 660674 372204 660676
rect 407604 660674 408204 660676
rect 443604 660674 444204 660676
rect 479604 660674 480204 660676
rect 515604 660674 516204 660676
rect 551604 660674 552204 660676
rect 590840 660674 591440 660676
rect -5676 657676 -5076 657678
rect 8004 657676 8604 657678
rect 44004 657676 44604 657678
rect 80004 657676 80604 657678
rect 116004 657676 116604 657678
rect 152004 657676 152604 657678
rect 188004 657676 188604 657678
rect 224004 657676 224604 657678
rect 260004 657676 260604 657678
rect 296004 657676 296604 657678
rect 332004 657676 332604 657678
rect 368004 657676 368604 657678
rect 404004 657676 404604 657678
rect 440004 657676 440604 657678
rect 476004 657676 476604 657678
rect 512004 657676 512604 657678
rect 548004 657676 548604 657678
rect 589000 657676 589600 657678
rect -6596 657654 590520 657676
rect -6596 657418 -5494 657654
rect -5258 657418 8186 657654
rect 8422 657418 44186 657654
rect 44422 657418 80186 657654
rect 80422 657418 116186 657654
rect 116422 657418 152186 657654
rect 152422 657418 188186 657654
rect 188422 657418 224186 657654
rect 224422 657418 260186 657654
rect 260422 657418 296186 657654
rect 296422 657418 332186 657654
rect 332422 657418 368186 657654
rect 368422 657418 404186 657654
rect 404422 657418 440186 657654
rect 440422 657418 476186 657654
rect 476422 657418 512186 657654
rect 512422 657418 548186 657654
rect 548422 657418 589182 657654
rect 589418 657418 590520 657654
rect -6596 657334 590520 657418
rect -6596 657098 -5494 657334
rect -5258 657098 8186 657334
rect 8422 657098 44186 657334
rect 44422 657098 80186 657334
rect 80422 657098 116186 657334
rect 116422 657098 152186 657334
rect 152422 657098 188186 657334
rect 188422 657098 224186 657334
rect 224422 657098 260186 657334
rect 260422 657098 296186 657334
rect 296422 657098 332186 657334
rect 332422 657098 368186 657334
rect 368422 657098 404186 657334
rect 404422 657098 440186 657334
rect 440422 657098 476186 657334
rect 476422 657098 512186 657334
rect 512422 657098 548186 657334
rect 548422 657098 589182 657334
rect 589418 657098 590520 657334
rect -6596 657076 590520 657098
rect -5676 657074 -5076 657076
rect 8004 657074 8604 657076
rect 44004 657074 44604 657076
rect 80004 657074 80604 657076
rect 116004 657074 116604 657076
rect 152004 657074 152604 657076
rect 188004 657074 188604 657076
rect 224004 657074 224604 657076
rect 260004 657074 260604 657076
rect 296004 657074 296604 657076
rect 332004 657074 332604 657076
rect 368004 657074 368604 657076
rect 404004 657074 404604 657076
rect 440004 657074 440604 657076
rect 476004 657074 476604 657076
rect 512004 657074 512604 657076
rect 548004 657074 548604 657076
rect 589000 657074 589600 657076
rect -3836 654076 -3236 654078
rect 4404 654076 5004 654078
rect 40404 654076 41004 654078
rect 76404 654076 77004 654078
rect 112404 654076 113004 654078
rect 148404 654076 149004 654078
rect 184404 654076 185004 654078
rect 220404 654076 221004 654078
rect 256404 654076 257004 654078
rect 292404 654076 293004 654078
rect 328404 654076 329004 654078
rect 364404 654076 365004 654078
rect 400404 654076 401004 654078
rect 436404 654076 437004 654078
rect 472404 654076 473004 654078
rect 508404 654076 509004 654078
rect 544404 654076 545004 654078
rect 580404 654076 581004 654078
rect 587160 654076 587760 654078
rect -4756 654054 588680 654076
rect -4756 653818 -3654 654054
rect -3418 653818 4586 654054
rect 4822 653818 40586 654054
rect 40822 653818 76586 654054
rect 76822 653818 112586 654054
rect 112822 653818 148586 654054
rect 148822 653818 184586 654054
rect 184822 653818 220586 654054
rect 220822 653818 256586 654054
rect 256822 653818 292586 654054
rect 292822 653818 328586 654054
rect 328822 653818 364586 654054
rect 364822 653818 400586 654054
rect 400822 653818 436586 654054
rect 436822 653818 472586 654054
rect 472822 653818 508586 654054
rect 508822 653818 544586 654054
rect 544822 653818 580586 654054
rect 580822 653818 587342 654054
rect 587578 653818 588680 654054
rect -4756 653734 588680 653818
rect -4756 653498 -3654 653734
rect -3418 653498 4586 653734
rect 4822 653498 40586 653734
rect 40822 653498 76586 653734
rect 76822 653498 112586 653734
rect 112822 653498 148586 653734
rect 148822 653498 184586 653734
rect 184822 653498 220586 653734
rect 220822 653498 256586 653734
rect 256822 653498 292586 653734
rect 292822 653498 328586 653734
rect 328822 653498 364586 653734
rect 364822 653498 400586 653734
rect 400822 653498 436586 653734
rect 436822 653498 472586 653734
rect 472822 653498 508586 653734
rect 508822 653498 544586 653734
rect 544822 653498 580586 653734
rect 580822 653498 587342 653734
rect 587578 653498 588680 653734
rect -4756 653476 588680 653498
rect -3836 653474 -3236 653476
rect 4404 653474 5004 653476
rect 40404 653474 41004 653476
rect 76404 653474 77004 653476
rect 112404 653474 113004 653476
rect 148404 653474 149004 653476
rect 184404 653474 185004 653476
rect 220404 653474 221004 653476
rect 256404 653474 257004 653476
rect 292404 653474 293004 653476
rect 328404 653474 329004 653476
rect 364404 653474 365004 653476
rect 400404 653474 401004 653476
rect 436404 653474 437004 653476
rect 472404 653474 473004 653476
rect 508404 653474 509004 653476
rect 544404 653474 545004 653476
rect 580404 653474 581004 653476
rect 587160 653474 587760 653476
rect -1996 650476 -1396 650478
rect 804 650476 1404 650478
rect 36804 650476 37404 650478
rect 72804 650476 73404 650478
rect 108804 650476 109404 650478
rect 144804 650476 145404 650478
rect 180804 650476 181404 650478
rect 216804 650476 217404 650478
rect 252804 650476 253404 650478
rect 288804 650476 289404 650478
rect 324804 650476 325404 650478
rect 360804 650476 361404 650478
rect 396804 650476 397404 650478
rect 432804 650476 433404 650478
rect 468804 650476 469404 650478
rect 504804 650476 505404 650478
rect 540804 650476 541404 650478
rect 576804 650476 577404 650478
rect 585320 650476 585920 650478
rect -2916 650454 586840 650476
rect -2916 650218 -1814 650454
rect -1578 650218 986 650454
rect 1222 650218 36986 650454
rect 37222 650218 72986 650454
rect 73222 650218 108986 650454
rect 109222 650218 144986 650454
rect 145222 650218 180986 650454
rect 181222 650218 216986 650454
rect 217222 650218 252986 650454
rect 253222 650218 288986 650454
rect 289222 650218 324986 650454
rect 325222 650218 360986 650454
rect 361222 650218 396986 650454
rect 397222 650218 432986 650454
rect 433222 650218 468986 650454
rect 469222 650218 504986 650454
rect 505222 650218 540986 650454
rect 541222 650218 576986 650454
rect 577222 650218 585502 650454
rect 585738 650218 586840 650454
rect -2916 650134 586840 650218
rect -2916 649898 -1814 650134
rect -1578 649898 986 650134
rect 1222 649898 36986 650134
rect 37222 649898 72986 650134
rect 73222 649898 108986 650134
rect 109222 649898 144986 650134
rect 145222 649898 180986 650134
rect 181222 649898 216986 650134
rect 217222 649898 252986 650134
rect 253222 649898 288986 650134
rect 289222 649898 324986 650134
rect 325222 649898 360986 650134
rect 361222 649898 396986 650134
rect 397222 649898 432986 650134
rect 433222 649898 468986 650134
rect 469222 649898 504986 650134
rect 505222 649898 540986 650134
rect 541222 649898 576986 650134
rect 577222 649898 585502 650134
rect 585738 649898 586840 650134
rect -2916 649876 586840 649898
rect -1996 649874 -1396 649876
rect 804 649874 1404 649876
rect 36804 649874 37404 649876
rect 72804 649874 73404 649876
rect 108804 649874 109404 649876
rect 144804 649874 145404 649876
rect 180804 649874 181404 649876
rect 216804 649874 217404 649876
rect 252804 649874 253404 649876
rect 288804 649874 289404 649876
rect 324804 649874 325404 649876
rect 360804 649874 361404 649876
rect 396804 649874 397404 649876
rect 432804 649874 433404 649876
rect 468804 649874 469404 649876
rect 504804 649874 505404 649876
rect 540804 649874 541404 649876
rect 576804 649874 577404 649876
rect 585320 649874 585920 649876
rect -8436 643276 -7836 643278
rect 29604 643276 30204 643278
rect 65604 643276 66204 643278
rect 101604 643276 102204 643278
rect 137604 643276 138204 643278
rect 173604 643276 174204 643278
rect 209604 643276 210204 643278
rect 245604 643276 246204 643278
rect 281604 643276 282204 643278
rect 317604 643276 318204 643278
rect 353604 643276 354204 643278
rect 389604 643276 390204 643278
rect 425604 643276 426204 643278
rect 461604 643276 462204 643278
rect 497604 643276 498204 643278
rect 533604 643276 534204 643278
rect 569604 643276 570204 643278
rect 591760 643276 592360 643278
rect -8436 643254 592360 643276
rect -8436 643018 -8254 643254
rect -8018 643018 29786 643254
rect 30022 643018 65786 643254
rect 66022 643018 101786 643254
rect 102022 643018 137786 643254
rect 138022 643018 173786 643254
rect 174022 643018 209786 643254
rect 210022 643018 245786 643254
rect 246022 643018 281786 643254
rect 282022 643018 317786 643254
rect 318022 643018 353786 643254
rect 354022 643018 389786 643254
rect 390022 643018 425786 643254
rect 426022 643018 461786 643254
rect 462022 643018 497786 643254
rect 498022 643018 533786 643254
rect 534022 643018 569786 643254
rect 570022 643018 591942 643254
rect 592178 643018 592360 643254
rect -8436 642934 592360 643018
rect -8436 642698 -8254 642934
rect -8018 642698 29786 642934
rect 30022 642698 65786 642934
rect 66022 642698 101786 642934
rect 102022 642698 137786 642934
rect 138022 642698 173786 642934
rect 174022 642698 209786 642934
rect 210022 642698 245786 642934
rect 246022 642698 281786 642934
rect 282022 642698 317786 642934
rect 318022 642698 353786 642934
rect 354022 642698 389786 642934
rect 390022 642698 425786 642934
rect 426022 642698 461786 642934
rect 462022 642698 497786 642934
rect 498022 642698 533786 642934
rect 534022 642698 569786 642934
rect 570022 642698 591942 642934
rect 592178 642698 592360 642934
rect -8436 642676 592360 642698
rect -8436 642674 -7836 642676
rect 29604 642674 30204 642676
rect 65604 642674 66204 642676
rect 101604 642674 102204 642676
rect 137604 642674 138204 642676
rect 173604 642674 174204 642676
rect 209604 642674 210204 642676
rect 245604 642674 246204 642676
rect 281604 642674 282204 642676
rect 317604 642674 318204 642676
rect 353604 642674 354204 642676
rect 389604 642674 390204 642676
rect 425604 642674 426204 642676
rect 461604 642674 462204 642676
rect 497604 642674 498204 642676
rect 533604 642674 534204 642676
rect 569604 642674 570204 642676
rect 591760 642674 592360 642676
rect -6596 639676 -5996 639678
rect 26004 639676 26604 639678
rect 62004 639676 62604 639678
rect 98004 639676 98604 639678
rect 134004 639676 134604 639678
rect 170004 639676 170604 639678
rect 206004 639676 206604 639678
rect 242004 639676 242604 639678
rect 278004 639676 278604 639678
rect 314004 639676 314604 639678
rect 350004 639676 350604 639678
rect 386004 639676 386604 639678
rect 422004 639676 422604 639678
rect 458004 639676 458604 639678
rect 494004 639676 494604 639678
rect 530004 639676 530604 639678
rect 566004 639676 566604 639678
rect 589920 639676 590520 639678
rect -6596 639654 590520 639676
rect -6596 639418 -6414 639654
rect -6178 639418 26186 639654
rect 26422 639418 62186 639654
rect 62422 639418 98186 639654
rect 98422 639418 134186 639654
rect 134422 639418 170186 639654
rect 170422 639418 206186 639654
rect 206422 639418 242186 639654
rect 242422 639418 278186 639654
rect 278422 639418 314186 639654
rect 314422 639418 350186 639654
rect 350422 639418 386186 639654
rect 386422 639418 422186 639654
rect 422422 639418 458186 639654
rect 458422 639418 494186 639654
rect 494422 639418 530186 639654
rect 530422 639418 566186 639654
rect 566422 639418 590102 639654
rect 590338 639418 590520 639654
rect -6596 639334 590520 639418
rect -6596 639098 -6414 639334
rect -6178 639098 26186 639334
rect 26422 639098 62186 639334
rect 62422 639098 98186 639334
rect 98422 639098 134186 639334
rect 134422 639098 170186 639334
rect 170422 639098 206186 639334
rect 206422 639098 242186 639334
rect 242422 639098 278186 639334
rect 278422 639098 314186 639334
rect 314422 639098 350186 639334
rect 350422 639098 386186 639334
rect 386422 639098 422186 639334
rect 422422 639098 458186 639334
rect 458422 639098 494186 639334
rect 494422 639098 530186 639334
rect 530422 639098 566186 639334
rect 566422 639098 590102 639334
rect 590338 639098 590520 639334
rect -6596 639076 590520 639098
rect -6596 639074 -5996 639076
rect 26004 639074 26604 639076
rect 62004 639074 62604 639076
rect 98004 639074 98604 639076
rect 134004 639074 134604 639076
rect 170004 639074 170604 639076
rect 206004 639074 206604 639076
rect 242004 639074 242604 639076
rect 278004 639074 278604 639076
rect 314004 639074 314604 639076
rect 350004 639074 350604 639076
rect 386004 639074 386604 639076
rect 422004 639074 422604 639076
rect 458004 639074 458604 639076
rect 494004 639074 494604 639076
rect 530004 639074 530604 639076
rect 566004 639074 566604 639076
rect 589920 639074 590520 639076
rect -4756 636076 -4156 636078
rect 22404 636076 23004 636078
rect 58404 636076 59004 636078
rect 94404 636076 95004 636078
rect 130404 636076 131004 636078
rect 166404 636076 167004 636078
rect 202404 636076 203004 636078
rect 238404 636076 239004 636078
rect 274404 636076 275004 636078
rect 310404 636076 311004 636078
rect 346404 636076 347004 636078
rect 382404 636076 383004 636078
rect 418404 636076 419004 636078
rect 454404 636076 455004 636078
rect 490404 636076 491004 636078
rect 526404 636076 527004 636078
rect 562404 636076 563004 636078
rect 588080 636076 588680 636078
rect -4756 636054 588680 636076
rect -4756 635818 -4574 636054
rect -4338 635818 22586 636054
rect 22822 635818 58586 636054
rect 58822 635818 94586 636054
rect 94822 635818 130586 636054
rect 130822 635818 166586 636054
rect 166822 635818 202586 636054
rect 202822 635818 238586 636054
rect 238822 635818 274586 636054
rect 274822 635818 310586 636054
rect 310822 635818 346586 636054
rect 346822 635818 382586 636054
rect 382822 635818 418586 636054
rect 418822 635818 454586 636054
rect 454822 635818 490586 636054
rect 490822 635818 526586 636054
rect 526822 635818 562586 636054
rect 562822 635818 588262 636054
rect 588498 635818 588680 636054
rect -4756 635734 588680 635818
rect -4756 635498 -4574 635734
rect -4338 635498 22586 635734
rect 22822 635498 58586 635734
rect 58822 635498 94586 635734
rect 94822 635498 130586 635734
rect 130822 635498 166586 635734
rect 166822 635498 202586 635734
rect 202822 635498 238586 635734
rect 238822 635498 274586 635734
rect 274822 635498 310586 635734
rect 310822 635498 346586 635734
rect 346822 635498 382586 635734
rect 382822 635498 418586 635734
rect 418822 635498 454586 635734
rect 454822 635498 490586 635734
rect 490822 635498 526586 635734
rect 526822 635498 562586 635734
rect 562822 635498 588262 635734
rect 588498 635498 588680 635734
rect -4756 635476 588680 635498
rect -4756 635474 -4156 635476
rect 22404 635474 23004 635476
rect 58404 635474 59004 635476
rect 94404 635474 95004 635476
rect 130404 635474 131004 635476
rect 166404 635474 167004 635476
rect 202404 635474 203004 635476
rect 238404 635474 239004 635476
rect 274404 635474 275004 635476
rect 310404 635474 311004 635476
rect 346404 635474 347004 635476
rect 382404 635474 383004 635476
rect 418404 635474 419004 635476
rect 454404 635474 455004 635476
rect 490404 635474 491004 635476
rect 526404 635474 527004 635476
rect 562404 635474 563004 635476
rect 588080 635474 588680 635476
rect -2916 632476 -2316 632478
rect 18804 632476 19404 632478
rect 54804 632476 55404 632478
rect 90804 632476 91404 632478
rect 126804 632476 127404 632478
rect 162804 632476 163404 632478
rect 198804 632476 199404 632478
rect 234804 632476 235404 632478
rect 270804 632476 271404 632478
rect 306804 632476 307404 632478
rect 342804 632476 343404 632478
rect 378804 632476 379404 632478
rect 414804 632476 415404 632478
rect 450804 632476 451404 632478
rect 486804 632476 487404 632478
rect 522804 632476 523404 632478
rect 558804 632476 559404 632478
rect 586240 632476 586840 632478
rect -2916 632454 586840 632476
rect -2916 632218 -2734 632454
rect -2498 632218 18986 632454
rect 19222 632218 54986 632454
rect 55222 632218 90986 632454
rect 91222 632218 126986 632454
rect 127222 632218 162986 632454
rect 163222 632218 198986 632454
rect 199222 632218 234986 632454
rect 235222 632218 270986 632454
rect 271222 632218 306986 632454
rect 307222 632218 342986 632454
rect 343222 632218 378986 632454
rect 379222 632218 414986 632454
rect 415222 632218 450986 632454
rect 451222 632218 486986 632454
rect 487222 632218 522986 632454
rect 523222 632218 558986 632454
rect 559222 632218 586422 632454
rect 586658 632218 586840 632454
rect -2916 632134 586840 632218
rect -2916 631898 -2734 632134
rect -2498 631898 18986 632134
rect 19222 631898 54986 632134
rect 55222 631898 90986 632134
rect 91222 631898 126986 632134
rect 127222 631898 162986 632134
rect 163222 631898 198986 632134
rect 199222 631898 234986 632134
rect 235222 631898 270986 632134
rect 271222 631898 306986 632134
rect 307222 631898 342986 632134
rect 343222 631898 378986 632134
rect 379222 631898 414986 632134
rect 415222 631898 450986 632134
rect 451222 631898 486986 632134
rect 487222 631898 522986 632134
rect 523222 631898 558986 632134
rect 559222 631898 586422 632134
rect 586658 631898 586840 632134
rect -2916 631876 586840 631898
rect -2916 631874 -2316 631876
rect 18804 631874 19404 631876
rect 54804 631874 55404 631876
rect 90804 631874 91404 631876
rect 126804 631874 127404 631876
rect 162804 631874 163404 631876
rect 198804 631874 199404 631876
rect 234804 631874 235404 631876
rect 270804 631874 271404 631876
rect 306804 631874 307404 631876
rect 342804 631874 343404 631876
rect 378804 631874 379404 631876
rect 414804 631874 415404 631876
rect 450804 631874 451404 631876
rect 486804 631874 487404 631876
rect 522804 631874 523404 631876
rect 558804 631874 559404 631876
rect 586240 631874 586840 631876
rect -7516 625276 -6916 625278
rect 11604 625276 12204 625278
rect 47604 625276 48204 625278
rect 83604 625276 84204 625278
rect 119604 625276 120204 625278
rect 155604 625276 156204 625278
rect 191604 625276 192204 625278
rect 227604 625276 228204 625278
rect 263604 625276 264204 625278
rect 299604 625276 300204 625278
rect 335604 625276 336204 625278
rect 371604 625276 372204 625278
rect 407604 625276 408204 625278
rect 443604 625276 444204 625278
rect 479604 625276 480204 625278
rect 515604 625276 516204 625278
rect 551604 625276 552204 625278
rect 590840 625276 591440 625278
rect -8436 625254 592360 625276
rect -8436 625018 -7334 625254
rect -7098 625018 11786 625254
rect 12022 625018 47786 625254
rect 48022 625018 83786 625254
rect 84022 625018 119786 625254
rect 120022 625018 155786 625254
rect 156022 625018 191786 625254
rect 192022 625018 227786 625254
rect 228022 625018 263786 625254
rect 264022 625018 299786 625254
rect 300022 625018 335786 625254
rect 336022 625018 371786 625254
rect 372022 625018 407786 625254
rect 408022 625018 443786 625254
rect 444022 625018 479786 625254
rect 480022 625018 515786 625254
rect 516022 625018 551786 625254
rect 552022 625018 591022 625254
rect 591258 625018 592360 625254
rect -8436 624934 592360 625018
rect -8436 624698 -7334 624934
rect -7098 624698 11786 624934
rect 12022 624698 47786 624934
rect 48022 624698 83786 624934
rect 84022 624698 119786 624934
rect 120022 624698 155786 624934
rect 156022 624698 191786 624934
rect 192022 624698 227786 624934
rect 228022 624698 263786 624934
rect 264022 624698 299786 624934
rect 300022 624698 335786 624934
rect 336022 624698 371786 624934
rect 372022 624698 407786 624934
rect 408022 624698 443786 624934
rect 444022 624698 479786 624934
rect 480022 624698 515786 624934
rect 516022 624698 551786 624934
rect 552022 624698 591022 624934
rect 591258 624698 592360 624934
rect -8436 624676 592360 624698
rect -7516 624674 -6916 624676
rect 11604 624674 12204 624676
rect 47604 624674 48204 624676
rect 83604 624674 84204 624676
rect 119604 624674 120204 624676
rect 155604 624674 156204 624676
rect 191604 624674 192204 624676
rect 227604 624674 228204 624676
rect 263604 624674 264204 624676
rect 299604 624674 300204 624676
rect 335604 624674 336204 624676
rect 371604 624674 372204 624676
rect 407604 624674 408204 624676
rect 443604 624674 444204 624676
rect 479604 624674 480204 624676
rect 515604 624674 516204 624676
rect 551604 624674 552204 624676
rect 590840 624674 591440 624676
rect -5676 621676 -5076 621678
rect 8004 621676 8604 621678
rect 44004 621676 44604 621678
rect 80004 621676 80604 621678
rect 116004 621676 116604 621678
rect 152004 621676 152604 621678
rect 188004 621676 188604 621678
rect 224004 621676 224604 621678
rect 260004 621676 260604 621678
rect 296004 621676 296604 621678
rect 332004 621676 332604 621678
rect 368004 621676 368604 621678
rect 404004 621676 404604 621678
rect 440004 621676 440604 621678
rect 476004 621676 476604 621678
rect 512004 621676 512604 621678
rect 548004 621676 548604 621678
rect 589000 621676 589600 621678
rect -6596 621654 590520 621676
rect -6596 621418 -5494 621654
rect -5258 621418 8186 621654
rect 8422 621418 44186 621654
rect 44422 621418 80186 621654
rect 80422 621418 116186 621654
rect 116422 621418 152186 621654
rect 152422 621418 188186 621654
rect 188422 621418 224186 621654
rect 224422 621418 260186 621654
rect 260422 621418 296186 621654
rect 296422 621418 332186 621654
rect 332422 621418 368186 621654
rect 368422 621418 404186 621654
rect 404422 621418 440186 621654
rect 440422 621418 476186 621654
rect 476422 621418 512186 621654
rect 512422 621418 548186 621654
rect 548422 621418 589182 621654
rect 589418 621418 590520 621654
rect -6596 621334 590520 621418
rect -6596 621098 -5494 621334
rect -5258 621098 8186 621334
rect 8422 621098 44186 621334
rect 44422 621098 80186 621334
rect 80422 621098 116186 621334
rect 116422 621098 152186 621334
rect 152422 621098 188186 621334
rect 188422 621098 224186 621334
rect 224422 621098 260186 621334
rect 260422 621098 296186 621334
rect 296422 621098 332186 621334
rect 332422 621098 368186 621334
rect 368422 621098 404186 621334
rect 404422 621098 440186 621334
rect 440422 621098 476186 621334
rect 476422 621098 512186 621334
rect 512422 621098 548186 621334
rect 548422 621098 589182 621334
rect 589418 621098 590520 621334
rect -6596 621076 590520 621098
rect -5676 621074 -5076 621076
rect 8004 621074 8604 621076
rect 44004 621074 44604 621076
rect 80004 621074 80604 621076
rect 116004 621074 116604 621076
rect 152004 621074 152604 621076
rect 188004 621074 188604 621076
rect 224004 621074 224604 621076
rect 260004 621074 260604 621076
rect 296004 621074 296604 621076
rect 332004 621074 332604 621076
rect 368004 621074 368604 621076
rect 404004 621074 404604 621076
rect 440004 621074 440604 621076
rect 476004 621074 476604 621076
rect 512004 621074 512604 621076
rect 548004 621074 548604 621076
rect 589000 621074 589600 621076
rect -3836 618076 -3236 618078
rect 4404 618076 5004 618078
rect 40404 618076 41004 618078
rect 76404 618076 77004 618078
rect 112404 618076 113004 618078
rect 148404 618076 149004 618078
rect 184404 618076 185004 618078
rect 220404 618076 221004 618078
rect 256404 618076 257004 618078
rect 292404 618076 293004 618078
rect 328404 618076 329004 618078
rect 364404 618076 365004 618078
rect 400404 618076 401004 618078
rect 436404 618076 437004 618078
rect 472404 618076 473004 618078
rect 508404 618076 509004 618078
rect 544404 618076 545004 618078
rect 580404 618076 581004 618078
rect 587160 618076 587760 618078
rect -4756 618054 588680 618076
rect -4756 617818 -3654 618054
rect -3418 617818 4586 618054
rect 4822 617818 40586 618054
rect 40822 617818 76586 618054
rect 76822 617818 112586 618054
rect 112822 617818 148586 618054
rect 148822 617818 184586 618054
rect 184822 617818 220586 618054
rect 220822 617818 256586 618054
rect 256822 617818 292586 618054
rect 292822 617818 328586 618054
rect 328822 617818 364586 618054
rect 364822 617818 400586 618054
rect 400822 617818 436586 618054
rect 436822 617818 472586 618054
rect 472822 617818 508586 618054
rect 508822 617818 544586 618054
rect 544822 617818 580586 618054
rect 580822 617818 587342 618054
rect 587578 617818 588680 618054
rect -4756 617734 588680 617818
rect -4756 617498 -3654 617734
rect -3418 617498 4586 617734
rect 4822 617498 40586 617734
rect 40822 617498 76586 617734
rect 76822 617498 112586 617734
rect 112822 617498 148586 617734
rect 148822 617498 184586 617734
rect 184822 617498 220586 617734
rect 220822 617498 256586 617734
rect 256822 617498 292586 617734
rect 292822 617498 328586 617734
rect 328822 617498 364586 617734
rect 364822 617498 400586 617734
rect 400822 617498 436586 617734
rect 436822 617498 472586 617734
rect 472822 617498 508586 617734
rect 508822 617498 544586 617734
rect 544822 617498 580586 617734
rect 580822 617498 587342 617734
rect 587578 617498 588680 617734
rect -4756 617476 588680 617498
rect -3836 617474 -3236 617476
rect 4404 617474 5004 617476
rect 40404 617474 41004 617476
rect 76404 617474 77004 617476
rect 112404 617474 113004 617476
rect 148404 617474 149004 617476
rect 184404 617474 185004 617476
rect 220404 617474 221004 617476
rect 256404 617474 257004 617476
rect 292404 617474 293004 617476
rect 328404 617474 329004 617476
rect 364404 617474 365004 617476
rect 400404 617474 401004 617476
rect 436404 617474 437004 617476
rect 472404 617474 473004 617476
rect 508404 617474 509004 617476
rect 544404 617474 545004 617476
rect 580404 617474 581004 617476
rect 587160 617474 587760 617476
rect -1996 614476 -1396 614478
rect 804 614476 1404 614478
rect 36804 614476 37404 614478
rect 72804 614476 73404 614478
rect 108804 614476 109404 614478
rect 144804 614476 145404 614478
rect 180804 614476 181404 614478
rect 216804 614476 217404 614478
rect 252804 614476 253404 614478
rect 288804 614476 289404 614478
rect 324804 614476 325404 614478
rect 360804 614476 361404 614478
rect 396804 614476 397404 614478
rect 432804 614476 433404 614478
rect 468804 614476 469404 614478
rect 504804 614476 505404 614478
rect 540804 614476 541404 614478
rect 576804 614476 577404 614478
rect 585320 614476 585920 614478
rect -2916 614454 586840 614476
rect -2916 614218 -1814 614454
rect -1578 614218 986 614454
rect 1222 614218 36986 614454
rect 37222 614218 72986 614454
rect 73222 614218 108986 614454
rect 109222 614218 144986 614454
rect 145222 614218 180986 614454
rect 181222 614218 216986 614454
rect 217222 614218 252986 614454
rect 253222 614218 288986 614454
rect 289222 614218 324986 614454
rect 325222 614218 360986 614454
rect 361222 614218 396986 614454
rect 397222 614218 432986 614454
rect 433222 614218 468986 614454
rect 469222 614218 504986 614454
rect 505222 614218 540986 614454
rect 541222 614218 576986 614454
rect 577222 614218 585502 614454
rect 585738 614218 586840 614454
rect -2916 614134 586840 614218
rect -2916 613898 -1814 614134
rect -1578 613898 986 614134
rect 1222 613898 36986 614134
rect 37222 613898 72986 614134
rect 73222 613898 108986 614134
rect 109222 613898 144986 614134
rect 145222 613898 180986 614134
rect 181222 613898 216986 614134
rect 217222 613898 252986 614134
rect 253222 613898 288986 614134
rect 289222 613898 324986 614134
rect 325222 613898 360986 614134
rect 361222 613898 396986 614134
rect 397222 613898 432986 614134
rect 433222 613898 468986 614134
rect 469222 613898 504986 614134
rect 505222 613898 540986 614134
rect 541222 613898 576986 614134
rect 577222 613898 585502 614134
rect 585738 613898 586840 614134
rect -2916 613876 586840 613898
rect -1996 613874 -1396 613876
rect 804 613874 1404 613876
rect 36804 613874 37404 613876
rect 72804 613874 73404 613876
rect 108804 613874 109404 613876
rect 144804 613874 145404 613876
rect 180804 613874 181404 613876
rect 216804 613874 217404 613876
rect 252804 613874 253404 613876
rect 288804 613874 289404 613876
rect 324804 613874 325404 613876
rect 360804 613874 361404 613876
rect 396804 613874 397404 613876
rect 432804 613874 433404 613876
rect 468804 613874 469404 613876
rect 504804 613874 505404 613876
rect 540804 613874 541404 613876
rect 576804 613874 577404 613876
rect 585320 613874 585920 613876
rect -8436 607276 -7836 607278
rect 29604 607276 30204 607278
rect 65604 607276 66204 607278
rect 101604 607276 102204 607278
rect 137604 607276 138204 607278
rect 173604 607276 174204 607278
rect 209604 607276 210204 607278
rect 245604 607276 246204 607278
rect 281604 607276 282204 607278
rect 317604 607276 318204 607278
rect 353604 607276 354204 607278
rect 389604 607276 390204 607278
rect 425604 607276 426204 607278
rect 461604 607276 462204 607278
rect 497604 607276 498204 607278
rect 533604 607276 534204 607278
rect 569604 607276 570204 607278
rect 591760 607276 592360 607278
rect -8436 607254 592360 607276
rect -8436 607018 -8254 607254
rect -8018 607018 29786 607254
rect 30022 607018 65786 607254
rect 66022 607018 101786 607254
rect 102022 607018 137786 607254
rect 138022 607018 173786 607254
rect 174022 607018 209786 607254
rect 210022 607018 245786 607254
rect 246022 607018 281786 607254
rect 282022 607018 317786 607254
rect 318022 607018 353786 607254
rect 354022 607018 389786 607254
rect 390022 607018 425786 607254
rect 426022 607018 461786 607254
rect 462022 607018 497786 607254
rect 498022 607018 533786 607254
rect 534022 607018 569786 607254
rect 570022 607018 591942 607254
rect 592178 607018 592360 607254
rect -8436 606934 592360 607018
rect -8436 606698 -8254 606934
rect -8018 606698 29786 606934
rect 30022 606698 65786 606934
rect 66022 606698 101786 606934
rect 102022 606698 137786 606934
rect 138022 606698 173786 606934
rect 174022 606698 209786 606934
rect 210022 606698 245786 606934
rect 246022 606698 281786 606934
rect 282022 606698 317786 606934
rect 318022 606698 353786 606934
rect 354022 606698 389786 606934
rect 390022 606698 425786 606934
rect 426022 606698 461786 606934
rect 462022 606698 497786 606934
rect 498022 606698 533786 606934
rect 534022 606698 569786 606934
rect 570022 606698 591942 606934
rect 592178 606698 592360 606934
rect -8436 606676 592360 606698
rect -8436 606674 -7836 606676
rect 29604 606674 30204 606676
rect 65604 606674 66204 606676
rect 101604 606674 102204 606676
rect 137604 606674 138204 606676
rect 173604 606674 174204 606676
rect 209604 606674 210204 606676
rect 245604 606674 246204 606676
rect 281604 606674 282204 606676
rect 317604 606674 318204 606676
rect 353604 606674 354204 606676
rect 389604 606674 390204 606676
rect 425604 606674 426204 606676
rect 461604 606674 462204 606676
rect 497604 606674 498204 606676
rect 533604 606674 534204 606676
rect 569604 606674 570204 606676
rect 591760 606674 592360 606676
rect -6596 603676 -5996 603678
rect 26004 603676 26604 603678
rect 62004 603676 62604 603678
rect 98004 603676 98604 603678
rect 134004 603676 134604 603678
rect 170004 603676 170604 603678
rect 206004 603676 206604 603678
rect 242004 603676 242604 603678
rect 278004 603676 278604 603678
rect 314004 603676 314604 603678
rect 350004 603676 350604 603678
rect 386004 603676 386604 603678
rect 422004 603676 422604 603678
rect 458004 603676 458604 603678
rect 494004 603676 494604 603678
rect 530004 603676 530604 603678
rect 566004 603676 566604 603678
rect 589920 603676 590520 603678
rect -6596 603654 590520 603676
rect -6596 603418 -6414 603654
rect -6178 603418 26186 603654
rect 26422 603418 62186 603654
rect 62422 603418 98186 603654
rect 98422 603418 134186 603654
rect 134422 603418 170186 603654
rect 170422 603418 206186 603654
rect 206422 603418 242186 603654
rect 242422 603418 278186 603654
rect 278422 603418 314186 603654
rect 314422 603418 350186 603654
rect 350422 603418 386186 603654
rect 386422 603418 422186 603654
rect 422422 603418 458186 603654
rect 458422 603418 494186 603654
rect 494422 603418 530186 603654
rect 530422 603418 566186 603654
rect 566422 603418 590102 603654
rect 590338 603418 590520 603654
rect -6596 603334 590520 603418
rect -6596 603098 -6414 603334
rect -6178 603098 26186 603334
rect 26422 603098 62186 603334
rect 62422 603098 98186 603334
rect 98422 603098 134186 603334
rect 134422 603098 170186 603334
rect 170422 603098 206186 603334
rect 206422 603098 242186 603334
rect 242422 603098 278186 603334
rect 278422 603098 314186 603334
rect 314422 603098 350186 603334
rect 350422 603098 386186 603334
rect 386422 603098 422186 603334
rect 422422 603098 458186 603334
rect 458422 603098 494186 603334
rect 494422 603098 530186 603334
rect 530422 603098 566186 603334
rect 566422 603098 590102 603334
rect 590338 603098 590520 603334
rect -6596 603076 590520 603098
rect -6596 603074 -5996 603076
rect 26004 603074 26604 603076
rect 62004 603074 62604 603076
rect 98004 603074 98604 603076
rect 134004 603074 134604 603076
rect 170004 603074 170604 603076
rect 206004 603074 206604 603076
rect 242004 603074 242604 603076
rect 278004 603074 278604 603076
rect 314004 603074 314604 603076
rect 350004 603074 350604 603076
rect 386004 603074 386604 603076
rect 422004 603074 422604 603076
rect 458004 603074 458604 603076
rect 494004 603074 494604 603076
rect 530004 603074 530604 603076
rect 566004 603074 566604 603076
rect 589920 603074 590520 603076
rect -4756 600076 -4156 600078
rect 22404 600076 23004 600078
rect 58404 600076 59004 600078
rect 94404 600076 95004 600078
rect 130404 600076 131004 600078
rect 166404 600076 167004 600078
rect 202404 600076 203004 600078
rect 238404 600076 239004 600078
rect 274404 600076 275004 600078
rect 310404 600076 311004 600078
rect 346404 600076 347004 600078
rect 382404 600076 383004 600078
rect 418404 600076 419004 600078
rect 454404 600076 455004 600078
rect 490404 600076 491004 600078
rect 526404 600076 527004 600078
rect 562404 600076 563004 600078
rect 588080 600076 588680 600078
rect -4756 600054 588680 600076
rect -4756 599818 -4574 600054
rect -4338 599818 22586 600054
rect 22822 599818 58586 600054
rect 58822 599818 94586 600054
rect 94822 599818 130586 600054
rect 130822 599818 166586 600054
rect 166822 599818 202586 600054
rect 202822 599818 238586 600054
rect 238822 599818 274586 600054
rect 274822 599818 310586 600054
rect 310822 599818 346586 600054
rect 346822 599818 382586 600054
rect 382822 599818 418586 600054
rect 418822 599818 454586 600054
rect 454822 599818 490586 600054
rect 490822 599818 526586 600054
rect 526822 599818 562586 600054
rect 562822 599818 588262 600054
rect 588498 599818 588680 600054
rect -4756 599734 588680 599818
rect -4756 599498 -4574 599734
rect -4338 599498 22586 599734
rect 22822 599498 58586 599734
rect 58822 599498 94586 599734
rect 94822 599498 130586 599734
rect 130822 599498 166586 599734
rect 166822 599498 202586 599734
rect 202822 599498 238586 599734
rect 238822 599498 274586 599734
rect 274822 599498 310586 599734
rect 310822 599498 346586 599734
rect 346822 599498 382586 599734
rect 382822 599498 418586 599734
rect 418822 599498 454586 599734
rect 454822 599498 490586 599734
rect 490822 599498 526586 599734
rect 526822 599498 562586 599734
rect 562822 599498 588262 599734
rect 588498 599498 588680 599734
rect -4756 599476 588680 599498
rect -4756 599474 -4156 599476
rect 22404 599474 23004 599476
rect 58404 599474 59004 599476
rect 94404 599474 95004 599476
rect 130404 599474 131004 599476
rect 166404 599474 167004 599476
rect 202404 599474 203004 599476
rect 238404 599474 239004 599476
rect 274404 599474 275004 599476
rect 310404 599474 311004 599476
rect 346404 599474 347004 599476
rect 382404 599474 383004 599476
rect 418404 599474 419004 599476
rect 454404 599474 455004 599476
rect 490404 599474 491004 599476
rect 526404 599474 527004 599476
rect 562404 599474 563004 599476
rect 588080 599474 588680 599476
rect -2916 596476 -2316 596478
rect 18804 596476 19404 596478
rect 54804 596476 55404 596478
rect 90804 596476 91404 596478
rect 126804 596476 127404 596478
rect 162804 596476 163404 596478
rect 198804 596476 199404 596478
rect 234804 596476 235404 596478
rect 270804 596476 271404 596478
rect 306804 596476 307404 596478
rect 342804 596476 343404 596478
rect 378804 596476 379404 596478
rect 414804 596476 415404 596478
rect 450804 596476 451404 596478
rect 486804 596476 487404 596478
rect 522804 596476 523404 596478
rect 558804 596476 559404 596478
rect 586240 596476 586840 596478
rect -2916 596454 586840 596476
rect -2916 596218 -2734 596454
rect -2498 596218 18986 596454
rect 19222 596218 54986 596454
rect 55222 596218 90986 596454
rect 91222 596218 126986 596454
rect 127222 596218 162986 596454
rect 163222 596218 198986 596454
rect 199222 596218 234986 596454
rect 235222 596218 270986 596454
rect 271222 596218 306986 596454
rect 307222 596218 342986 596454
rect 343222 596218 378986 596454
rect 379222 596218 414986 596454
rect 415222 596218 450986 596454
rect 451222 596218 486986 596454
rect 487222 596218 522986 596454
rect 523222 596218 558986 596454
rect 559222 596218 586422 596454
rect 586658 596218 586840 596454
rect -2916 596134 586840 596218
rect -2916 595898 -2734 596134
rect -2498 595898 18986 596134
rect 19222 595898 54986 596134
rect 55222 595898 90986 596134
rect 91222 595898 126986 596134
rect 127222 595898 162986 596134
rect 163222 595898 198986 596134
rect 199222 595898 234986 596134
rect 235222 595898 270986 596134
rect 271222 595898 306986 596134
rect 307222 595898 342986 596134
rect 343222 595898 378986 596134
rect 379222 595898 414986 596134
rect 415222 595898 450986 596134
rect 451222 595898 486986 596134
rect 487222 595898 522986 596134
rect 523222 595898 558986 596134
rect 559222 595898 586422 596134
rect 586658 595898 586840 596134
rect -2916 595876 586840 595898
rect -2916 595874 -2316 595876
rect 18804 595874 19404 595876
rect 54804 595874 55404 595876
rect 90804 595874 91404 595876
rect 126804 595874 127404 595876
rect 162804 595874 163404 595876
rect 198804 595874 199404 595876
rect 234804 595874 235404 595876
rect 270804 595874 271404 595876
rect 306804 595874 307404 595876
rect 342804 595874 343404 595876
rect 378804 595874 379404 595876
rect 414804 595874 415404 595876
rect 450804 595874 451404 595876
rect 486804 595874 487404 595876
rect 522804 595874 523404 595876
rect 558804 595874 559404 595876
rect 586240 595874 586840 595876
rect -7516 589276 -6916 589278
rect 11604 589276 12204 589278
rect 47604 589276 48204 589278
rect 83604 589276 84204 589278
rect 119604 589276 120204 589278
rect 155604 589276 156204 589278
rect 191604 589276 192204 589278
rect 227604 589276 228204 589278
rect 263604 589276 264204 589278
rect 299604 589276 300204 589278
rect 335604 589276 336204 589278
rect 371604 589276 372204 589278
rect 407604 589276 408204 589278
rect 443604 589276 444204 589278
rect 479604 589276 480204 589278
rect 515604 589276 516204 589278
rect 551604 589276 552204 589278
rect 590840 589276 591440 589278
rect -8436 589254 592360 589276
rect -8436 589018 -7334 589254
rect -7098 589018 11786 589254
rect 12022 589018 47786 589254
rect 48022 589018 83786 589254
rect 84022 589018 119786 589254
rect 120022 589018 155786 589254
rect 156022 589018 191786 589254
rect 192022 589018 227786 589254
rect 228022 589018 263786 589254
rect 264022 589018 299786 589254
rect 300022 589018 335786 589254
rect 336022 589018 371786 589254
rect 372022 589018 407786 589254
rect 408022 589018 443786 589254
rect 444022 589018 479786 589254
rect 480022 589018 515786 589254
rect 516022 589018 551786 589254
rect 552022 589018 591022 589254
rect 591258 589018 592360 589254
rect -8436 588934 592360 589018
rect -8436 588698 -7334 588934
rect -7098 588698 11786 588934
rect 12022 588698 47786 588934
rect 48022 588698 83786 588934
rect 84022 588698 119786 588934
rect 120022 588698 155786 588934
rect 156022 588698 191786 588934
rect 192022 588698 227786 588934
rect 228022 588698 263786 588934
rect 264022 588698 299786 588934
rect 300022 588698 335786 588934
rect 336022 588698 371786 588934
rect 372022 588698 407786 588934
rect 408022 588698 443786 588934
rect 444022 588698 479786 588934
rect 480022 588698 515786 588934
rect 516022 588698 551786 588934
rect 552022 588698 591022 588934
rect 591258 588698 592360 588934
rect -8436 588676 592360 588698
rect -7516 588674 -6916 588676
rect 11604 588674 12204 588676
rect 47604 588674 48204 588676
rect 83604 588674 84204 588676
rect 119604 588674 120204 588676
rect 155604 588674 156204 588676
rect 191604 588674 192204 588676
rect 227604 588674 228204 588676
rect 263604 588674 264204 588676
rect 299604 588674 300204 588676
rect 335604 588674 336204 588676
rect 371604 588674 372204 588676
rect 407604 588674 408204 588676
rect 443604 588674 444204 588676
rect 479604 588674 480204 588676
rect 515604 588674 516204 588676
rect 551604 588674 552204 588676
rect 590840 588674 591440 588676
rect -5676 585676 -5076 585678
rect 8004 585676 8604 585678
rect 44004 585676 44604 585678
rect 80004 585676 80604 585678
rect 116004 585676 116604 585678
rect 152004 585676 152604 585678
rect 188004 585676 188604 585678
rect 224004 585676 224604 585678
rect 260004 585676 260604 585678
rect 296004 585676 296604 585678
rect 332004 585676 332604 585678
rect 368004 585676 368604 585678
rect 404004 585676 404604 585678
rect 440004 585676 440604 585678
rect 476004 585676 476604 585678
rect 512004 585676 512604 585678
rect 548004 585676 548604 585678
rect 589000 585676 589600 585678
rect -6596 585654 590520 585676
rect -6596 585418 -5494 585654
rect -5258 585418 8186 585654
rect 8422 585418 44186 585654
rect 44422 585418 80186 585654
rect 80422 585418 116186 585654
rect 116422 585418 152186 585654
rect 152422 585418 188186 585654
rect 188422 585418 224186 585654
rect 224422 585418 260186 585654
rect 260422 585418 296186 585654
rect 296422 585418 332186 585654
rect 332422 585418 368186 585654
rect 368422 585418 404186 585654
rect 404422 585418 440186 585654
rect 440422 585418 476186 585654
rect 476422 585418 512186 585654
rect 512422 585418 548186 585654
rect 548422 585418 589182 585654
rect 589418 585418 590520 585654
rect -6596 585334 590520 585418
rect -6596 585098 -5494 585334
rect -5258 585098 8186 585334
rect 8422 585098 44186 585334
rect 44422 585098 80186 585334
rect 80422 585098 116186 585334
rect 116422 585098 152186 585334
rect 152422 585098 188186 585334
rect 188422 585098 224186 585334
rect 224422 585098 260186 585334
rect 260422 585098 296186 585334
rect 296422 585098 332186 585334
rect 332422 585098 368186 585334
rect 368422 585098 404186 585334
rect 404422 585098 440186 585334
rect 440422 585098 476186 585334
rect 476422 585098 512186 585334
rect 512422 585098 548186 585334
rect 548422 585098 589182 585334
rect 589418 585098 590520 585334
rect -6596 585076 590520 585098
rect -5676 585074 -5076 585076
rect 8004 585074 8604 585076
rect 44004 585074 44604 585076
rect 80004 585074 80604 585076
rect 116004 585074 116604 585076
rect 152004 585074 152604 585076
rect 188004 585074 188604 585076
rect 224004 585074 224604 585076
rect 260004 585074 260604 585076
rect 296004 585074 296604 585076
rect 332004 585074 332604 585076
rect 368004 585074 368604 585076
rect 404004 585074 404604 585076
rect 440004 585074 440604 585076
rect 476004 585074 476604 585076
rect 512004 585074 512604 585076
rect 548004 585074 548604 585076
rect 589000 585074 589600 585076
rect -3836 582076 -3236 582078
rect 4404 582076 5004 582078
rect 40404 582076 41004 582078
rect 76404 582076 77004 582078
rect 112404 582076 113004 582078
rect 148404 582076 149004 582078
rect 184404 582076 185004 582078
rect 220404 582076 221004 582078
rect 256404 582076 257004 582078
rect 292404 582076 293004 582078
rect 328404 582076 329004 582078
rect 364404 582076 365004 582078
rect 400404 582076 401004 582078
rect 436404 582076 437004 582078
rect 472404 582076 473004 582078
rect 508404 582076 509004 582078
rect 544404 582076 545004 582078
rect 580404 582076 581004 582078
rect 587160 582076 587760 582078
rect -4756 582054 588680 582076
rect -4756 581818 -3654 582054
rect -3418 581818 4586 582054
rect 4822 581818 40586 582054
rect 40822 581818 76586 582054
rect 76822 581818 112586 582054
rect 112822 581818 148586 582054
rect 148822 581818 184586 582054
rect 184822 581818 220586 582054
rect 220822 581818 256586 582054
rect 256822 581818 292586 582054
rect 292822 581818 328586 582054
rect 328822 581818 364586 582054
rect 364822 581818 400586 582054
rect 400822 581818 436586 582054
rect 436822 581818 472586 582054
rect 472822 581818 508586 582054
rect 508822 581818 544586 582054
rect 544822 581818 580586 582054
rect 580822 581818 587342 582054
rect 587578 581818 588680 582054
rect -4756 581734 588680 581818
rect -4756 581498 -3654 581734
rect -3418 581498 4586 581734
rect 4822 581498 40586 581734
rect 40822 581498 76586 581734
rect 76822 581498 112586 581734
rect 112822 581498 148586 581734
rect 148822 581498 184586 581734
rect 184822 581498 220586 581734
rect 220822 581498 256586 581734
rect 256822 581498 292586 581734
rect 292822 581498 328586 581734
rect 328822 581498 364586 581734
rect 364822 581498 400586 581734
rect 400822 581498 436586 581734
rect 436822 581498 472586 581734
rect 472822 581498 508586 581734
rect 508822 581498 544586 581734
rect 544822 581498 580586 581734
rect 580822 581498 587342 581734
rect 587578 581498 588680 581734
rect -4756 581476 588680 581498
rect -3836 581474 -3236 581476
rect 4404 581474 5004 581476
rect 40404 581474 41004 581476
rect 76404 581474 77004 581476
rect 112404 581474 113004 581476
rect 148404 581474 149004 581476
rect 184404 581474 185004 581476
rect 220404 581474 221004 581476
rect 256404 581474 257004 581476
rect 292404 581474 293004 581476
rect 328404 581474 329004 581476
rect 364404 581474 365004 581476
rect 400404 581474 401004 581476
rect 436404 581474 437004 581476
rect 472404 581474 473004 581476
rect 508404 581474 509004 581476
rect 544404 581474 545004 581476
rect 580404 581474 581004 581476
rect 587160 581474 587760 581476
rect -1996 578476 -1396 578478
rect 804 578476 1404 578478
rect 36804 578476 37404 578478
rect 72804 578476 73404 578478
rect 108804 578476 109404 578478
rect 144804 578476 145404 578478
rect 180804 578476 181404 578478
rect 216804 578476 217404 578478
rect 252804 578476 253404 578478
rect 288804 578476 289404 578478
rect 324804 578476 325404 578478
rect 360804 578476 361404 578478
rect 396804 578476 397404 578478
rect 432804 578476 433404 578478
rect 468804 578476 469404 578478
rect 504804 578476 505404 578478
rect 540804 578476 541404 578478
rect 576804 578476 577404 578478
rect 585320 578476 585920 578478
rect -2916 578454 586840 578476
rect -2916 578218 -1814 578454
rect -1578 578218 986 578454
rect 1222 578218 36986 578454
rect 37222 578218 72986 578454
rect 73222 578218 108986 578454
rect 109222 578218 144986 578454
rect 145222 578218 180986 578454
rect 181222 578218 216986 578454
rect 217222 578218 252986 578454
rect 253222 578218 288986 578454
rect 289222 578218 324986 578454
rect 325222 578218 360986 578454
rect 361222 578218 396986 578454
rect 397222 578218 432986 578454
rect 433222 578218 468986 578454
rect 469222 578218 504986 578454
rect 505222 578218 540986 578454
rect 541222 578218 576986 578454
rect 577222 578218 585502 578454
rect 585738 578218 586840 578454
rect -2916 578134 586840 578218
rect -2916 577898 -1814 578134
rect -1578 577898 986 578134
rect 1222 577898 36986 578134
rect 37222 577898 72986 578134
rect 73222 577898 108986 578134
rect 109222 577898 144986 578134
rect 145222 577898 180986 578134
rect 181222 577898 216986 578134
rect 217222 577898 252986 578134
rect 253222 577898 288986 578134
rect 289222 577898 324986 578134
rect 325222 577898 360986 578134
rect 361222 577898 396986 578134
rect 397222 577898 432986 578134
rect 433222 577898 468986 578134
rect 469222 577898 504986 578134
rect 505222 577898 540986 578134
rect 541222 577898 576986 578134
rect 577222 577898 585502 578134
rect 585738 577898 586840 578134
rect -2916 577876 586840 577898
rect -1996 577874 -1396 577876
rect 804 577874 1404 577876
rect 36804 577874 37404 577876
rect 72804 577874 73404 577876
rect 108804 577874 109404 577876
rect 144804 577874 145404 577876
rect 180804 577874 181404 577876
rect 216804 577874 217404 577876
rect 252804 577874 253404 577876
rect 288804 577874 289404 577876
rect 324804 577874 325404 577876
rect 360804 577874 361404 577876
rect 396804 577874 397404 577876
rect 432804 577874 433404 577876
rect 468804 577874 469404 577876
rect 504804 577874 505404 577876
rect 540804 577874 541404 577876
rect 576804 577874 577404 577876
rect 585320 577874 585920 577876
rect -8436 571276 -7836 571278
rect 29604 571276 30204 571278
rect 65604 571276 66204 571278
rect 101604 571276 102204 571278
rect 137604 571276 138204 571278
rect 173604 571276 174204 571278
rect 209604 571276 210204 571278
rect 245604 571276 246204 571278
rect 281604 571276 282204 571278
rect 317604 571276 318204 571278
rect 353604 571276 354204 571278
rect 389604 571276 390204 571278
rect 425604 571276 426204 571278
rect 461604 571276 462204 571278
rect 497604 571276 498204 571278
rect 533604 571276 534204 571278
rect 569604 571276 570204 571278
rect 591760 571276 592360 571278
rect -8436 571254 592360 571276
rect -8436 571018 -8254 571254
rect -8018 571018 29786 571254
rect 30022 571018 65786 571254
rect 66022 571018 101786 571254
rect 102022 571018 137786 571254
rect 138022 571018 173786 571254
rect 174022 571018 209786 571254
rect 210022 571018 245786 571254
rect 246022 571018 281786 571254
rect 282022 571018 317786 571254
rect 318022 571018 353786 571254
rect 354022 571018 389786 571254
rect 390022 571018 425786 571254
rect 426022 571018 461786 571254
rect 462022 571018 497786 571254
rect 498022 571018 533786 571254
rect 534022 571018 569786 571254
rect 570022 571018 591942 571254
rect 592178 571018 592360 571254
rect -8436 570934 592360 571018
rect -8436 570698 -8254 570934
rect -8018 570698 29786 570934
rect 30022 570698 65786 570934
rect 66022 570698 101786 570934
rect 102022 570698 137786 570934
rect 138022 570698 173786 570934
rect 174022 570698 209786 570934
rect 210022 570698 245786 570934
rect 246022 570698 281786 570934
rect 282022 570698 317786 570934
rect 318022 570698 353786 570934
rect 354022 570698 389786 570934
rect 390022 570698 425786 570934
rect 426022 570698 461786 570934
rect 462022 570698 497786 570934
rect 498022 570698 533786 570934
rect 534022 570698 569786 570934
rect 570022 570698 591942 570934
rect 592178 570698 592360 570934
rect -8436 570676 592360 570698
rect -8436 570674 -7836 570676
rect 29604 570674 30204 570676
rect 65604 570674 66204 570676
rect 101604 570674 102204 570676
rect 137604 570674 138204 570676
rect 173604 570674 174204 570676
rect 209604 570674 210204 570676
rect 245604 570674 246204 570676
rect 281604 570674 282204 570676
rect 317604 570674 318204 570676
rect 353604 570674 354204 570676
rect 389604 570674 390204 570676
rect 425604 570674 426204 570676
rect 461604 570674 462204 570676
rect 497604 570674 498204 570676
rect 533604 570674 534204 570676
rect 569604 570674 570204 570676
rect 591760 570674 592360 570676
rect -6596 567676 -5996 567678
rect 26004 567676 26604 567678
rect 62004 567676 62604 567678
rect 98004 567676 98604 567678
rect 134004 567676 134604 567678
rect 170004 567676 170604 567678
rect 206004 567676 206604 567678
rect 242004 567676 242604 567678
rect 278004 567676 278604 567678
rect 314004 567676 314604 567678
rect 350004 567676 350604 567678
rect 386004 567676 386604 567678
rect 422004 567676 422604 567678
rect 458004 567676 458604 567678
rect 494004 567676 494604 567678
rect 530004 567676 530604 567678
rect 566004 567676 566604 567678
rect 589920 567676 590520 567678
rect -6596 567654 590520 567676
rect -6596 567418 -6414 567654
rect -6178 567418 26186 567654
rect 26422 567418 62186 567654
rect 62422 567418 98186 567654
rect 98422 567418 134186 567654
rect 134422 567418 170186 567654
rect 170422 567418 206186 567654
rect 206422 567418 242186 567654
rect 242422 567418 278186 567654
rect 278422 567418 314186 567654
rect 314422 567418 350186 567654
rect 350422 567418 386186 567654
rect 386422 567418 422186 567654
rect 422422 567418 458186 567654
rect 458422 567418 494186 567654
rect 494422 567418 530186 567654
rect 530422 567418 566186 567654
rect 566422 567418 590102 567654
rect 590338 567418 590520 567654
rect -6596 567334 590520 567418
rect -6596 567098 -6414 567334
rect -6178 567098 26186 567334
rect 26422 567098 62186 567334
rect 62422 567098 98186 567334
rect 98422 567098 134186 567334
rect 134422 567098 170186 567334
rect 170422 567098 206186 567334
rect 206422 567098 242186 567334
rect 242422 567098 278186 567334
rect 278422 567098 314186 567334
rect 314422 567098 350186 567334
rect 350422 567098 386186 567334
rect 386422 567098 422186 567334
rect 422422 567098 458186 567334
rect 458422 567098 494186 567334
rect 494422 567098 530186 567334
rect 530422 567098 566186 567334
rect 566422 567098 590102 567334
rect 590338 567098 590520 567334
rect -6596 567076 590520 567098
rect -6596 567074 -5996 567076
rect 26004 567074 26604 567076
rect 62004 567074 62604 567076
rect 98004 567074 98604 567076
rect 134004 567074 134604 567076
rect 170004 567074 170604 567076
rect 206004 567074 206604 567076
rect 242004 567074 242604 567076
rect 278004 567074 278604 567076
rect 314004 567074 314604 567076
rect 350004 567074 350604 567076
rect 386004 567074 386604 567076
rect 422004 567074 422604 567076
rect 458004 567074 458604 567076
rect 494004 567074 494604 567076
rect 530004 567074 530604 567076
rect 566004 567074 566604 567076
rect 589920 567074 590520 567076
rect -4756 564076 -4156 564078
rect 22404 564076 23004 564078
rect 58404 564076 59004 564078
rect 94404 564076 95004 564078
rect 130404 564076 131004 564078
rect 166404 564076 167004 564078
rect 202404 564076 203004 564078
rect 238404 564076 239004 564078
rect 274404 564076 275004 564078
rect 310404 564076 311004 564078
rect 346404 564076 347004 564078
rect 382404 564076 383004 564078
rect 418404 564076 419004 564078
rect 454404 564076 455004 564078
rect 490404 564076 491004 564078
rect 526404 564076 527004 564078
rect 562404 564076 563004 564078
rect 588080 564076 588680 564078
rect -4756 564054 588680 564076
rect -4756 563818 -4574 564054
rect -4338 563818 22586 564054
rect 22822 563818 58586 564054
rect 58822 563818 94586 564054
rect 94822 563818 130586 564054
rect 130822 563818 166586 564054
rect 166822 563818 202586 564054
rect 202822 563818 238586 564054
rect 238822 563818 274586 564054
rect 274822 563818 310586 564054
rect 310822 563818 346586 564054
rect 346822 563818 382586 564054
rect 382822 563818 418586 564054
rect 418822 563818 454586 564054
rect 454822 563818 490586 564054
rect 490822 563818 526586 564054
rect 526822 563818 562586 564054
rect 562822 563818 588262 564054
rect 588498 563818 588680 564054
rect -4756 563734 588680 563818
rect -4756 563498 -4574 563734
rect -4338 563498 22586 563734
rect 22822 563498 58586 563734
rect 58822 563498 94586 563734
rect 94822 563498 130586 563734
rect 130822 563498 166586 563734
rect 166822 563498 202586 563734
rect 202822 563498 238586 563734
rect 238822 563498 274586 563734
rect 274822 563498 310586 563734
rect 310822 563498 346586 563734
rect 346822 563498 382586 563734
rect 382822 563498 418586 563734
rect 418822 563498 454586 563734
rect 454822 563498 490586 563734
rect 490822 563498 526586 563734
rect 526822 563498 562586 563734
rect 562822 563498 588262 563734
rect 588498 563498 588680 563734
rect -4756 563476 588680 563498
rect -4756 563474 -4156 563476
rect 22404 563474 23004 563476
rect 58404 563474 59004 563476
rect 94404 563474 95004 563476
rect 130404 563474 131004 563476
rect 166404 563474 167004 563476
rect 202404 563474 203004 563476
rect 238404 563474 239004 563476
rect 274404 563474 275004 563476
rect 310404 563474 311004 563476
rect 346404 563474 347004 563476
rect 382404 563474 383004 563476
rect 418404 563474 419004 563476
rect 454404 563474 455004 563476
rect 490404 563474 491004 563476
rect 526404 563474 527004 563476
rect 562404 563474 563004 563476
rect 588080 563474 588680 563476
rect 233796 562860 235404 562996
rect 5084 562818 18100 562860
rect 5084 562582 5126 562818
rect 5362 562582 18100 562818
rect 5084 562540 18100 562582
rect 17780 561500 18100 562540
rect 31028 562540 37236 562860
rect 31028 561500 31348 562540
rect 17780 561180 31348 561500
rect 36916 561500 37236 562540
rect 75556 562180 76060 562860
rect 120636 562818 125740 562860
rect 120636 562582 120678 562818
rect 120914 562582 125462 562818
rect 125698 562582 125740 562818
rect 120636 562540 125740 562582
rect 139956 562818 145060 562860
rect 139956 562582 139998 562818
rect 140234 562582 145060 562818
rect 139956 562540 145060 562582
rect 159276 562818 164380 562860
rect 159276 562582 159318 562818
rect 159554 562582 164102 562818
rect 164338 562582 164380 562818
rect 159276 562540 164380 562582
rect 167188 562818 173948 562860
rect 167188 562582 167230 562818
rect 167466 562582 173948 562818
rect 167188 562540 173948 562582
rect 178596 562818 183700 562860
rect 178596 562582 178638 562818
rect 178874 562582 183422 562818
rect 183658 562582 183700 562818
rect 178596 562540 183700 562582
rect 196628 562818 205228 562860
rect 196628 562582 196670 562818
rect 196906 562582 204950 562818
rect 205186 562582 205228 562818
rect 196628 562540 205228 562582
rect 210980 562540 220868 562860
rect 66172 561860 76060 562180
rect 66172 561500 66492 561860
rect 36916 561458 50668 561500
rect 36916 561222 50390 561458
rect 50626 561222 50668 561458
rect 36916 561180 50668 561222
rect 51452 561458 66492 561500
rect 51452 561222 51494 561458
rect 51730 561222 66492 561458
rect 51452 561180 66492 561222
rect 75740 561500 76060 561860
rect 144740 561500 145060 562540
rect 173628 561500 173948 562540
rect 210980 561500 211300 562540
rect 75740 561458 85812 561500
rect 75740 561222 85534 561458
rect 85770 561222 85812 561458
rect 75740 561180 85812 561222
rect 90092 561458 108628 561500
rect 90092 561222 90134 561458
rect 90370 561222 108350 561458
rect 108586 561222 108628 561458
rect 90092 561180 108628 561222
rect 109596 561458 117828 561500
rect 109596 561222 109638 561458
rect 109874 561222 117550 561458
rect 117786 561222 117828 561458
rect 109596 561180 117828 561222
rect 134988 561458 135860 561500
rect 134988 561222 135030 561458
rect 135266 561222 135582 561458
rect 135818 561222 135860 561458
rect 134988 561180 135860 561222
rect 144740 561458 147636 561500
rect 144740 561222 147358 561458
rect 147594 561222 147636 561458
rect 144740 561180 147636 561222
rect 154308 561458 155180 561500
rect 154308 561222 154350 561458
rect 154586 561222 154902 561458
rect 155138 561222 155180 561458
rect 154308 561180 155180 561222
rect 173628 561458 176340 561500
rect 173628 561222 176062 561458
rect 176298 561222 176340 561458
rect 173628 561180 176340 561222
rect 192948 561458 193820 561500
rect 192948 561222 192990 561458
rect 193226 561222 193542 561458
rect 193778 561222 193820 561458
rect 192948 561180 193820 561222
rect 207484 561458 211300 561500
rect 207484 561222 207526 561458
rect 207762 561222 211300 561458
rect 207484 561180 211300 561222
rect 220548 561500 220868 562540
rect 233796 562676 244420 562860
rect 233796 562180 234116 562676
rect 235084 562540 244420 562676
rect 253484 562818 263924 562860
rect 253484 562582 253526 562818
rect 253762 562582 263924 562818
rect 253484 562540 263924 562582
rect 275748 562818 285084 562860
rect 275748 562582 275790 562818
rect 276026 562582 285084 562818
rect 275748 562540 285084 562582
rect 293044 562818 299804 562860
rect 293044 562582 293086 562818
rect 293322 562582 299804 562818
rect 293044 562540 299804 562582
rect 225332 562138 234116 562180
rect 225332 561902 225374 562138
rect 225610 561902 234116 562138
rect 225332 561860 234116 561902
rect 244100 562180 244420 562540
rect 263604 562180 263924 562540
rect 284764 562180 285084 562540
rect 244100 562138 252700 562180
rect 244100 561902 252422 562138
rect 252658 561902 252700 562138
rect 244100 561860 252700 561902
rect 263604 562138 266500 562180
rect 263604 561902 266222 562138
rect 266458 561902 266500 562138
rect 263604 561860 266500 561902
rect 284764 562138 288580 562180
rect 284764 561902 288302 562138
rect 288538 561902 288580 562138
rect 284764 561860 288580 561902
rect 299484 561500 299804 562540
rect 317148 562180 317652 562860
rect 334996 562818 336972 562860
rect 334996 562582 335038 562818
rect 335274 562582 336694 562818
rect 336930 562582 336972 562818
rect 334996 562540 336972 562582
rect 349532 562818 357580 562860
rect 349532 562582 357302 562818
rect 357538 562582 357580 562818
rect 349532 562540 357580 562582
rect 370324 562818 376900 562860
rect 370324 562582 370366 562818
rect 370602 562582 376900 562818
rect 370324 562540 376900 562582
rect 349532 562180 349852 562540
rect 376580 562180 376900 562540
rect 379340 562540 386468 562860
rect 379340 562180 379660 562540
rect 307580 561860 317652 562180
rect 337204 562138 349852 562180
rect 337204 561902 337246 562138
rect 337482 561902 349852 562138
rect 337204 561860 349852 561902
rect 366828 562138 369540 562180
rect 366828 561902 366870 562138
rect 367106 561902 369262 562138
rect 369498 561902 369540 562138
rect 366828 561860 369540 561902
rect 376580 561860 379660 562180
rect 307580 561500 307900 561860
rect 220548 561458 223812 561500
rect 220548 561222 223534 561458
rect 223770 561222 223812 561458
rect 220548 561180 223812 561222
rect 299484 561180 307900 561500
rect 317332 561500 317652 561860
rect 386148 561500 386468 562540
rect 388356 562818 393460 562860
rect 388356 562582 393182 562818
rect 393418 562582 393460 562818
rect 388356 562540 393460 562582
rect 411172 562818 424556 562860
rect 411172 562582 424278 562818
rect 424514 562582 424556 562818
rect 411172 562540 424556 562582
rect 428284 562818 436332 562860
rect 428284 562582 428326 562818
rect 428562 562582 436054 562818
rect 436290 562582 436332 562818
rect 428284 562540 436332 562582
rect 388356 561500 388676 562540
rect 411172 562180 411492 562540
rect 406204 562138 411492 562180
rect 406204 561902 406246 562138
rect 406482 561902 411492 562138
rect 406204 561860 411492 561902
rect 317332 561458 318756 561500
rect 317332 561222 318478 561458
rect 318714 561222 318756 561458
rect 317332 561180 318756 561222
rect 319172 561458 325932 561500
rect 319172 561222 319214 561458
rect 319450 561222 325654 561458
rect 325890 561222 325932 561458
rect 319172 561180 325932 561222
rect 386148 561180 388676 561500
rect -2916 560476 -2316 560478
rect 18804 560476 19404 560478
rect 54804 560476 55404 560478
rect 90804 560476 91404 560478
rect 126804 560476 127404 560478
rect 162804 560476 163404 560478
rect 198804 560476 199404 560478
rect 234804 560476 235404 560478
rect 270804 560476 271404 560478
rect 306804 560476 307404 560478
rect 342804 560476 343404 560478
rect 378804 560476 379404 560478
rect 414804 560476 415404 560478
rect 450804 560476 451404 560478
rect 486804 560476 487404 560478
rect 522804 560476 523404 560478
rect 558804 560476 559404 560478
rect 586240 560476 586840 560478
rect -2916 560454 586840 560476
rect -2916 560218 -2734 560454
rect -2498 560218 18986 560454
rect 19222 560218 54986 560454
rect 55222 560218 90986 560454
rect 91222 560218 126986 560454
rect 127222 560218 162986 560454
rect 163222 560218 198986 560454
rect 199222 560218 234986 560454
rect 235222 560218 270986 560454
rect 271222 560218 306986 560454
rect 307222 560218 342986 560454
rect 343222 560218 378986 560454
rect 379222 560218 414986 560454
rect 415222 560218 450986 560454
rect 451222 560218 486986 560454
rect 487222 560218 522986 560454
rect 523222 560218 558986 560454
rect 559222 560218 586422 560454
rect 586658 560218 586840 560454
rect -2916 560134 586840 560218
rect -2916 559898 -2734 560134
rect -2498 559898 18986 560134
rect 19222 559898 54986 560134
rect 55222 559898 90986 560134
rect 91222 559898 126986 560134
rect 127222 559898 162986 560134
rect 163222 559898 198986 560134
rect 199222 559898 234986 560134
rect 235222 559898 270986 560134
rect 271222 559898 306986 560134
rect 307222 559898 342986 560134
rect 343222 559898 378986 560134
rect 379222 559898 414986 560134
rect 415222 559898 450986 560134
rect 451222 559898 486986 560134
rect 487222 559898 522986 560134
rect 523222 559898 558986 560134
rect 559222 559898 586422 560134
rect 586658 559898 586840 560134
rect -2916 559876 586840 559898
rect -2916 559874 -2316 559876
rect 18804 559874 19404 559876
rect 54804 559874 55404 559876
rect 90804 559874 91404 559876
rect 126804 559874 127404 559876
rect 162804 559874 163404 559876
rect 198804 559874 199404 559876
rect 234804 559874 235404 559876
rect 270804 559874 271404 559876
rect 306804 559874 307404 559876
rect 342804 559874 343404 559876
rect 378804 559874 379404 559876
rect 414804 559874 415404 559876
rect 450804 559874 451404 559876
rect 486804 559874 487404 559876
rect 522804 559874 523404 559876
rect 558804 559874 559404 559876
rect 586240 559874 586840 559876
rect -7516 553276 -6916 553278
rect 11604 553276 12204 553278
rect 47604 553276 48204 553278
rect 83604 553276 84204 553278
rect 119604 553276 120204 553278
rect 155604 553276 156204 553278
rect 191604 553276 192204 553278
rect 227604 553276 228204 553278
rect 263604 553276 264204 553278
rect 299604 553276 300204 553278
rect 335604 553276 336204 553278
rect 371604 553276 372204 553278
rect 407604 553276 408204 553278
rect 443604 553276 444204 553278
rect 479604 553276 480204 553278
rect 515604 553276 516204 553278
rect 551604 553276 552204 553278
rect 590840 553276 591440 553278
rect -8436 553254 592360 553276
rect -8436 553018 -7334 553254
rect -7098 553018 11786 553254
rect 12022 553018 47786 553254
rect 48022 553018 83786 553254
rect 84022 553018 119786 553254
rect 120022 553018 155786 553254
rect 156022 553018 191786 553254
rect 192022 553018 227786 553254
rect 228022 553018 263786 553254
rect 264022 553018 299786 553254
rect 300022 553018 335786 553254
rect 336022 553018 371786 553254
rect 372022 553018 407786 553254
rect 408022 553018 443786 553254
rect 444022 553018 479786 553254
rect 480022 553018 515786 553254
rect 516022 553018 551786 553254
rect 552022 553018 591022 553254
rect 591258 553018 592360 553254
rect -8436 552934 592360 553018
rect -8436 552698 -7334 552934
rect -7098 552698 11786 552934
rect 12022 552698 47786 552934
rect 48022 552698 83786 552934
rect 84022 552698 119786 552934
rect 120022 552698 155786 552934
rect 156022 552698 191786 552934
rect 192022 552698 227786 552934
rect 228022 552698 263786 552934
rect 264022 552698 299786 552934
rect 300022 552698 335786 552934
rect 336022 552698 371786 552934
rect 372022 552698 407786 552934
rect 408022 552698 443786 552934
rect 444022 552698 479786 552934
rect 480022 552698 515786 552934
rect 516022 552698 551786 552934
rect 552022 552698 591022 552934
rect 591258 552698 592360 552934
rect -8436 552676 592360 552698
rect -7516 552674 -6916 552676
rect 11604 552674 12204 552676
rect 47604 552674 48204 552676
rect 83604 552674 84204 552676
rect 119604 552674 120204 552676
rect 155604 552674 156204 552676
rect 191604 552674 192204 552676
rect 227604 552674 228204 552676
rect 263604 552674 264204 552676
rect 299604 552674 300204 552676
rect 335604 552674 336204 552676
rect 371604 552674 372204 552676
rect 407604 552674 408204 552676
rect 443604 552674 444204 552676
rect 479604 552674 480204 552676
rect 515604 552674 516204 552676
rect 551604 552674 552204 552676
rect 590840 552674 591440 552676
rect -5676 549676 -5076 549678
rect 8004 549676 8604 549678
rect 44004 549676 44604 549678
rect 80004 549676 80604 549678
rect 116004 549676 116604 549678
rect 152004 549676 152604 549678
rect 188004 549676 188604 549678
rect 224004 549676 224604 549678
rect 260004 549676 260604 549678
rect 296004 549676 296604 549678
rect 332004 549676 332604 549678
rect 368004 549676 368604 549678
rect 404004 549676 404604 549678
rect 440004 549676 440604 549678
rect 476004 549676 476604 549678
rect 512004 549676 512604 549678
rect 548004 549676 548604 549678
rect 589000 549676 589600 549678
rect -6596 549654 590520 549676
rect -6596 549418 -5494 549654
rect -5258 549418 8186 549654
rect 8422 549418 44186 549654
rect 44422 549418 80186 549654
rect 80422 549418 116186 549654
rect 116422 549418 152186 549654
rect 152422 549418 188186 549654
rect 188422 549418 224186 549654
rect 224422 549418 260186 549654
rect 260422 549418 296186 549654
rect 296422 549418 332186 549654
rect 332422 549418 368186 549654
rect 368422 549418 404186 549654
rect 404422 549418 440186 549654
rect 440422 549418 476186 549654
rect 476422 549418 512186 549654
rect 512422 549418 548186 549654
rect 548422 549418 589182 549654
rect 589418 549418 590520 549654
rect -6596 549334 590520 549418
rect -6596 549098 -5494 549334
rect -5258 549098 8186 549334
rect 8422 549098 44186 549334
rect 44422 549098 80186 549334
rect 80422 549098 116186 549334
rect 116422 549098 152186 549334
rect 152422 549098 188186 549334
rect 188422 549098 224186 549334
rect 224422 549098 260186 549334
rect 260422 549098 296186 549334
rect 296422 549098 332186 549334
rect 332422 549098 368186 549334
rect 368422 549098 404186 549334
rect 404422 549098 440186 549334
rect 440422 549098 476186 549334
rect 476422 549098 512186 549334
rect 512422 549098 548186 549334
rect 548422 549098 589182 549334
rect 589418 549098 590520 549334
rect -6596 549076 590520 549098
rect -5676 549074 -5076 549076
rect 8004 549074 8604 549076
rect 44004 549074 44604 549076
rect 80004 549074 80604 549076
rect 116004 549074 116604 549076
rect 152004 549074 152604 549076
rect 188004 549074 188604 549076
rect 224004 549074 224604 549076
rect 260004 549074 260604 549076
rect 296004 549074 296604 549076
rect 332004 549074 332604 549076
rect 368004 549074 368604 549076
rect 404004 549074 404604 549076
rect 440004 549074 440604 549076
rect 476004 549074 476604 549076
rect 512004 549074 512604 549076
rect 548004 549074 548604 549076
rect 589000 549074 589600 549076
rect -3836 546076 -3236 546078
rect 4404 546076 5004 546078
rect 40404 546076 41004 546078
rect 76404 546076 77004 546078
rect 112404 546076 113004 546078
rect 148404 546076 149004 546078
rect 184404 546076 185004 546078
rect 220404 546076 221004 546078
rect 256404 546076 257004 546078
rect 292404 546076 293004 546078
rect 328404 546076 329004 546078
rect 364404 546076 365004 546078
rect 400404 546076 401004 546078
rect 436404 546076 437004 546078
rect 472404 546076 473004 546078
rect 508404 546076 509004 546078
rect 544404 546076 545004 546078
rect 580404 546076 581004 546078
rect 587160 546076 587760 546078
rect -4756 546054 588680 546076
rect -4756 545818 -3654 546054
rect -3418 545818 4586 546054
rect 4822 545818 40586 546054
rect 40822 545818 76586 546054
rect 76822 545818 112586 546054
rect 112822 545818 148586 546054
rect 148822 545818 184586 546054
rect 184822 545818 220586 546054
rect 220822 545818 256586 546054
rect 256822 545818 292586 546054
rect 292822 545818 328586 546054
rect 328822 545818 364586 546054
rect 364822 545818 400586 546054
rect 400822 545818 436586 546054
rect 436822 545818 472586 546054
rect 472822 545818 508586 546054
rect 508822 545818 544586 546054
rect 544822 545818 580586 546054
rect 580822 545818 587342 546054
rect 587578 545818 588680 546054
rect -4756 545734 588680 545818
rect -4756 545498 -3654 545734
rect -3418 545498 4586 545734
rect 4822 545498 40586 545734
rect 40822 545498 76586 545734
rect 76822 545498 112586 545734
rect 112822 545498 148586 545734
rect 148822 545498 184586 545734
rect 184822 545498 220586 545734
rect 220822 545498 256586 545734
rect 256822 545498 292586 545734
rect 292822 545498 328586 545734
rect 328822 545498 364586 545734
rect 364822 545498 400586 545734
rect 400822 545498 436586 545734
rect 436822 545498 472586 545734
rect 472822 545498 508586 545734
rect 508822 545498 544586 545734
rect 544822 545498 580586 545734
rect 580822 545498 587342 545734
rect 587578 545498 588680 545734
rect -4756 545476 588680 545498
rect -3836 545474 -3236 545476
rect 4404 545474 5004 545476
rect 40404 545474 41004 545476
rect 76404 545474 77004 545476
rect 112404 545474 113004 545476
rect 148404 545474 149004 545476
rect 184404 545474 185004 545476
rect 220404 545474 221004 545476
rect 256404 545474 257004 545476
rect 292404 545474 293004 545476
rect 328404 545474 329004 545476
rect 364404 545474 365004 545476
rect 400404 545474 401004 545476
rect 436404 545474 437004 545476
rect 472404 545474 473004 545476
rect 508404 545474 509004 545476
rect 544404 545474 545004 545476
rect 580404 545474 581004 545476
rect 587160 545474 587760 545476
rect -1996 542476 -1396 542478
rect 804 542476 1404 542478
rect 36804 542476 37404 542478
rect 72804 542476 73404 542478
rect 108804 542476 109404 542478
rect 144804 542476 145404 542478
rect 180804 542476 181404 542478
rect 216804 542476 217404 542478
rect 252804 542476 253404 542478
rect 288804 542476 289404 542478
rect 324804 542476 325404 542478
rect 360804 542476 361404 542478
rect 396804 542476 397404 542478
rect 432804 542476 433404 542478
rect 468804 542476 469404 542478
rect 504804 542476 505404 542478
rect 540804 542476 541404 542478
rect 576804 542476 577404 542478
rect 585320 542476 585920 542478
rect -2916 542454 586840 542476
rect -2916 542218 -1814 542454
rect -1578 542218 986 542454
rect 1222 542218 36986 542454
rect 37222 542218 72986 542454
rect 73222 542218 108986 542454
rect 109222 542218 144986 542454
rect 145222 542218 180986 542454
rect 181222 542218 216986 542454
rect 217222 542218 252986 542454
rect 253222 542218 288986 542454
rect 289222 542218 324986 542454
rect 325222 542218 360986 542454
rect 361222 542218 396986 542454
rect 397222 542218 432986 542454
rect 433222 542218 468986 542454
rect 469222 542218 504986 542454
rect 505222 542218 540986 542454
rect 541222 542218 576986 542454
rect 577222 542218 585502 542454
rect 585738 542218 586840 542454
rect -2916 542134 586840 542218
rect -2916 541898 -1814 542134
rect -1578 541898 986 542134
rect 1222 541898 36986 542134
rect 37222 541898 72986 542134
rect 73222 541898 108986 542134
rect 109222 541898 144986 542134
rect 145222 541898 180986 542134
rect 181222 541898 216986 542134
rect 217222 541898 252986 542134
rect 253222 541898 288986 542134
rect 289222 541898 324986 542134
rect 325222 541898 360986 542134
rect 361222 541898 396986 542134
rect 397222 541898 432986 542134
rect 433222 541898 468986 542134
rect 469222 541898 504986 542134
rect 505222 541898 540986 542134
rect 541222 541898 576986 542134
rect 577222 541898 585502 542134
rect 585738 541898 586840 542134
rect -2916 541876 586840 541898
rect -1996 541874 -1396 541876
rect 804 541874 1404 541876
rect 36804 541874 37404 541876
rect 72804 541874 73404 541876
rect 108804 541874 109404 541876
rect 144804 541874 145404 541876
rect 180804 541874 181404 541876
rect 216804 541874 217404 541876
rect 252804 541874 253404 541876
rect 288804 541874 289404 541876
rect 324804 541874 325404 541876
rect 360804 541874 361404 541876
rect 396804 541874 397404 541876
rect 432804 541874 433404 541876
rect 468804 541874 469404 541876
rect 504804 541874 505404 541876
rect 540804 541874 541404 541876
rect 576804 541874 577404 541876
rect 585320 541874 585920 541876
rect -8436 535276 -7836 535278
rect 29604 535276 30204 535278
rect 65604 535276 66204 535278
rect 101604 535276 102204 535278
rect 137604 535276 138204 535278
rect 173604 535276 174204 535278
rect 209604 535276 210204 535278
rect 245604 535276 246204 535278
rect 281604 535276 282204 535278
rect 317604 535276 318204 535278
rect 353604 535276 354204 535278
rect 389604 535276 390204 535278
rect 425604 535276 426204 535278
rect 461604 535276 462204 535278
rect 497604 535276 498204 535278
rect 533604 535276 534204 535278
rect 569604 535276 570204 535278
rect 591760 535276 592360 535278
rect -8436 535254 592360 535276
rect -8436 535018 -8254 535254
rect -8018 535018 29786 535254
rect 30022 535018 65786 535254
rect 66022 535018 101786 535254
rect 102022 535018 137786 535254
rect 138022 535018 173786 535254
rect 174022 535018 209786 535254
rect 210022 535018 245786 535254
rect 246022 535018 281786 535254
rect 282022 535018 317786 535254
rect 318022 535018 353786 535254
rect 354022 535018 389786 535254
rect 390022 535018 425786 535254
rect 426022 535018 461786 535254
rect 462022 535018 497786 535254
rect 498022 535018 533786 535254
rect 534022 535018 569786 535254
rect 570022 535018 591942 535254
rect 592178 535018 592360 535254
rect -8436 534934 592360 535018
rect -8436 534698 -8254 534934
rect -8018 534698 29786 534934
rect 30022 534698 65786 534934
rect 66022 534698 101786 534934
rect 102022 534698 137786 534934
rect 138022 534698 173786 534934
rect 174022 534698 209786 534934
rect 210022 534698 245786 534934
rect 246022 534698 281786 534934
rect 282022 534698 317786 534934
rect 318022 534698 353786 534934
rect 354022 534698 389786 534934
rect 390022 534698 425786 534934
rect 426022 534698 461786 534934
rect 462022 534698 497786 534934
rect 498022 534698 533786 534934
rect 534022 534698 569786 534934
rect 570022 534698 591942 534934
rect 592178 534698 592360 534934
rect -8436 534676 592360 534698
rect -8436 534674 -7836 534676
rect 29604 534674 30204 534676
rect 65604 534674 66204 534676
rect 101604 534674 102204 534676
rect 137604 534674 138204 534676
rect 173604 534674 174204 534676
rect 209604 534674 210204 534676
rect 245604 534674 246204 534676
rect 281604 534674 282204 534676
rect 317604 534674 318204 534676
rect 353604 534674 354204 534676
rect 389604 534674 390204 534676
rect 425604 534674 426204 534676
rect 461604 534674 462204 534676
rect 497604 534674 498204 534676
rect 533604 534674 534204 534676
rect 569604 534674 570204 534676
rect 591760 534674 592360 534676
rect -6596 531676 -5996 531678
rect 26004 531676 26604 531678
rect 62004 531676 62604 531678
rect 98004 531676 98604 531678
rect 134004 531676 134604 531678
rect 170004 531676 170604 531678
rect 206004 531676 206604 531678
rect 242004 531676 242604 531678
rect 278004 531676 278604 531678
rect 314004 531676 314604 531678
rect 350004 531676 350604 531678
rect 386004 531676 386604 531678
rect 422004 531676 422604 531678
rect 458004 531676 458604 531678
rect 494004 531676 494604 531678
rect 530004 531676 530604 531678
rect 566004 531676 566604 531678
rect 589920 531676 590520 531678
rect -6596 531654 590520 531676
rect -6596 531418 -6414 531654
rect -6178 531418 26186 531654
rect 26422 531418 62186 531654
rect 62422 531418 98186 531654
rect 98422 531418 134186 531654
rect 134422 531418 170186 531654
rect 170422 531418 206186 531654
rect 206422 531418 242186 531654
rect 242422 531418 278186 531654
rect 278422 531418 314186 531654
rect 314422 531418 350186 531654
rect 350422 531418 386186 531654
rect 386422 531418 422186 531654
rect 422422 531418 458186 531654
rect 458422 531418 494186 531654
rect 494422 531418 530186 531654
rect 530422 531418 566186 531654
rect 566422 531418 590102 531654
rect 590338 531418 590520 531654
rect -6596 531334 590520 531418
rect -6596 531098 -6414 531334
rect -6178 531098 26186 531334
rect 26422 531098 62186 531334
rect 62422 531098 98186 531334
rect 98422 531098 134186 531334
rect 134422 531098 170186 531334
rect 170422 531098 206186 531334
rect 206422 531098 242186 531334
rect 242422 531098 278186 531334
rect 278422 531098 314186 531334
rect 314422 531098 350186 531334
rect 350422 531098 386186 531334
rect 386422 531098 422186 531334
rect 422422 531098 458186 531334
rect 458422 531098 494186 531334
rect 494422 531098 530186 531334
rect 530422 531098 566186 531334
rect 566422 531098 590102 531334
rect 590338 531098 590520 531334
rect -6596 531076 590520 531098
rect -6596 531074 -5996 531076
rect 26004 531074 26604 531076
rect 62004 531074 62604 531076
rect 98004 531074 98604 531076
rect 134004 531074 134604 531076
rect 170004 531074 170604 531076
rect 206004 531074 206604 531076
rect 242004 531074 242604 531076
rect 278004 531074 278604 531076
rect 314004 531074 314604 531076
rect 350004 531074 350604 531076
rect 386004 531074 386604 531076
rect 422004 531074 422604 531076
rect 458004 531074 458604 531076
rect 494004 531074 494604 531076
rect 530004 531074 530604 531076
rect 566004 531074 566604 531076
rect 589920 531074 590520 531076
rect -4756 528076 -4156 528078
rect 22404 528076 23004 528078
rect 58404 528076 59004 528078
rect 94404 528076 95004 528078
rect 130404 528076 131004 528078
rect 166404 528076 167004 528078
rect 202404 528076 203004 528078
rect 238404 528076 239004 528078
rect 274404 528076 275004 528078
rect 310404 528076 311004 528078
rect 346404 528076 347004 528078
rect 382404 528076 383004 528078
rect 418404 528076 419004 528078
rect 454404 528076 455004 528078
rect 490404 528076 491004 528078
rect 526404 528076 527004 528078
rect 562404 528076 563004 528078
rect 588080 528076 588680 528078
rect -4756 528054 588680 528076
rect -4756 527818 -4574 528054
rect -4338 527818 22586 528054
rect 22822 527818 58586 528054
rect 58822 527818 94586 528054
rect 94822 527818 130586 528054
rect 130822 527818 166586 528054
rect 166822 527818 202586 528054
rect 202822 527818 238586 528054
rect 238822 527818 274586 528054
rect 274822 527818 310586 528054
rect 310822 527818 346586 528054
rect 346822 527818 382586 528054
rect 382822 527818 418586 528054
rect 418822 527818 454586 528054
rect 454822 527818 490586 528054
rect 490822 527818 526586 528054
rect 526822 527818 562586 528054
rect 562822 527818 588262 528054
rect 588498 527818 588680 528054
rect -4756 527734 588680 527818
rect -4756 527498 -4574 527734
rect -4338 527498 22586 527734
rect 22822 527498 58586 527734
rect 58822 527498 94586 527734
rect 94822 527498 130586 527734
rect 130822 527498 166586 527734
rect 166822 527498 202586 527734
rect 202822 527498 238586 527734
rect 238822 527498 274586 527734
rect 274822 527498 310586 527734
rect 310822 527498 346586 527734
rect 346822 527498 382586 527734
rect 382822 527498 418586 527734
rect 418822 527498 454586 527734
rect 454822 527498 490586 527734
rect 490822 527498 526586 527734
rect 526822 527498 562586 527734
rect 562822 527498 588262 527734
rect 588498 527498 588680 527734
rect -4756 527476 588680 527498
rect -4756 527474 -4156 527476
rect 22404 527474 23004 527476
rect 58404 527474 59004 527476
rect 94404 527474 95004 527476
rect 130404 527474 131004 527476
rect 166404 527474 167004 527476
rect 202404 527474 203004 527476
rect 238404 527474 239004 527476
rect 274404 527474 275004 527476
rect 310404 527474 311004 527476
rect 346404 527474 347004 527476
rect 382404 527474 383004 527476
rect 418404 527474 419004 527476
rect 454404 527474 455004 527476
rect 490404 527474 491004 527476
rect 526404 527474 527004 527476
rect 562404 527474 563004 527476
rect 588080 527474 588680 527476
rect -2916 524476 -2316 524478
rect 18804 524476 19404 524478
rect 54804 524476 55404 524478
rect 90804 524476 91404 524478
rect 126804 524476 127404 524478
rect 162804 524476 163404 524478
rect 198804 524476 199404 524478
rect 234804 524476 235404 524478
rect 270804 524476 271404 524478
rect 306804 524476 307404 524478
rect 342804 524476 343404 524478
rect 378804 524476 379404 524478
rect 414804 524476 415404 524478
rect 450804 524476 451404 524478
rect 486804 524476 487404 524478
rect 522804 524476 523404 524478
rect 558804 524476 559404 524478
rect 586240 524476 586840 524478
rect -2916 524454 586840 524476
rect -2916 524218 -2734 524454
rect -2498 524218 18986 524454
rect 19222 524218 54986 524454
rect 55222 524218 90986 524454
rect 91222 524218 126986 524454
rect 127222 524218 162986 524454
rect 163222 524218 198986 524454
rect 199222 524218 234986 524454
rect 235222 524218 270986 524454
rect 271222 524218 306986 524454
rect 307222 524218 342986 524454
rect 343222 524218 378986 524454
rect 379222 524218 414986 524454
rect 415222 524218 450986 524454
rect 451222 524218 486986 524454
rect 487222 524218 522986 524454
rect 523222 524218 558986 524454
rect 559222 524218 586422 524454
rect 586658 524218 586840 524454
rect -2916 524134 586840 524218
rect -2916 523898 -2734 524134
rect -2498 523898 18986 524134
rect 19222 523898 54986 524134
rect 55222 523898 90986 524134
rect 91222 523898 126986 524134
rect 127222 523898 162986 524134
rect 163222 523898 198986 524134
rect 199222 523898 234986 524134
rect 235222 523898 270986 524134
rect 271222 523898 306986 524134
rect 307222 523898 342986 524134
rect 343222 523898 378986 524134
rect 379222 523898 414986 524134
rect 415222 523898 450986 524134
rect 451222 523898 486986 524134
rect 487222 523898 522986 524134
rect 523222 523898 558986 524134
rect 559222 523898 586422 524134
rect 586658 523898 586840 524134
rect -2916 523876 586840 523898
rect -2916 523874 -2316 523876
rect 18804 523874 19404 523876
rect 54804 523874 55404 523876
rect 90804 523874 91404 523876
rect 126804 523874 127404 523876
rect 162804 523874 163404 523876
rect 198804 523874 199404 523876
rect 234804 523874 235404 523876
rect 270804 523874 271404 523876
rect 306804 523874 307404 523876
rect 342804 523874 343404 523876
rect 378804 523874 379404 523876
rect 414804 523874 415404 523876
rect 450804 523874 451404 523876
rect 486804 523874 487404 523876
rect 522804 523874 523404 523876
rect 558804 523874 559404 523876
rect 586240 523874 586840 523876
rect -7516 517276 -6916 517278
rect 11604 517276 12204 517278
rect 47604 517276 48204 517278
rect 83604 517276 84204 517278
rect 119604 517276 120204 517278
rect 155604 517276 156204 517278
rect 191604 517276 192204 517278
rect 227604 517276 228204 517278
rect 263604 517276 264204 517278
rect 299604 517276 300204 517278
rect 335604 517276 336204 517278
rect 371604 517276 372204 517278
rect 407604 517276 408204 517278
rect 443604 517276 444204 517278
rect 479604 517276 480204 517278
rect 515604 517276 516204 517278
rect 551604 517276 552204 517278
rect 590840 517276 591440 517278
rect -8436 517254 592360 517276
rect -8436 517018 -7334 517254
rect -7098 517018 11786 517254
rect 12022 517018 47786 517254
rect 48022 517018 83786 517254
rect 84022 517018 119786 517254
rect 120022 517018 155786 517254
rect 156022 517018 191786 517254
rect 192022 517018 227786 517254
rect 228022 517018 263786 517254
rect 264022 517018 299786 517254
rect 300022 517018 335786 517254
rect 336022 517018 371786 517254
rect 372022 517018 407786 517254
rect 408022 517018 443786 517254
rect 444022 517018 479786 517254
rect 480022 517018 515786 517254
rect 516022 517018 551786 517254
rect 552022 517018 591022 517254
rect 591258 517018 592360 517254
rect -8436 516934 592360 517018
rect -8436 516698 -7334 516934
rect -7098 516698 11786 516934
rect 12022 516698 47786 516934
rect 48022 516698 83786 516934
rect 84022 516698 119786 516934
rect 120022 516698 155786 516934
rect 156022 516698 191786 516934
rect 192022 516698 227786 516934
rect 228022 516698 263786 516934
rect 264022 516698 299786 516934
rect 300022 516698 335786 516934
rect 336022 516698 371786 516934
rect 372022 516698 407786 516934
rect 408022 516698 443786 516934
rect 444022 516698 479786 516934
rect 480022 516698 515786 516934
rect 516022 516698 551786 516934
rect 552022 516698 591022 516934
rect 591258 516698 592360 516934
rect -8436 516676 592360 516698
rect -7516 516674 -6916 516676
rect 11604 516674 12204 516676
rect 47604 516674 48204 516676
rect 83604 516674 84204 516676
rect 119604 516674 120204 516676
rect 155604 516674 156204 516676
rect 191604 516674 192204 516676
rect 227604 516674 228204 516676
rect 263604 516674 264204 516676
rect 299604 516674 300204 516676
rect 335604 516674 336204 516676
rect 371604 516674 372204 516676
rect 407604 516674 408204 516676
rect 443604 516674 444204 516676
rect 479604 516674 480204 516676
rect 515604 516674 516204 516676
rect 551604 516674 552204 516676
rect 590840 516674 591440 516676
rect -5676 513676 -5076 513678
rect 8004 513676 8604 513678
rect 44004 513676 44604 513678
rect 80004 513676 80604 513678
rect 116004 513676 116604 513678
rect 152004 513676 152604 513678
rect 188004 513676 188604 513678
rect 224004 513676 224604 513678
rect 260004 513676 260604 513678
rect 296004 513676 296604 513678
rect 332004 513676 332604 513678
rect 368004 513676 368604 513678
rect 404004 513676 404604 513678
rect 440004 513676 440604 513678
rect 476004 513676 476604 513678
rect 512004 513676 512604 513678
rect 548004 513676 548604 513678
rect 589000 513676 589600 513678
rect -6596 513654 590520 513676
rect -6596 513418 -5494 513654
rect -5258 513418 8186 513654
rect 8422 513418 44186 513654
rect 44422 513418 80186 513654
rect 80422 513418 116186 513654
rect 116422 513418 152186 513654
rect 152422 513418 188186 513654
rect 188422 513418 224186 513654
rect 224422 513418 260186 513654
rect 260422 513418 296186 513654
rect 296422 513418 332186 513654
rect 332422 513418 368186 513654
rect 368422 513418 404186 513654
rect 404422 513418 440186 513654
rect 440422 513418 476186 513654
rect 476422 513418 512186 513654
rect 512422 513418 548186 513654
rect 548422 513418 589182 513654
rect 589418 513418 590520 513654
rect -6596 513334 590520 513418
rect -6596 513098 -5494 513334
rect -5258 513098 8186 513334
rect 8422 513098 44186 513334
rect 44422 513098 80186 513334
rect 80422 513098 116186 513334
rect 116422 513098 152186 513334
rect 152422 513098 188186 513334
rect 188422 513098 224186 513334
rect 224422 513098 260186 513334
rect 260422 513098 296186 513334
rect 296422 513098 332186 513334
rect 332422 513098 368186 513334
rect 368422 513098 404186 513334
rect 404422 513098 440186 513334
rect 440422 513098 476186 513334
rect 476422 513098 512186 513334
rect 512422 513098 548186 513334
rect 548422 513098 589182 513334
rect 589418 513098 590520 513334
rect -6596 513076 590520 513098
rect -5676 513074 -5076 513076
rect 8004 513074 8604 513076
rect 44004 513074 44604 513076
rect 80004 513074 80604 513076
rect 116004 513074 116604 513076
rect 152004 513074 152604 513076
rect 188004 513074 188604 513076
rect 224004 513074 224604 513076
rect 260004 513074 260604 513076
rect 296004 513074 296604 513076
rect 332004 513074 332604 513076
rect 368004 513074 368604 513076
rect 404004 513074 404604 513076
rect 440004 513074 440604 513076
rect 476004 513074 476604 513076
rect 512004 513074 512604 513076
rect 548004 513074 548604 513076
rect 589000 513074 589600 513076
rect -3836 510076 -3236 510078
rect 4404 510076 5004 510078
rect 40404 510076 41004 510078
rect 76404 510076 77004 510078
rect 112404 510076 113004 510078
rect 148404 510076 149004 510078
rect 184404 510076 185004 510078
rect 220404 510076 221004 510078
rect 256404 510076 257004 510078
rect 292404 510076 293004 510078
rect 328404 510076 329004 510078
rect 364404 510076 365004 510078
rect 400404 510076 401004 510078
rect 436404 510076 437004 510078
rect 472404 510076 473004 510078
rect 508404 510076 509004 510078
rect 544404 510076 545004 510078
rect 580404 510076 581004 510078
rect 587160 510076 587760 510078
rect -4756 510054 588680 510076
rect -4756 509818 -3654 510054
rect -3418 509818 4586 510054
rect 4822 509818 40586 510054
rect 40822 509818 76586 510054
rect 76822 509818 112586 510054
rect 112822 509818 148586 510054
rect 148822 509818 184586 510054
rect 184822 509818 220586 510054
rect 220822 509818 256586 510054
rect 256822 509818 292586 510054
rect 292822 509818 328586 510054
rect 328822 509818 364586 510054
rect 364822 509818 400586 510054
rect 400822 509818 436586 510054
rect 436822 509818 472586 510054
rect 472822 509818 508586 510054
rect 508822 509818 544586 510054
rect 544822 509818 580586 510054
rect 580822 509818 587342 510054
rect 587578 509818 588680 510054
rect -4756 509734 588680 509818
rect -4756 509498 -3654 509734
rect -3418 509498 4586 509734
rect 4822 509498 40586 509734
rect 40822 509498 76586 509734
rect 76822 509498 112586 509734
rect 112822 509498 148586 509734
rect 148822 509498 184586 509734
rect 184822 509498 220586 509734
rect 220822 509498 256586 509734
rect 256822 509498 292586 509734
rect 292822 509498 328586 509734
rect 328822 509498 364586 509734
rect 364822 509498 400586 509734
rect 400822 509498 436586 509734
rect 436822 509498 472586 509734
rect 472822 509498 508586 509734
rect 508822 509498 544586 509734
rect 544822 509498 580586 509734
rect 580822 509498 587342 509734
rect 587578 509498 588680 509734
rect -4756 509476 588680 509498
rect -3836 509474 -3236 509476
rect 4404 509474 5004 509476
rect 40404 509474 41004 509476
rect 76404 509474 77004 509476
rect 112404 509474 113004 509476
rect 148404 509474 149004 509476
rect 184404 509474 185004 509476
rect 220404 509474 221004 509476
rect 256404 509474 257004 509476
rect 292404 509474 293004 509476
rect 328404 509474 329004 509476
rect 364404 509474 365004 509476
rect 400404 509474 401004 509476
rect 436404 509474 437004 509476
rect 472404 509474 473004 509476
rect 508404 509474 509004 509476
rect 544404 509474 545004 509476
rect 580404 509474 581004 509476
rect 587160 509474 587760 509476
rect -1996 506476 -1396 506478
rect 804 506476 1404 506478
rect 36804 506476 37404 506478
rect 72804 506476 73404 506478
rect 108804 506476 109404 506478
rect 144804 506476 145404 506478
rect 180804 506476 181404 506478
rect 216804 506476 217404 506478
rect 252804 506476 253404 506478
rect 288804 506476 289404 506478
rect 324804 506476 325404 506478
rect 360804 506476 361404 506478
rect 396804 506476 397404 506478
rect 432804 506476 433404 506478
rect 468804 506476 469404 506478
rect 504804 506476 505404 506478
rect 540804 506476 541404 506478
rect 576804 506476 577404 506478
rect 585320 506476 585920 506478
rect -2916 506454 586840 506476
rect -2916 506218 -1814 506454
rect -1578 506218 986 506454
rect 1222 506218 36986 506454
rect 37222 506218 72986 506454
rect 73222 506218 108986 506454
rect 109222 506218 144986 506454
rect 145222 506218 180986 506454
rect 181222 506218 216986 506454
rect 217222 506218 252986 506454
rect 253222 506218 288986 506454
rect 289222 506218 324986 506454
rect 325222 506218 360986 506454
rect 361222 506218 396986 506454
rect 397222 506218 432986 506454
rect 433222 506218 468986 506454
rect 469222 506218 504986 506454
rect 505222 506218 540986 506454
rect 541222 506218 576986 506454
rect 577222 506218 585502 506454
rect 585738 506218 586840 506454
rect -2916 506134 586840 506218
rect -2916 505898 -1814 506134
rect -1578 505898 986 506134
rect 1222 505898 36986 506134
rect 37222 505898 72986 506134
rect 73222 505898 108986 506134
rect 109222 505898 144986 506134
rect 145222 505898 180986 506134
rect 181222 505898 216986 506134
rect 217222 505898 252986 506134
rect 253222 505898 288986 506134
rect 289222 505898 324986 506134
rect 325222 505898 360986 506134
rect 361222 505898 396986 506134
rect 397222 505898 432986 506134
rect 433222 505898 468986 506134
rect 469222 505898 504986 506134
rect 505222 505898 540986 506134
rect 541222 505898 576986 506134
rect 577222 505898 585502 506134
rect 585738 505898 586840 506134
rect -2916 505876 586840 505898
rect -1996 505874 -1396 505876
rect 804 505874 1404 505876
rect 36804 505874 37404 505876
rect 72804 505874 73404 505876
rect 108804 505874 109404 505876
rect 144804 505874 145404 505876
rect 180804 505874 181404 505876
rect 216804 505874 217404 505876
rect 252804 505874 253404 505876
rect 288804 505874 289404 505876
rect 324804 505874 325404 505876
rect 360804 505874 361404 505876
rect 396804 505874 397404 505876
rect 432804 505874 433404 505876
rect 468804 505874 469404 505876
rect 504804 505874 505404 505876
rect 540804 505874 541404 505876
rect 576804 505874 577404 505876
rect 585320 505874 585920 505876
rect -8436 499276 -7836 499278
rect 29604 499276 30204 499278
rect 65604 499276 66204 499278
rect 101604 499276 102204 499278
rect 137604 499276 138204 499278
rect 173604 499276 174204 499278
rect 209604 499276 210204 499278
rect 245604 499276 246204 499278
rect 281604 499276 282204 499278
rect 317604 499276 318204 499278
rect 353604 499276 354204 499278
rect 389604 499276 390204 499278
rect 425604 499276 426204 499278
rect 461604 499276 462204 499278
rect 497604 499276 498204 499278
rect 533604 499276 534204 499278
rect 569604 499276 570204 499278
rect 591760 499276 592360 499278
rect -8436 499254 592360 499276
rect -8436 499018 -8254 499254
rect -8018 499018 29786 499254
rect 30022 499018 65786 499254
rect 66022 499018 101786 499254
rect 102022 499018 137786 499254
rect 138022 499018 173786 499254
rect 174022 499018 209786 499254
rect 210022 499018 245786 499254
rect 246022 499018 281786 499254
rect 282022 499018 317786 499254
rect 318022 499018 353786 499254
rect 354022 499018 389786 499254
rect 390022 499018 425786 499254
rect 426022 499018 461786 499254
rect 462022 499018 497786 499254
rect 498022 499018 533786 499254
rect 534022 499018 569786 499254
rect 570022 499018 591942 499254
rect 592178 499018 592360 499254
rect -8436 498934 592360 499018
rect -8436 498698 -8254 498934
rect -8018 498698 29786 498934
rect 30022 498698 65786 498934
rect 66022 498698 101786 498934
rect 102022 498698 137786 498934
rect 138022 498698 173786 498934
rect 174022 498698 209786 498934
rect 210022 498698 245786 498934
rect 246022 498698 281786 498934
rect 282022 498698 317786 498934
rect 318022 498698 353786 498934
rect 354022 498698 389786 498934
rect 390022 498698 425786 498934
rect 426022 498698 461786 498934
rect 462022 498698 497786 498934
rect 498022 498698 533786 498934
rect 534022 498698 569786 498934
rect 570022 498698 591942 498934
rect 592178 498698 592360 498934
rect -8436 498676 592360 498698
rect -8436 498674 -7836 498676
rect 29604 498674 30204 498676
rect 65604 498674 66204 498676
rect 101604 498674 102204 498676
rect 137604 498674 138204 498676
rect 173604 498674 174204 498676
rect 209604 498674 210204 498676
rect 245604 498674 246204 498676
rect 281604 498674 282204 498676
rect 317604 498674 318204 498676
rect 353604 498674 354204 498676
rect 389604 498674 390204 498676
rect 425604 498674 426204 498676
rect 461604 498674 462204 498676
rect 497604 498674 498204 498676
rect 533604 498674 534204 498676
rect 569604 498674 570204 498676
rect 591760 498674 592360 498676
rect -6596 495676 -5996 495678
rect 26004 495676 26604 495678
rect 62004 495676 62604 495678
rect 98004 495676 98604 495678
rect 134004 495676 134604 495678
rect 170004 495676 170604 495678
rect 206004 495676 206604 495678
rect 242004 495676 242604 495678
rect 278004 495676 278604 495678
rect 314004 495676 314604 495678
rect 350004 495676 350604 495678
rect 386004 495676 386604 495678
rect 422004 495676 422604 495678
rect 458004 495676 458604 495678
rect 494004 495676 494604 495678
rect 530004 495676 530604 495678
rect 566004 495676 566604 495678
rect 589920 495676 590520 495678
rect -6596 495654 590520 495676
rect -6596 495418 -6414 495654
rect -6178 495418 26186 495654
rect 26422 495418 62186 495654
rect 62422 495418 98186 495654
rect 98422 495418 134186 495654
rect 134422 495418 170186 495654
rect 170422 495418 206186 495654
rect 206422 495418 242186 495654
rect 242422 495418 278186 495654
rect 278422 495418 314186 495654
rect 314422 495418 350186 495654
rect 350422 495418 386186 495654
rect 386422 495418 422186 495654
rect 422422 495418 458186 495654
rect 458422 495418 494186 495654
rect 494422 495418 530186 495654
rect 530422 495418 566186 495654
rect 566422 495418 590102 495654
rect 590338 495418 590520 495654
rect -6596 495334 590520 495418
rect -6596 495098 -6414 495334
rect -6178 495098 26186 495334
rect 26422 495098 62186 495334
rect 62422 495098 98186 495334
rect 98422 495098 134186 495334
rect 134422 495098 170186 495334
rect 170422 495098 206186 495334
rect 206422 495098 242186 495334
rect 242422 495098 278186 495334
rect 278422 495098 314186 495334
rect 314422 495098 350186 495334
rect 350422 495098 386186 495334
rect 386422 495098 422186 495334
rect 422422 495098 458186 495334
rect 458422 495098 494186 495334
rect 494422 495098 530186 495334
rect 530422 495098 566186 495334
rect 566422 495098 590102 495334
rect 590338 495098 590520 495334
rect -6596 495076 590520 495098
rect -6596 495074 -5996 495076
rect 26004 495074 26604 495076
rect 62004 495074 62604 495076
rect 98004 495074 98604 495076
rect 134004 495074 134604 495076
rect 170004 495074 170604 495076
rect 206004 495074 206604 495076
rect 242004 495074 242604 495076
rect 278004 495074 278604 495076
rect 314004 495074 314604 495076
rect 350004 495074 350604 495076
rect 386004 495074 386604 495076
rect 422004 495074 422604 495076
rect 458004 495074 458604 495076
rect 494004 495074 494604 495076
rect 530004 495074 530604 495076
rect 566004 495074 566604 495076
rect 589920 495074 590520 495076
rect -4756 492076 -4156 492078
rect 22404 492076 23004 492078
rect 58404 492076 59004 492078
rect 94404 492076 95004 492078
rect 130404 492076 131004 492078
rect 166404 492076 167004 492078
rect 202404 492076 203004 492078
rect 238404 492076 239004 492078
rect 274404 492076 275004 492078
rect 310404 492076 311004 492078
rect 346404 492076 347004 492078
rect 382404 492076 383004 492078
rect 418404 492076 419004 492078
rect 454404 492076 455004 492078
rect 490404 492076 491004 492078
rect 526404 492076 527004 492078
rect 562404 492076 563004 492078
rect 588080 492076 588680 492078
rect -4756 492054 588680 492076
rect -4756 491818 -4574 492054
rect -4338 491818 22586 492054
rect 22822 491818 58586 492054
rect 58822 491818 94586 492054
rect 94822 491818 130586 492054
rect 130822 491818 166586 492054
rect 166822 491818 202586 492054
rect 202822 491818 238586 492054
rect 238822 491818 274586 492054
rect 274822 491818 310586 492054
rect 310822 491818 346586 492054
rect 346822 491818 382586 492054
rect 382822 491818 418586 492054
rect 418822 491818 454586 492054
rect 454822 491818 490586 492054
rect 490822 491818 526586 492054
rect 526822 491818 562586 492054
rect 562822 491818 588262 492054
rect 588498 491818 588680 492054
rect -4756 491734 588680 491818
rect -4756 491498 -4574 491734
rect -4338 491498 22586 491734
rect 22822 491498 58586 491734
rect 58822 491498 94586 491734
rect 94822 491498 130586 491734
rect 130822 491498 166586 491734
rect 166822 491498 202586 491734
rect 202822 491498 238586 491734
rect 238822 491498 274586 491734
rect 274822 491498 310586 491734
rect 310822 491498 346586 491734
rect 346822 491498 382586 491734
rect 382822 491498 418586 491734
rect 418822 491498 454586 491734
rect 454822 491498 490586 491734
rect 490822 491498 526586 491734
rect 526822 491498 562586 491734
rect 562822 491498 588262 491734
rect 588498 491498 588680 491734
rect -4756 491476 588680 491498
rect -4756 491474 -4156 491476
rect 22404 491474 23004 491476
rect 58404 491474 59004 491476
rect 94404 491474 95004 491476
rect 130404 491474 131004 491476
rect 166404 491474 167004 491476
rect 202404 491474 203004 491476
rect 238404 491474 239004 491476
rect 274404 491474 275004 491476
rect 310404 491474 311004 491476
rect 346404 491474 347004 491476
rect 382404 491474 383004 491476
rect 418404 491474 419004 491476
rect 454404 491474 455004 491476
rect 490404 491474 491004 491476
rect 526404 491474 527004 491476
rect 562404 491474 563004 491476
rect 588080 491474 588680 491476
rect -2916 488476 -2316 488478
rect 18804 488476 19404 488478
rect 54804 488476 55404 488478
rect 90804 488476 91404 488478
rect 126804 488476 127404 488478
rect 162804 488476 163404 488478
rect 198804 488476 199404 488478
rect 234804 488476 235404 488478
rect 270804 488476 271404 488478
rect 306804 488476 307404 488478
rect 342804 488476 343404 488478
rect 378804 488476 379404 488478
rect 414804 488476 415404 488478
rect 450804 488476 451404 488478
rect 486804 488476 487404 488478
rect 522804 488476 523404 488478
rect 558804 488476 559404 488478
rect 586240 488476 586840 488478
rect -2916 488454 586840 488476
rect -2916 488218 -2734 488454
rect -2498 488218 18986 488454
rect 19222 488218 54986 488454
rect 55222 488218 90986 488454
rect 91222 488218 126986 488454
rect 127222 488218 162986 488454
rect 163222 488218 198986 488454
rect 199222 488218 234986 488454
rect 235222 488218 270986 488454
rect 271222 488218 306986 488454
rect 307222 488218 342986 488454
rect 343222 488218 378986 488454
rect 379222 488218 414986 488454
rect 415222 488218 450986 488454
rect 451222 488218 486986 488454
rect 487222 488218 522986 488454
rect 523222 488218 558986 488454
rect 559222 488218 586422 488454
rect 586658 488218 586840 488454
rect -2916 488134 586840 488218
rect -2916 487898 -2734 488134
rect -2498 487898 18986 488134
rect 19222 487898 54986 488134
rect 55222 487898 90986 488134
rect 91222 487898 126986 488134
rect 127222 487898 162986 488134
rect 163222 487898 198986 488134
rect 199222 487898 234986 488134
rect 235222 487898 270986 488134
rect 271222 487898 306986 488134
rect 307222 487898 342986 488134
rect 343222 487898 378986 488134
rect 379222 487898 414986 488134
rect 415222 487898 450986 488134
rect 451222 487898 486986 488134
rect 487222 487898 522986 488134
rect 523222 487898 558986 488134
rect 559222 487898 586422 488134
rect 586658 487898 586840 488134
rect -2916 487876 586840 487898
rect -2916 487874 -2316 487876
rect 18804 487874 19404 487876
rect 54804 487874 55404 487876
rect 90804 487874 91404 487876
rect 126804 487874 127404 487876
rect 162804 487874 163404 487876
rect 198804 487874 199404 487876
rect 234804 487874 235404 487876
rect 270804 487874 271404 487876
rect 306804 487874 307404 487876
rect 342804 487874 343404 487876
rect 378804 487874 379404 487876
rect 414804 487874 415404 487876
rect 450804 487874 451404 487876
rect 486804 487874 487404 487876
rect 522804 487874 523404 487876
rect 558804 487874 559404 487876
rect 586240 487874 586840 487876
rect -7516 481276 -6916 481278
rect 11604 481276 12204 481278
rect 47604 481276 48204 481278
rect 83604 481276 84204 481278
rect 119604 481276 120204 481278
rect 155604 481276 156204 481278
rect 191604 481276 192204 481278
rect 227604 481276 228204 481278
rect 263604 481276 264204 481278
rect 299604 481276 300204 481278
rect 335604 481276 336204 481278
rect 371604 481276 372204 481278
rect 407604 481276 408204 481278
rect 443604 481276 444204 481278
rect 479604 481276 480204 481278
rect 515604 481276 516204 481278
rect 551604 481276 552204 481278
rect 590840 481276 591440 481278
rect -8436 481254 592360 481276
rect -8436 481018 -7334 481254
rect -7098 481018 11786 481254
rect 12022 481018 47786 481254
rect 48022 481018 83786 481254
rect 84022 481018 119786 481254
rect 120022 481018 155786 481254
rect 156022 481018 191786 481254
rect 192022 481018 227786 481254
rect 228022 481018 263786 481254
rect 264022 481018 299786 481254
rect 300022 481018 335786 481254
rect 336022 481018 371786 481254
rect 372022 481018 407786 481254
rect 408022 481018 443786 481254
rect 444022 481018 479786 481254
rect 480022 481018 515786 481254
rect 516022 481018 551786 481254
rect 552022 481018 591022 481254
rect 591258 481018 592360 481254
rect -8436 480934 592360 481018
rect -8436 480698 -7334 480934
rect -7098 480698 11786 480934
rect 12022 480698 47786 480934
rect 48022 480698 83786 480934
rect 84022 480698 119786 480934
rect 120022 480698 155786 480934
rect 156022 480698 191786 480934
rect 192022 480698 227786 480934
rect 228022 480698 263786 480934
rect 264022 480698 299786 480934
rect 300022 480698 335786 480934
rect 336022 480698 371786 480934
rect 372022 480698 407786 480934
rect 408022 480698 443786 480934
rect 444022 480698 479786 480934
rect 480022 480698 515786 480934
rect 516022 480698 551786 480934
rect 552022 480698 591022 480934
rect 591258 480698 592360 480934
rect -8436 480676 592360 480698
rect -7516 480674 -6916 480676
rect 11604 480674 12204 480676
rect 47604 480674 48204 480676
rect 83604 480674 84204 480676
rect 119604 480674 120204 480676
rect 155604 480674 156204 480676
rect 191604 480674 192204 480676
rect 227604 480674 228204 480676
rect 263604 480674 264204 480676
rect 299604 480674 300204 480676
rect 335604 480674 336204 480676
rect 371604 480674 372204 480676
rect 407604 480674 408204 480676
rect 443604 480674 444204 480676
rect 479604 480674 480204 480676
rect 515604 480674 516204 480676
rect 551604 480674 552204 480676
rect 590840 480674 591440 480676
rect -5676 477676 -5076 477678
rect 8004 477676 8604 477678
rect 44004 477676 44604 477678
rect 80004 477676 80604 477678
rect 116004 477676 116604 477678
rect 152004 477676 152604 477678
rect 188004 477676 188604 477678
rect 224004 477676 224604 477678
rect 260004 477676 260604 477678
rect 296004 477676 296604 477678
rect 332004 477676 332604 477678
rect 368004 477676 368604 477678
rect 404004 477676 404604 477678
rect 440004 477676 440604 477678
rect 476004 477676 476604 477678
rect 512004 477676 512604 477678
rect 548004 477676 548604 477678
rect 589000 477676 589600 477678
rect -6596 477654 590520 477676
rect -6596 477418 -5494 477654
rect -5258 477418 8186 477654
rect 8422 477418 44186 477654
rect 44422 477418 80186 477654
rect 80422 477418 116186 477654
rect 116422 477418 152186 477654
rect 152422 477418 188186 477654
rect 188422 477418 224186 477654
rect 224422 477418 260186 477654
rect 260422 477418 296186 477654
rect 296422 477418 332186 477654
rect 332422 477418 368186 477654
rect 368422 477418 404186 477654
rect 404422 477418 440186 477654
rect 440422 477418 476186 477654
rect 476422 477418 512186 477654
rect 512422 477418 548186 477654
rect 548422 477418 589182 477654
rect 589418 477418 590520 477654
rect -6596 477334 590520 477418
rect -6596 477098 -5494 477334
rect -5258 477098 8186 477334
rect 8422 477098 44186 477334
rect 44422 477098 80186 477334
rect 80422 477098 116186 477334
rect 116422 477098 152186 477334
rect 152422 477098 188186 477334
rect 188422 477098 224186 477334
rect 224422 477098 260186 477334
rect 260422 477098 296186 477334
rect 296422 477098 332186 477334
rect 332422 477098 368186 477334
rect 368422 477098 404186 477334
rect 404422 477098 440186 477334
rect 440422 477098 476186 477334
rect 476422 477098 512186 477334
rect 512422 477098 548186 477334
rect 548422 477098 589182 477334
rect 589418 477098 590520 477334
rect -6596 477076 590520 477098
rect -5676 477074 -5076 477076
rect 8004 477074 8604 477076
rect 44004 477074 44604 477076
rect 80004 477074 80604 477076
rect 116004 477074 116604 477076
rect 152004 477074 152604 477076
rect 188004 477074 188604 477076
rect 224004 477074 224604 477076
rect 260004 477074 260604 477076
rect 296004 477074 296604 477076
rect 332004 477074 332604 477076
rect 368004 477074 368604 477076
rect 404004 477074 404604 477076
rect 440004 477074 440604 477076
rect 476004 477074 476604 477076
rect 512004 477074 512604 477076
rect 548004 477074 548604 477076
rect 589000 477074 589600 477076
rect -3836 474076 -3236 474078
rect 4404 474076 5004 474078
rect 40404 474076 41004 474078
rect 76404 474076 77004 474078
rect 112404 474076 113004 474078
rect 148404 474076 149004 474078
rect 184404 474076 185004 474078
rect 220404 474076 221004 474078
rect 256404 474076 257004 474078
rect 292404 474076 293004 474078
rect 328404 474076 329004 474078
rect 364404 474076 365004 474078
rect 400404 474076 401004 474078
rect 436404 474076 437004 474078
rect 472404 474076 473004 474078
rect 508404 474076 509004 474078
rect 544404 474076 545004 474078
rect 580404 474076 581004 474078
rect 587160 474076 587760 474078
rect -4756 474054 588680 474076
rect -4756 473818 -3654 474054
rect -3418 473818 4586 474054
rect 4822 473818 40586 474054
rect 40822 473818 76586 474054
rect 76822 473818 112586 474054
rect 112822 473818 148586 474054
rect 148822 473818 184586 474054
rect 184822 473818 220586 474054
rect 220822 473818 256586 474054
rect 256822 473818 292586 474054
rect 292822 473818 328586 474054
rect 328822 473818 364586 474054
rect 364822 473818 400586 474054
rect 400822 473818 436586 474054
rect 436822 473818 472586 474054
rect 472822 473818 508586 474054
rect 508822 473818 544586 474054
rect 544822 473818 580586 474054
rect 580822 473818 587342 474054
rect 587578 473818 588680 474054
rect -4756 473734 588680 473818
rect -4756 473498 -3654 473734
rect -3418 473498 4586 473734
rect 4822 473498 40586 473734
rect 40822 473498 76586 473734
rect 76822 473498 112586 473734
rect 112822 473498 148586 473734
rect 148822 473498 184586 473734
rect 184822 473498 220586 473734
rect 220822 473498 256586 473734
rect 256822 473498 292586 473734
rect 292822 473498 328586 473734
rect 328822 473498 364586 473734
rect 364822 473498 400586 473734
rect 400822 473498 436586 473734
rect 436822 473498 472586 473734
rect 472822 473498 508586 473734
rect 508822 473498 544586 473734
rect 544822 473498 580586 473734
rect 580822 473498 587342 473734
rect 587578 473498 588680 473734
rect -4756 473476 588680 473498
rect -3836 473474 -3236 473476
rect 4404 473474 5004 473476
rect 40404 473474 41004 473476
rect 76404 473474 77004 473476
rect 112404 473474 113004 473476
rect 148404 473474 149004 473476
rect 184404 473474 185004 473476
rect 220404 473474 221004 473476
rect 256404 473474 257004 473476
rect 292404 473474 293004 473476
rect 328404 473474 329004 473476
rect 364404 473474 365004 473476
rect 400404 473474 401004 473476
rect 436404 473474 437004 473476
rect 472404 473474 473004 473476
rect 508404 473474 509004 473476
rect 544404 473474 545004 473476
rect 580404 473474 581004 473476
rect 587160 473474 587760 473476
rect -1996 470476 -1396 470478
rect 804 470476 1404 470478
rect 36804 470476 37404 470478
rect 72804 470476 73404 470478
rect 108804 470476 109404 470478
rect 144804 470476 145404 470478
rect 180804 470476 181404 470478
rect 216804 470476 217404 470478
rect 252804 470476 253404 470478
rect 288804 470476 289404 470478
rect 324804 470476 325404 470478
rect 360804 470476 361404 470478
rect 396804 470476 397404 470478
rect 432804 470476 433404 470478
rect 468804 470476 469404 470478
rect 504804 470476 505404 470478
rect 540804 470476 541404 470478
rect 576804 470476 577404 470478
rect 585320 470476 585920 470478
rect -2916 470454 586840 470476
rect -2916 470218 -1814 470454
rect -1578 470218 986 470454
rect 1222 470218 36986 470454
rect 37222 470218 72986 470454
rect 73222 470218 108986 470454
rect 109222 470218 144986 470454
rect 145222 470218 180986 470454
rect 181222 470218 216986 470454
rect 217222 470218 252986 470454
rect 253222 470218 288986 470454
rect 289222 470218 324986 470454
rect 325222 470218 360986 470454
rect 361222 470218 396986 470454
rect 397222 470218 432986 470454
rect 433222 470218 468986 470454
rect 469222 470218 504986 470454
rect 505222 470218 540986 470454
rect 541222 470218 576986 470454
rect 577222 470218 585502 470454
rect 585738 470218 586840 470454
rect -2916 470134 586840 470218
rect -2916 469898 -1814 470134
rect -1578 469898 986 470134
rect 1222 469898 36986 470134
rect 37222 469898 72986 470134
rect 73222 469898 108986 470134
rect 109222 469898 144986 470134
rect 145222 469898 180986 470134
rect 181222 469898 216986 470134
rect 217222 469898 252986 470134
rect 253222 469898 288986 470134
rect 289222 469898 324986 470134
rect 325222 469898 360986 470134
rect 361222 469898 396986 470134
rect 397222 469898 432986 470134
rect 433222 469898 468986 470134
rect 469222 469898 504986 470134
rect 505222 469898 540986 470134
rect 541222 469898 576986 470134
rect 577222 469898 585502 470134
rect 585738 469898 586840 470134
rect -2916 469876 586840 469898
rect -1996 469874 -1396 469876
rect 804 469874 1404 469876
rect 36804 469874 37404 469876
rect 72804 469874 73404 469876
rect 108804 469874 109404 469876
rect 144804 469874 145404 469876
rect 180804 469874 181404 469876
rect 216804 469874 217404 469876
rect 252804 469874 253404 469876
rect 288804 469874 289404 469876
rect 324804 469874 325404 469876
rect 360804 469874 361404 469876
rect 396804 469874 397404 469876
rect 432804 469874 433404 469876
rect 468804 469874 469404 469876
rect 504804 469874 505404 469876
rect 540804 469874 541404 469876
rect 576804 469874 577404 469876
rect 585320 469874 585920 469876
rect -8436 463276 -7836 463278
rect 29604 463276 30204 463278
rect 65604 463276 66204 463278
rect 101604 463276 102204 463278
rect 137604 463276 138204 463278
rect 173604 463276 174204 463278
rect 209604 463276 210204 463278
rect 245604 463276 246204 463278
rect 281604 463276 282204 463278
rect 317604 463276 318204 463278
rect 353604 463276 354204 463278
rect 389604 463276 390204 463278
rect 425604 463276 426204 463278
rect 461604 463276 462204 463278
rect 497604 463276 498204 463278
rect 533604 463276 534204 463278
rect 569604 463276 570204 463278
rect 591760 463276 592360 463278
rect -8436 463254 592360 463276
rect -8436 463018 -8254 463254
rect -8018 463018 29786 463254
rect 30022 463018 65786 463254
rect 66022 463018 101786 463254
rect 102022 463018 137786 463254
rect 138022 463018 173786 463254
rect 174022 463018 209786 463254
rect 210022 463018 245786 463254
rect 246022 463018 281786 463254
rect 282022 463018 317786 463254
rect 318022 463018 353786 463254
rect 354022 463018 389786 463254
rect 390022 463018 425786 463254
rect 426022 463018 461786 463254
rect 462022 463018 497786 463254
rect 498022 463018 533786 463254
rect 534022 463018 569786 463254
rect 570022 463018 591942 463254
rect 592178 463018 592360 463254
rect -8436 462934 592360 463018
rect -8436 462698 -8254 462934
rect -8018 462698 29786 462934
rect 30022 462698 65786 462934
rect 66022 462698 101786 462934
rect 102022 462698 137786 462934
rect 138022 462698 173786 462934
rect 174022 462698 209786 462934
rect 210022 462698 245786 462934
rect 246022 462698 281786 462934
rect 282022 462698 317786 462934
rect 318022 462698 353786 462934
rect 354022 462698 389786 462934
rect 390022 462698 425786 462934
rect 426022 462698 461786 462934
rect 462022 462698 497786 462934
rect 498022 462698 533786 462934
rect 534022 462698 569786 462934
rect 570022 462698 591942 462934
rect 592178 462698 592360 462934
rect -8436 462676 592360 462698
rect -8436 462674 -7836 462676
rect 29604 462674 30204 462676
rect 65604 462674 66204 462676
rect 101604 462674 102204 462676
rect 137604 462674 138204 462676
rect 173604 462674 174204 462676
rect 209604 462674 210204 462676
rect 245604 462674 246204 462676
rect 281604 462674 282204 462676
rect 317604 462674 318204 462676
rect 353604 462674 354204 462676
rect 389604 462674 390204 462676
rect 425604 462674 426204 462676
rect 461604 462674 462204 462676
rect 497604 462674 498204 462676
rect 533604 462674 534204 462676
rect 569604 462674 570204 462676
rect 591760 462674 592360 462676
rect -6596 459676 -5996 459678
rect 26004 459676 26604 459678
rect 62004 459676 62604 459678
rect 98004 459676 98604 459678
rect 134004 459676 134604 459678
rect 170004 459676 170604 459678
rect 206004 459676 206604 459678
rect 242004 459676 242604 459678
rect 278004 459676 278604 459678
rect 314004 459676 314604 459678
rect 350004 459676 350604 459678
rect 386004 459676 386604 459678
rect 422004 459676 422604 459678
rect 458004 459676 458604 459678
rect 494004 459676 494604 459678
rect 530004 459676 530604 459678
rect 566004 459676 566604 459678
rect 589920 459676 590520 459678
rect -6596 459654 590520 459676
rect -6596 459418 -6414 459654
rect -6178 459418 26186 459654
rect 26422 459418 62186 459654
rect 62422 459418 98186 459654
rect 98422 459418 134186 459654
rect 134422 459418 170186 459654
rect 170422 459418 206186 459654
rect 206422 459418 242186 459654
rect 242422 459418 278186 459654
rect 278422 459418 314186 459654
rect 314422 459418 350186 459654
rect 350422 459418 386186 459654
rect 386422 459418 422186 459654
rect 422422 459418 458186 459654
rect 458422 459418 494186 459654
rect 494422 459418 530186 459654
rect 530422 459418 566186 459654
rect 566422 459418 590102 459654
rect 590338 459418 590520 459654
rect -6596 459334 590520 459418
rect -6596 459098 -6414 459334
rect -6178 459098 26186 459334
rect 26422 459098 62186 459334
rect 62422 459098 98186 459334
rect 98422 459098 134186 459334
rect 134422 459098 170186 459334
rect 170422 459098 206186 459334
rect 206422 459098 242186 459334
rect 242422 459098 278186 459334
rect 278422 459098 314186 459334
rect 314422 459098 350186 459334
rect 350422 459098 386186 459334
rect 386422 459098 422186 459334
rect 422422 459098 458186 459334
rect 458422 459098 494186 459334
rect 494422 459098 530186 459334
rect 530422 459098 566186 459334
rect 566422 459098 590102 459334
rect 590338 459098 590520 459334
rect -6596 459076 590520 459098
rect -6596 459074 -5996 459076
rect 26004 459074 26604 459076
rect 62004 459074 62604 459076
rect 98004 459074 98604 459076
rect 134004 459074 134604 459076
rect 170004 459074 170604 459076
rect 206004 459074 206604 459076
rect 242004 459074 242604 459076
rect 278004 459074 278604 459076
rect 314004 459074 314604 459076
rect 350004 459074 350604 459076
rect 386004 459074 386604 459076
rect 422004 459074 422604 459076
rect 458004 459074 458604 459076
rect 494004 459074 494604 459076
rect 530004 459074 530604 459076
rect 566004 459074 566604 459076
rect 589920 459074 590520 459076
rect -4756 456076 -4156 456078
rect 22404 456076 23004 456078
rect 58404 456076 59004 456078
rect 94404 456076 95004 456078
rect 130404 456076 131004 456078
rect 166404 456076 167004 456078
rect 202404 456076 203004 456078
rect 238404 456076 239004 456078
rect 274404 456076 275004 456078
rect 310404 456076 311004 456078
rect 346404 456076 347004 456078
rect 382404 456076 383004 456078
rect 418404 456076 419004 456078
rect 454404 456076 455004 456078
rect 490404 456076 491004 456078
rect 526404 456076 527004 456078
rect 562404 456076 563004 456078
rect 588080 456076 588680 456078
rect -4756 456054 588680 456076
rect -4756 455818 -4574 456054
rect -4338 455818 22586 456054
rect 22822 455818 58586 456054
rect 58822 455818 94586 456054
rect 94822 455818 130586 456054
rect 130822 455818 166586 456054
rect 166822 455818 202586 456054
rect 202822 455818 238586 456054
rect 238822 455818 274586 456054
rect 274822 455818 310586 456054
rect 310822 455818 346586 456054
rect 346822 455818 382586 456054
rect 382822 455818 418586 456054
rect 418822 455818 454586 456054
rect 454822 455818 490586 456054
rect 490822 455818 526586 456054
rect 526822 455818 562586 456054
rect 562822 455818 588262 456054
rect 588498 455818 588680 456054
rect -4756 455734 588680 455818
rect -4756 455498 -4574 455734
rect -4338 455498 22586 455734
rect 22822 455498 58586 455734
rect 58822 455498 94586 455734
rect 94822 455498 130586 455734
rect 130822 455498 166586 455734
rect 166822 455498 202586 455734
rect 202822 455498 238586 455734
rect 238822 455498 274586 455734
rect 274822 455498 310586 455734
rect 310822 455498 346586 455734
rect 346822 455498 382586 455734
rect 382822 455498 418586 455734
rect 418822 455498 454586 455734
rect 454822 455498 490586 455734
rect 490822 455498 526586 455734
rect 526822 455498 562586 455734
rect 562822 455498 588262 455734
rect 588498 455498 588680 455734
rect -4756 455476 588680 455498
rect -4756 455474 -4156 455476
rect 22404 455474 23004 455476
rect 58404 455474 59004 455476
rect 94404 455474 95004 455476
rect 130404 455474 131004 455476
rect 166404 455474 167004 455476
rect 202404 455474 203004 455476
rect 238404 455474 239004 455476
rect 274404 455474 275004 455476
rect 310404 455474 311004 455476
rect 346404 455474 347004 455476
rect 382404 455474 383004 455476
rect 418404 455474 419004 455476
rect 454404 455474 455004 455476
rect 490404 455474 491004 455476
rect 526404 455474 527004 455476
rect 562404 455474 563004 455476
rect 588080 455474 588680 455476
rect -2916 452476 -2316 452478
rect 18804 452476 19404 452478
rect 54804 452476 55404 452478
rect 90804 452476 91404 452478
rect 126804 452476 127404 452478
rect 162804 452476 163404 452478
rect 198804 452476 199404 452478
rect 234804 452476 235404 452478
rect 270804 452476 271404 452478
rect 306804 452476 307404 452478
rect 342804 452476 343404 452478
rect 378804 452476 379404 452478
rect 414804 452476 415404 452478
rect 450804 452476 451404 452478
rect 486804 452476 487404 452478
rect 522804 452476 523404 452478
rect 558804 452476 559404 452478
rect 586240 452476 586840 452478
rect -2916 452454 586840 452476
rect -2916 452218 -2734 452454
rect -2498 452218 18986 452454
rect 19222 452218 54986 452454
rect 55222 452218 90986 452454
rect 91222 452218 126986 452454
rect 127222 452218 162986 452454
rect 163222 452218 198986 452454
rect 199222 452218 234986 452454
rect 235222 452218 270986 452454
rect 271222 452218 306986 452454
rect 307222 452218 342986 452454
rect 343222 452218 378986 452454
rect 379222 452218 414986 452454
rect 415222 452218 450986 452454
rect 451222 452218 486986 452454
rect 487222 452218 522986 452454
rect 523222 452218 558986 452454
rect 559222 452218 586422 452454
rect 586658 452218 586840 452454
rect -2916 452134 586840 452218
rect -2916 451898 -2734 452134
rect -2498 451898 18986 452134
rect 19222 451898 54986 452134
rect 55222 451898 90986 452134
rect 91222 451898 126986 452134
rect 127222 451898 162986 452134
rect 163222 451898 198986 452134
rect 199222 451898 234986 452134
rect 235222 451898 270986 452134
rect 271222 451898 306986 452134
rect 307222 451898 342986 452134
rect 343222 451898 378986 452134
rect 379222 451898 414986 452134
rect 415222 451898 450986 452134
rect 451222 451898 486986 452134
rect 487222 451898 522986 452134
rect 523222 451898 558986 452134
rect 559222 451898 586422 452134
rect 586658 451898 586840 452134
rect -2916 451876 586840 451898
rect -2916 451874 -2316 451876
rect 18804 451874 19404 451876
rect 54804 451874 55404 451876
rect 90804 451874 91404 451876
rect 126804 451874 127404 451876
rect 162804 451874 163404 451876
rect 198804 451874 199404 451876
rect 234804 451874 235404 451876
rect 270804 451874 271404 451876
rect 306804 451874 307404 451876
rect 342804 451874 343404 451876
rect 378804 451874 379404 451876
rect 414804 451874 415404 451876
rect 450804 451874 451404 451876
rect 486804 451874 487404 451876
rect 522804 451874 523404 451876
rect 558804 451874 559404 451876
rect 586240 451874 586840 451876
rect -7516 445276 -6916 445278
rect 11604 445276 12204 445278
rect 47604 445276 48204 445278
rect 83604 445276 84204 445278
rect 119604 445276 120204 445278
rect 155604 445276 156204 445278
rect 191604 445276 192204 445278
rect 227604 445276 228204 445278
rect 263604 445276 264204 445278
rect 299604 445276 300204 445278
rect 335604 445276 336204 445278
rect 371604 445276 372204 445278
rect 407604 445276 408204 445278
rect 443604 445276 444204 445278
rect 479604 445276 480204 445278
rect 515604 445276 516204 445278
rect 551604 445276 552204 445278
rect 590840 445276 591440 445278
rect -8436 445254 592360 445276
rect -8436 445018 -7334 445254
rect -7098 445018 11786 445254
rect 12022 445018 47786 445254
rect 48022 445018 83786 445254
rect 84022 445018 119786 445254
rect 120022 445018 155786 445254
rect 156022 445018 191786 445254
rect 192022 445018 227786 445254
rect 228022 445018 263786 445254
rect 264022 445018 299786 445254
rect 300022 445018 335786 445254
rect 336022 445018 371786 445254
rect 372022 445018 407786 445254
rect 408022 445018 443786 445254
rect 444022 445018 479786 445254
rect 480022 445018 515786 445254
rect 516022 445018 551786 445254
rect 552022 445018 591022 445254
rect 591258 445018 592360 445254
rect -8436 444934 592360 445018
rect -8436 444698 -7334 444934
rect -7098 444698 11786 444934
rect 12022 444698 47786 444934
rect 48022 444698 83786 444934
rect 84022 444698 119786 444934
rect 120022 444698 155786 444934
rect 156022 444698 191786 444934
rect 192022 444698 227786 444934
rect 228022 444698 263786 444934
rect 264022 444698 299786 444934
rect 300022 444698 335786 444934
rect 336022 444698 371786 444934
rect 372022 444698 407786 444934
rect 408022 444698 443786 444934
rect 444022 444698 479786 444934
rect 480022 444698 515786 444934
rect 516022 444698 551786 444934
rect 552022 444698 591022 444934
rect 591258 444698 592360 444934
rect -8436 444676 592360 444698
rect -7516 444674 -6916 444676
rect 11604 444674 12204 444676
rect 47604 444674 48204 444676
rect 83604 444674 84204 444676
rect 119604 444674 120204 444676
rect 155604 444674 156204 444676
rect 191604 444674 192204 444676
rect 227604 444674 228204 444676
rect 263604 444674 264204 444676
rect 299604 444674 300204 444676
rect 335604 444674 336204 444676
rect 371604 444674 372204 444676
rect 407604 444674 408204 444676
rect 443604 444674 444204 444676
rect 479604 444674 480204 444676
rect 515604 444674 516204 444676
rect 551604 444674 552204 444676
rect 590840 444674 591440 444676
rect -5676 441676 -5076 441678
rect 8004 441676 8604 441678
rect 44004 441676 44604 441678
rect 80004 441676 80604 441678
rect 116004 441676 116604 441678
rect 152004 441676 152604 441678
rect 188004 441676 188604 441678
rect 224004 441676 224604 441678
rect 260004 441676 260604 441678
rect 296004 441676 296604 441678
rect 332004 441676 332604 441678
rect 368004 441676 368604 441678
rect 404004 441676 404604 441678
rect 440004 441676 440604 441678
rect 476004 441676 476604 441678
rect 512004 441676 512604 441678
rect 548004 441676 548604 441678
rect 589000 441676 589600 441678
rect -6596 441654 590520 441676
rect -6596 441418 -5494 441654
rect -5258 441418 8186 441654
rect 8422 441418 44186 441654
rect 44422 441418 80186 441654
rect 80422 441418 116186 441654
rect 116422 441418 152186 441654
rect 152422 441418 188186 441654
rect 188422 441418 224186 441654
rect 224422 441418 260186 441654
rect 260422 441418 296186 441654
rect 296422 441418 332186 441654
rect 332422 441418 368186 441654
rect 368422 441418 404186 441654
rect 404422 441418 440186 441654
rect 440422 441418 476186 441654
rect 476422 441418 512186 441654
rect 512422 441418 548186 441654
rect 548422 441418 589182 441654
rect 589418 441418 590520 441654
rect -6596 441334 590520 441418
rect -6596 441098 -5494 441334
rect -5258 441098 8186 441334
rect 8422 441098 44186 441334
rect 44422 441098 80186 441334
rect 80422 441098 116186 441334
rect 116422 441098 152186 441334
rect 152422 441098 188186 441334
rect 188422 441098 224186 441334
rect 224422 441098 260186 441334
rect 260422 441098 296186 441334
rect 296422 441098 332186 441334
rect 332422 441098 368186 441334
rect 368422 441098 404186 441334
rect 404422 441098 440186 441334
rect 440422 441098 476186 441334
rect 476422 441098 512186 441334
rect 512422 441098 548186 441334
rect 548422 441098 589182 441334
rect 589418 441098 590520 441334
rect -6596 441076 590520 441098
rect -5676 441074 -5076 441076
rect 8004 441074 8604 441076
rect 44004 441074 44604 441076
rect 80004 441074 80604 441076
rect 116004 441074 116604 441076
rect 152004 441074 152604 441076
rect 188004 441074 188604 441076
rect 224004 441074 224604 441076
rect 260004 441074 260604 441076
rect 296004 441074 296604 441076
rect 332004 441074 332604 441076
rect 368004 441074 368604 441076
rect 404004 441074 404604 441076
rect 440004 441074 440604 441076
rect 476004 441074 476604 441076
rect 512004 441074 512604 441076
rect 548004 441074 548604 441076
rect 589000 441074 589600 441076
rect -3836 438076 -3236 438078
rect 4404 438076 5004 438078
rect 40404 438076 41004 438078
rect 76404 438076 77004 438078
rect 112404 438076 113004 438078
rect 148404 438076 149004 438078
rect 184404 438076 185004 438078
rect 220404 438076 221004 438078
rect 256404 438076 257004 438078
rect 292404 438076 293004 438078
rect 328404 438076 329004 438078
rect 364404 438076 365004 438078
rect 400404 438076 401004 438078
rect 436404 438076 437004 438078
rect 472404 438076 473004 438078
rect 508404 438076 509004 438078
rect 544404 438076 545004 438078
rect 580404 438076 581004 438078
rect 587160 438076 587760 438078
rect -4756 438054 588680 438076
rect -4756 437818 -3654 438054
rect -3418 437818 4586 438054
rect 4822 437818 40586 438054
rect 40822 437818 76586 438054
rect 76822 437818 112586 438054
rect 112822 437818 148586 438054
rect 148822 437818 184586 438054
rect 184822 437818 220586 438054
rect 220822 437818 256586 438054
rect 256822 437818 292586 438054
rect 292822 437818 328586 438054
rect 328822 437818 364586 438054
rect 364822 437818 400586 438054
rect 400822 437818 436586 438054
rect 436822 437818 472586 438054
rect 472822 437818 508586 438054
rect 508822 437818 544586 438054
rect 544822 437818 580586 438054
rect 580822 437818 587342 438054
rect 587578 437818 588680 438054
rect -4756 437734 588680 437818
rect -4756 437498 -3654 437734
rect -3418 437498 4586 437734
rect 4822 437498 40586 437734
rect 40822 437498 76586 437734
rect 76822 437498 112586 437734
rect 112822 437498 148586 437734
rect 148822 437498 184586 437734
rect 184822 437498 220586 437734
rect 220822 437498 256586 437734
rect 256822 437498 292586 437734
rect 292822 437498 328586 437734
rect 328822 437498 364586 437734
rect 364822 437498 400586 437734
rect 400822 437498 436586 437734
rect 436822 437498 472586 437734
rect 472822 437498 508586 437734
rect 508822 437498 544586 437734
rect 544822 437498 580586 437734
rect 580822 437498 587342 437734
rect 587578 437498 588680 437734
rect -4756 437476 588680 437498
rect -3836 437474 -3236 437476
rect 4404 437474 5004 437476
rect 40404 437474 41004 437476
rect 76404 437474 77004 437476
rect 112404 437474 113004 437476
rect 148404 437474 149004 437476
rect 184404 437474 185004 437476
rect 220404 437474 221004 437476
rect 256404 437474 257004 437476
rect 292404 437474 293004 437476
rect 328404 437474 329004 437476
rect 364404 437474 365004 437476
rect 400404 437474 401004 437476
rect 436404 437474 437004 437476
rect 472404 437474 473004 437476
rect 508404 437474 509004 437476
rect 544404 437474 545004 437476
rect 580404 437474 581004 437476
rect 587160 437474 587760 437476
rect -1996 434476 -1396 434478
rect 804 434476 1404 434478
rect 36804 434476 37404 434478
rect 72804 434476 73404 434478
rect 108804 434476 109404 434478
rect 144804 434476 145404 434478
rect 180804 434476 181404 434478
rect 216804 434476 217404 434478
rect 252804 434476 253404 434478
rect 288804 434476 289404 434478
rect 324804 434476 325404 434478
rect 360804 434476 361404 434478
rect 396804 434476 397404 434478
rect 432804 434476 433404 434478
rect 468804 434476 469404 434478
rect 504804 434476 505404 434478
rect 540804 434476 541404 434478
rect 576804 434476 577404 434478
rect 585320 434476 585920 434478
rect -2916 434454 586840 434476
rect -2916 434218 -1814 434454
rect -1578 434218 986 434454
rect 1222 434218 36986 434454
rect 37222 434218 72986 434454
rect 73222 434218 108986 434454
rect 109222 434218 144986 434454
rect 145222 434218 180986 434454
rect 181222 434218 216986 434454
rect 217222 434218 252986 434454
rect 253222 434218 288986 434454
rect 289222 434218 324986 434454
rect 325222 434218 360986 434454
rect 361222 434218 396986 434454
rect 397222 434218 432986 434454
rect 433222 434218 468986 434454
rect 469222 434218 504986 434454
rect 505222 434218 540986 434454
rect 541222 434218 576986 434454
rect 577222 434218 585502 434454
rect 585738 434218 586840 434454
rect -2916 434134 586840 434218
rect -2916 433898 -1814 434134
rect -1578 433898 986 434134
rect 1222 433898 36986 434134
rect 37222 433898 72986 434134
rect 73222 433898 108986 434134
rect 109222 433898 144986 434134
rect 145222 433898 180986 434134
rect 181222 433898 216986 434134
rect 217222 433898 252986 434134
rect 253222 433898 288986 434134
rect 289222 433898 324986 434134
rect 325222 433898 360986 434134
rect 361222 433898 396986 434134
rect 397222 433898 432986 434134
rect 433222 433898 468986 434134
rect 469222 433898 504986 434134
rect 505222 433898 540986 434134
rect 541222 433898 576986 434134
rect 577222 433898 585502 434134
rect 585738 433898 586840 434134
rect -2916 433876 586840 433898
rect -1996 433874 -1396 433876
rect 804 433874 1404 433876
rect 36804 433874 37404 433876
rect 72804 433874 73404 433876
rect 108804 433874 109404 433876
rect 144804 433874 145404 433876
rect 180804 433874 181404 433876
rect 216804 433874 217404 433876
rect 252804 433874 253404 433876
rect 288804 433874 289404 433876
rect 324804 433874 325404 433876
rect 360804 433874 361404 433876
rect 396804 433874 397404 433876
rect 432804 433874 433404 433876
rect 468804 433874 469404 433876
rect 504804 433874 505404 433876
rect 540804 433874 541404 433876
rect 576804 433874 577404 433876
rect 585320 433874 585920 433876
rect -8436 427276 -7836 427278
rect 29604 427276 30204 427278
rect 65604 427276 66204 427278
rect 101604 427276 102204 427278
rect 137604 427276 138204 427278
rect 173604 427276 174204 427278
rect 209604 427276 210204 427278
rect 245604 427276 246204 427278
rect 281604 427276 282204 427278
rect 317604 427276 318204 427278
rect 353604 427276 354204 427278
rect 389604 427276 390204 427278
rect 425604 427276 426204 427278
rect 461604 427276 462204 427278
rect 497604 427276 498204 427278
rect 533604 427276 534204 427278
rect 569604 427276 570204 427278
rect 591760 427276 592360 427278
rect -8436 427254 592360 427276
rect -8436 427018 -8254 427254
rect -8018 427018 29786 427254
rect 30022 427018 65786 427254
rect 66022 427018 101786 427254
rect 102022 427018 137786 427254
rect 138022 427018 173786 427254
rect 174022 427018 209786 427254
rect 210022 427018 245786 427254
rect 246022 427018 281786 427254
rect 282022 427018 317786 427254
rect 318022 427018 353786 427254
rect 354022 427018 389786 427254
rect 390022 427018 425786 427254
rect 426022 427018 461786 427254
rect 462022 427018 497786 427254
rect 498022 427018 533786 427254
rect 534022 427018 569786 427254
rect 570022 427018 591942 427254
rect 592178 427018 592360 427254
rect -8436 426934 592360 427018
rect -8436 426698 -8254 426934
rect -8018 426698 29786 426934
rect 30022 426698 65786 426934
rect 66022 426698 101786 426934
rect 102022 426698 137786 426934
rect 138022 426698 173786 426934
rect 174022 426698 209786 426934
rect 210022 426698 245786 426934
rect 246022 426698 281786 426934
rect 282022 426698 317786 426934
rect 318022 426698 353786 426934
rect 354022 426698 389786 426934
rect 390022 426698 425786 426934
rect 426022 426698 461786 426934
rect 462022 426698 497786 426934
rect 498022 426698 533786 426934
rect 534022 426698 569786 426934
rect 570022 426698 591942 426934
rect 592178 426698 592360 426934
rect -8436 426676 592360 426698
rect -8436 426674 -7836 426676
rect 29604 426674 30204 426676
rect 65604 426674 66204 426676
rect 101604 426674 102204 426676
rect 137604 426674 138204 426676
rect 173604 426674 174204 426676
rect 209604 426674 210204 426676
rect 245604 426674 246204 426676
rect 281604 426674 282204 426676
rect 317604 426674 318204 426676
rect 353604 426674 354204 426676
rect 389604 426674 390204 426676
rect 425604 426674 426204 426676
rect 461604 426674 462204 426676
rect 497604 426674 498204 426676
rect 533604 426674 534204 426676
rect 569604 426674 570204 426676
rect 591760 426674 592360 426676
rect -6596 423676 -5996 423678
rect 26004 423676 26604 423678
rect 62004 423676 62604 423678
rect 98004 423676 98604 423678
rect 134004 423676 134604 423678
rect 170004 423676 170604 423678
rect 206004 423676 206604 423678
rect 242004 423676 242604 423678
rect 278004 423676 278604 423678
rect 314004 423676 314604 423678
rect 350004 423676 350604 423678
rect 386004 423676 386604 423678
rect 422004 423676 422604 423678
rect 458004 423676 458604 423678
rect 494004 423676 494604 423678
rect 530004 423676 530604 423678
rect 566004 423676 566604 423678
rect 589920 423676 590520 423678
rect -6596 423654 590520 423676
rect -6596 423418 -6414 423654
rect -6178 423418 26186 423654
rect 26422 423418 62186 423654
rect 62422 423418 98186 423654
rect 98422 423418 134186 423654
rect 134422 423418 170186 423654
rect 170422 423418 206186 423654
rect 206422 423418 242186 423654
rect 242422 423418 278186 423654
rect 278422 423418 314186 423654
rect 314422 423418 350186 423654
rect 350422 423418 386186 423654
rect 386422 423418 422186 423654
rect 422422 423418 458186 423654
rect 458422 423418 494186 423654
rect 494422 423418 530186 423654
rect 530422 423418 566186 423654
rect 566422 423418 590102 423654
rect 590338 423418 590520 423654
rect -6596 423334 590520 423418
rect -6596 423098 -6414 423334
rect -6178 423098 26186 423334
rect 26422 423098 62186 423334
rect 62422 423098 98186 423334
rect 98422 423098 134186 423334
rect 134422 423098 170186 423334
rect 170422 423098 206186 423334
rect 206422 423098 242186 423334
rect 242422 423098 278186 423334
rect 278422 423098 314186 423334
rect 314422 423098 350186 423334
rect 350422 423098 386186 423334
rect 386422 423098 422186 423334
rect 422422 423098 458186 423334
rect 458422 423098 494186 423334
rect 494422 423098 530186 423334
rect 530422 423098 566186 423334
rect 566422 423098 590102 423334
rect 590338 423098 590520 423334
rect -6596 423076 590520 423098
rect -6596 423074 -5996 423076
rect 26004 423074 26604 423076
rect 62004 423074 62604 423076
rect 98004 423074 98604 423076
rect 134004 423074 134604 423076
rect 170004 423074 170604 423076
rect 206004 423074 206604 423076
rect 242004 423074 242604 423076
rect 278004 423074 278604 423076
rect 314004 423074 314604 423076
rect 350004 423074 350604 423076
rect 386004 423074 386604 423076
rect 422004 423074 422604 423076
rect 458004 423074 458604 423076
rect 494004 423074 494604 423076
rect 530004 423074 530604 423076
rect 566004 423074 566604 423076
rect 589920 423074 590520 423076
rect -4756 420076 -4156 420078
rect 22404 420076 23004 420078
rect 58404 420076 59004 420078
rect 94404 420076 95004 420078
rect 130404 420076 131004 420078
rect 166404 420076 167004 420078
rect 202404 420076 203004 420078
rect 238404 420076 239004 420078
rect 274404 420076 275004 420078
rect 310404 420076 311004 420078
rect 346404 420076 347004 420078
rect 382404 420076 383004 420078
rect 418404 420076 419004 420078
rect 454404 420076 455004 420078
rect 490404 420076 491004 420078
rect 526404 420076 527004 420078
rect 562404 420076 563004 420078
rect 588080 420076 588680 420078
rect -4756 420054 588680 420076
rect -4756 419818 -4574 420054
rect -4338 419818 22586 420054
rect 22822 419818 58586 420054
rect 58822 419818 94586 420054
rect 94822 419818 130586 420054
rect 130822 419818 166586 420054
rect 166822 419818 202586 420054
rect 202822 419818 238586 420054
rect 238822 419818 274586 420054
rect 274822 419818 310586 420054
rect 310822 419818 346586 420054
rect 346822 419818 382586 420054
rect 382822 419818 418586 420054
rect 418822 419818 454586 420054
rect 454822 419818 490586 420054
rect 490822 419818 526586 420054
rect 526822 419818 562586 420054
rect 562822 419818 588262 420054
rect 588498 419818 588680 420054
rect -4756 419734 588680 419818
rect -4756 419498 -4574 419734
rect -4338 419498 22586 419734
rect 22822 419498 58586 419734
rect 58822 419498 94586 419734
rect 94822 419498 130586 419734
rect 130822 419498 166586 419734
rect 166822 419498 202586 419734
rect 202822 419498 238586 419734
rect 238822 419498 274586 419734
rect 274822 419498 310586 419734
rect 310822 419498 346586 419734
rect 346822 419498 382586 419734
rect 382822 419498 418586 419734
rect 418822 419498 454586 419734
rect 454822 419498 490586 419734
rect 490822 419498 526586 419734
rect 526822 419498 562586 419734
rect 562822 419498 588262 419734
rect 588498 419498 588680 419734
rect -4756 419476 588680 419498
rect -4756 419474 -4156 419476
rect 22404 419474 23004 419476
rect 58404 419474 59004 419476
rect 94404 419474 95004 419476
rect 130404 419474 131004 419476
rect 166404 419474 167004 419476
rect 202404 419474 203004 419476
rect 238404 419474 239004 419476
rect 274404 419474 275004 419476
rect 310404 419474 311004 419476
rect 346404 419474 347004 419476
rect 382404 419474 383004 419476
rect 418404 419474 419004 419476
rect 454404 419474 455004 419476
rect 490404 419474 491004 419476
rect 526404 419474 527004 419476
rect 562404 419474 563004 419476
rect 588080 419474 588680 419476
rect -2916 416476 -2316 416478
rect 18804 416476 19404 416478
rect 54804 416476 55404 416478
rect 90804 416476 91404 416478
rect 126804 416476 127404 416478
rect 162804 416476 163404 416478
rect 198804 416476 199404 416478
rect 234804 416476 235404 416478
rect 270804 416476 271404 416478
rect 306804 416476 307404 416478
rect 342804 416476 343404 416478
rect 378804 416476 379404 416478
rect 414804 416476 415404 416478
rect 450804 416476 451404 416478
rect 486804 416476 487404 416478
rect 522804 416476 523404 416478
rect 558804 416476 559404 416478
rect 586240 416476 586840 416478
rect -2916 416454 586840 416476
rect -2916 416218 -2734 416454
rect -2498 416218 18986 416454
rect 19222 416218 54986 416454
rect 55222 416218 90986 416454
rect 91222 416218 126986 416454
rect 127222 416218 162986 416454
rect 163222 416218 198986 416454
rect 199222 416218 234986 416454
rect 235222 416218 270986 416454
rect 271222 416218 306986 416454
rect 307222 416218 342986 416454
rect 343222 416218 378986 416454
rect 379222 416218 414986 416454
rect 415222 416218 450986 416454
rect 451222 416218 486986 416454
rect 487222 416218 522986 416454
rect 523222 416218 558986 416454
rect 559222 416218 586422 416454
rect 586658 416218 586840 416454
rect -2916 416134 586840 416218
rect -2916 415898 -2734 416134
rect -2498 415898 18986 416134
rect 19222 415898 54986 416134
rect 55222 415898 90986 416134
rect 91222 415898 126986 416134
rect 127222 415898 162986 416134
rect 163222 415898 198986 416134
rect 199222 415898 234986 416134
rect 235222 415898 270986 416134
rect 271222 415898 306986 416134
rect 307222 415898 342986 416134
rect 343222 415898 378986 416134
rect 379222 415898 414986 416134
rect 415222 415898 450986 416134
rect 451222 415898 486986 416134
rect 487222 415898 522986 416134
rect 523222 415898 558986 416134
rect 559222 415898 586422 416134
rect 586658 415898 586840 416134
rect -2916 415876 586840 415898
rect -2916 415874 -2316 415876
rect 18804 415874 19404 415876
rect 54804 415874 55404 415876
rect 90804 415874 91404 415876
rect 126804 415874 127404 415876
rect 162804 415874 163404 415876
rect 198804 415874 199404 415876
rect 234804 415874 235404 415876
rect 270804 415874 271404 415876
rect 306804 415874 307404 415876
rect 342804 415874 343404 415876
rect 378804 415874 379404 415876
rect 414804 415874 415404 415876
rect 450804 415874 451404 415876
rect 486804 415874 487404 415876
rect 522804 415874 523404 415876
rect 558804 415874 559404 415876
rect 586240 415874 586840 415876
rect -7516 409276 -6916 409278
rect 11604 409276 12204 409278
rect 47604 409276 48204 409278
rect 83604 409276 84204 409278
rect 119604 409276 120204 409278
rect 155604 409276 156204 409278
rect 191604 409276 192204 409278
rect 227604 409276 228204 409278
rect 263604 409276 264204 409278
rect 299604 409276 300204 409278
rect 335604 409276 336204 409278
rect 371604 409276 372204 409278
rect 407604 409276 408204 409278
rect 443604 409276 444204 409278
rect 479604 409276 480204 409278
rect 515604 409276 516204 409278
rect 551604 409276 552204 409278
rect 590840 409276 591440 409278
rect -8436 409254 592360 409276
rect -8436 409018 -7334 409254
rect -7098 409018 11786 409254
rect 12022 409018 47786 409254
rect 48022 409018 83786 409254
rect 84022 409018 119786 409254
rect 120022 409018 155786 409254
rect 156022 409018 191786 409254
rect 192022 409018 227786 409254
rect 228022 409018 263786 409254
rect 264022 409018 299786 409254
rect 300022 409018 335786 409254
rect 336022 409018 371786 409254
rect 372022 409018 407786 409254
rect 408022 409018 443786 409254
rect 444022 409018 479786 409254
rect 480022 409018 515786 409254
rect 516022 409018 551786 409254
rect 552022 409018 591022 409254
rect 591258 409018 592360 409254
rect -8436 408934 592360 409018
rect -8436 408698 -7334 408934
rect -7098 408698 11786 408934
rect 12022 408698 47786 408934
rect 48022 408698 83786 408934
rect 84022 408698 119786 408934
rect 120022 408698 155786 408934
rect 156022 408698 191786 408934
rect 192022 408698 227786 408934
rect 228022 408698 263786 408934
rect 264022 408698 299786 408934
rect 300022 408698 335786 408934
rect 336022 408698 371786 408934
rect 372022 408698 407786 408934
rect 408022 408698 443786 408934
rect 444022 408698 479786 408934
rect 480022 408698 515786 408934
rect 516022 408698 551786 408934
rect 552022 408698 591022 408934
rect 591258 408698 592360 408934
rect -8436 408676 592360 408698
rect -7516 408674 -6916 408676
rect 11604 408674 12204 408676
rect 47604 408674 48204 408676
rect 83604 408674 84204 408676
rect 119604 408674 120204 408676
rect 155604 408674 156204 408676
rect 191604 408674 192204 408676
rect 227604 408674 228204 408676
rect 263604 408674 264204 408676
rect 299604 408674 300204 408676
rect 335604 408674 336204 408676
rect 371604 408674 372204 408676
rect 407604 408674 408204 408676
rect 443604 408674 444204 408676
rect 479604 408674 480204 408676
rect 515604 408674 516204 408676
rect 551604 408674 552204 408676
rect 590840 408674 591440 408676
rect -5676 405676 -5076 405678
rect 8004 405676 8604 405678
rect 44004 405676 44604 405678
rect 80004 405676 80604 405678
rect 116004 405676 116604 405678
rect 152004 405676 152604 405678
rect 188004 405676 188604 405678
rect 224004 405676 224604 405678
rect 260004 405676 260604 405678
rect 296004 405676 296604 405678
rect 332004 405676 332604 405678
rect 368004 405676 368604 405678
rect 404004 405676 404604 405678
rect 440004 405676 440604 405678
rect 476004 405676 476604 405678
rect 512004 405676 512604 405678
rect 548004 405676 548604 405678
rect 589000 405676 589600 405678
rect -6596 405654 590520 405676
rect -6596 405418 -5494 405654
rect -5258 405418 8186 405654
rect 8422 405418 44186 405654
rect 44422 405418 80186 405654
rect 80422 405418 116186 405654
rect 116422 405418 152186 405654
rect 152422 405418 188186 405654
rect 188422 405418 224186 405654
rect 224422 405418 260186 405654
rect 260422 405418 296186 405654
rect 296422 405418 332186 405654
rect 332422 405418 368186 405654
rect 368422 405418 404186 405654
rect 404422 405418 440186 405654
rect 440422 405418 476186 405654
rect 476422 405418 512186 405654
rect 512422 405418 548186 405654
rect 548422 405418 589182 405654
rect 589418 405418 590520 405654
rect -6596 405334 590520 405418
rect -6596 405098 -5494 405334
rect -5258 405098 8186 405334
rect 8422 405098 44186 405334
rect 44422 405098 80186 405334
rect 80422 405098 116186 405334
rect 116422 405098 152186 405334
rect 152422 405098 188186 405334
rect 188422 405098 224186 405334
rect 224422 405098 260186 405334
rect 260422 405098 296186 405334
rect 296422 405098 332186 405334
rect 332422 405098 368186 405334
rect 368422 405098 404186 405334
rect 404422 405098 440186 405334
rect 440422 405098 476186 405334
rect 476422 405098 512186 405334
rect 512422 405098 548186 405334
rect 548422 405098 589182 405334
rect 589418 405098 590520 405334
rect -6596 405076 590520 405098
rect -5676 405074 -5076 405076
rect 8004 405074 8604 405076
rect 44004 405074 44604 405076
rect 80004 405074 80604 405076
rect 116004 405074 116604 405076
rect 152004 405074 152604 405076
rect 188004 405074 188604 405076
rect 224004 405074 224604 405076
rect 260004 405074 260604 405076
rect 296004 405074 296604 405076
rect 332004 405074 332604 405076
rect 368004 405074 368604 405076
rect 404004 405074 404604 405076
rect 440004 405074 440604 405076
rect 476004 405074 476604 405076
rect 512004 405074 512604 405076
rect 548004 405074 548604 405076
rect 589000 405074 589600 405076
rect -3836 402076 -3236 402078
rect 4404 402076 5004 402078
rect 40404 402076 41004 402078
rect 76404 402076 77004 402078
rect 112404 402076 113004 402078
rect 148404 402076 149004 402078
rect 184404 402076 185004 402078
rect 220404 402076 221004 402078
rect 256404 402076 257004 402078
rect 292404 402076 293004 402078
rect 328404 402076 329004 402078
rect 364404 402076 365004 402078
rect 400404 402076 401004 402078
rect 436404 402076 437004 402078
rect 472404 402076 473004 402078
rect 508404 402076 509004 402078
rect 544404 402076 545004 402078
rect 580404 402076 581004 402078
rect 587160 402076 587760 402078
rect -4756 402054 588680 402076
rect -4756 401818 -3654 402054
rect -3418 401818 4586 402054
rect 4822 401818 40586 402054
rect 40822 401818 76586 402054
rect 76822 401818 112586 402054
rect 112822 401818 148586 402054
rect 148822 401818 184586 402054
rect 184822 401818 220586 402054
rect 220822 401818 256586 402054
rect 256822 401818 292586 402054
rect 292822 401818 328586 402054
rect 328822 401818 364586 402054
rect 364822 401818 400586 402054
rect 400822 401818 436586 402054
rect 436822 401818 472586 402054
rect 472822 401818 508586 402054
rect 508822 401818 544586 402054
rect 544822 401818 580586 402054
rect 580822 401818 587342 402054
rect 587578 401818 588680 402054
rect -4756 401734 588680 401818
rect -4756 401498 -3654 401734
rect -3418 401498 4586 401734
rect 4822 401498 40586 401734
rect 40822 401498 76586 401734
rect 76822 401498 112586 401734
rect 112822 401498 148586 401734
rect 148822 401498 184586 401734
rect 184822 401498 220586 401734
rect 220822 401498 256586 401734
rect 256822 401498 292586 401734
rect 292822 401498 328586 401734
rect 328822 401498 364586 401734
rect 364822 401498 400586 401734
rect 400822 401498 436586 401734
rect 436822 401498 472586 401734
rect 472822 401498 508586 401734
rect 508822 401498 544586 401734
rect 544822 401498 580586 401734
rect 580822 401498 587342 401734
rect 587578 401498 588680 401734
rect -4756 401476 588680 401498
rect -3836 401474 -3236 401476
rect 4404 401474 5004 401476
rect 40404 401474 41004 401476
rect 76404 401474 77004 401476
rect 112404 401474 113004 401476
rect 148404 401474 149004 401476
rect 184404 401474 185004 401476
rect 220404 401474 221004 401476
rect 256404 401474 257004 401476
rect 292404 401474 293004 401476
rect 328404 401474 329004 401476
rect 364404 401474 365004 401476
rect 400404 401474 401004 401476
rect 436404 401474 437004 401476
rect 472404 401474 473004 401476
rect 508404 401474 509004 401476
rect 544404 401474 545004 401476
rect 580404 401474 581004 401476
rect 587160 401474 587760 401476
rect -1996 398476 -1396 398478
rect 804 398476 1404 398478
rect 36804 398476 37404 398478
rect 72804 398476 73404 398478
rect 108804 398476 109404 398478
rect 144804 398476 145404 398478
rect 180804 398476 181404 398478
rect 216804 398476 217404 398478
rect 252804 398476 253404 398478
rect 288804 398476 289404 398478
rect 324804 398476 325404 398478
rect 360804 398476 361404 398478
rect 396804 398476 397404 398478
rect 432804 398476 433404 398478
rect 468804 398476 469404 398478
rect 504804 398476 505404 398478
rect 540804 398476 541404 398478
rect 576804 398476 577404 398478
rect 585320 398476 585920 398478
rect -2916 398454 586840 398476
rect -2916 398218 -1814 398454
rect -1578 398218 986 398454
rect 1222 398218 36986 398454
rect 37222 398218 72986 398454
rect 73222 398218 108986 398454
rect 109222 398218 144986 398454
rect 145222 398218 180986 398454
rect 181222 398218 216986 398454
rect 217222 398218 252986 398454
rect 253222 398218 288986 398454
rect 289222 398218 324986 398454
rect 325222 398218 360986 398454
rect 361222 398218 396986 398454
rect 397222 398218 432986 398454
rect 433222 398218 468986 398454
rect 469222 398218 504986 398454
rect 505222 398218 540986 398454
rect 541222 398218 576986 398454
rect 577222 398218 585502 398454
rect 585738 398218 586840 398454
rect -2916 398134 586840 398218
rect -2916 397898 -1814 398134
rect -1578 397898 986 398134
rect 1222 397898 36986 398134
rect 37222 397898 72986 398134
rect 73222 397898 108986 398134
rect 109222 397898 144986 398134
rect 145222 397898 180986 398134
rect 181222 397898 216986 398134
rect 217222 397898 252986 398134
rect 253222 397898 288986 398134
rect 289222 397898 324986 398134
rect 325222 397898 360986 398134
rect 361222 397898 396986 398134
rect 397222 397898 432986 398134
rect 433222 397898 468986 398134
rect 469222 397898 504986 398134
rect 505222 397898 540986 398134
rect 541222 397898 576986 398134
rect 577222 397898 585502 398134
rect 585738 397898 586840 398134
rect -2916 397876 586840 397898
rect -1996 397874 -1396 397876
rect 804 397874 1404 397876
rect 36804 397874 37404 397876
rect 72804 397874 73404 397876
rect 108804 397874 109404 397876
rect 144804 397874 145404 397876
rect 180804 397874 181404 397876
rect 216804 397874 217404 397876
rect 252804 397874 253404 397876
rect 288804 397874 289404 397876
rect 324804 397874 325404 397876
rect 360804 397874 361404 397876
rect 396804 397874 397404 397876
rect 432804 397874 433404 397876
rect 468804 397874 469404 397876
rect 504804 397874 505404 397876
rect 540804 397874 541404 397876
rect 576804 397874 577404 397876
rect 585320 397874 585920 397876
rect -8436 391276 -7836 391278
rect 29604 391276 30204 391278
rect 65604 391276 66204 391278
rect 101604 391276 102204 391278
rect 137604 391276 138204 391278
rect 173604 391276 174204 391278
rect 209604 391276 210204 391278
rect 245604 391276 246204 391278
rect 281604 391276 282204 391278
rect 317604 391276 318204 391278
rect 353604 391276 354204 391278
rect 389604 391276 390204 391278
rect 425604 391276 426204 391278
rect 461604 391276 462204 391278
rect 497604 391276 498204 391278
rect 533604 391276 534204 391278
rect 569604 391276 570204 391278
rect 591760 391276 592360 391278
rect -8436 391254 592360 391276
rect -8436 391018 -8254 391254
rect -8018 391018 29786 391254
rect 30022 391018 65786 391254
rect 66022 391018 101786 391254
rect 102022 391018 137786 391254
rect 138022 391018 173786 391254
rect 174022 391018 209786 391254
rect 210022 391018 245786 391254
rect 246022 391018 281786 391254
rect 282022 391018 317786 391254
rect 318022 391018 353786 391254
rect 354022 391018 389786 391254
rect 390022 391018 425786 391254
rect 426022 391018 461786 391254
rect 462022 391018 497786 391254
rect 498022 391018 533786 391254
rect 534022 391018 569786 391254
rect 570022 391018 591942 391254
rect 592178 391018 592360 391254
rect -8436 390934 592360 391018
rect -8436 390698 -8254 390934
rect -8018 390698 29786 390934
rect 30022 390698 65786 390934
rect 66022 390698 101786 390934
rect 102022 390698 137786 390934
rect 138022 390698 173786 390934
rect 174022 390698 209786 390934
rect 210022 390698 245786 390934
rect 246022 390698 281786 390934
rect 282022 390698 317786 390934
rect 318022 390698 353786 390934
rect 354022 390698 389786 390934
rect 390022 390698 425786 390934
rect 426022 390698 461786 390934
rect 462022 390698 497786 390934
rect 498022 390698 533786 390934
rect 534022 390698 569786 390934
rect 570022 390698 591942 390934
rect 592178 390698 592360 390934
rect -8436 390676 592360 390698
rect -8436 390674 -7836 390676
rect 29604 390674 30204 390676
rect 65604 390674 66204 390676
rect 101604 390674 102204 390676
rect 137604 390674 138204 390676
rect 173604 390674 174204 390676
rect 209604 390674 210204 390676
rect 245604 390674 246204 390676
rect 281604 390674 282204 390676
rect 317604 390674 318204 390676
rect 353604 390674 354204 390676
rect 389604 390674 390204 390676
rect 425604 390674 426204 390676
rect 461604 390674 462204 390676
rect 497604 390674 498204 390676
rect 533604 390674 534204 390676
rect 569604 390674 570204 390676
rect 591760 390674 592360 390676
rect -6596 387676 -5996 387678
rect 26004 387676 26604 387678
rect 62004 387676 62604 387678
rect 98004 387676 98604 387678
rect 134004 387676 134604 387678
rect 170004 387676 170604 387678
rect 206004 387676 206604 387678
rect 242004 387676 242604 387678
rect 278004 387676 278604 387678
rect 314004 387676 314604 387678
rect 350004 387676 350604 387678
rect 386004 387676 386604 387678
rect 422004 387676 422604 387678
rect 458004 387676 458604 387678
rect 494004 387676 494604 387678
rect 530004 387676 530604 387678
rect 566004 387676 566604 387678
rect 589920 387676 590520 387678
rect -6596 387654 590520 387676
rect -6596 387418 -6414 387654
rect -6178 387418 26186 387654
rect 26422 387418 62186 387654
rect 62422 387418 98186 387654
rect 98422 387418 134186 387654
rect 134422 387418 170186 387654
rect 170422 387418 206186 387654
rect 206422 387418 242186 387654
rect 242422 387418 278186 387654
rect 278422 387418 314186 387654
rect 314422 387418 350186 387654
rect 350422 387418 386186 387654
rect 386422 387418 422186 387654
rect 422422 387418 458186 387654
rect 458422 387418 494186 387654
rect 494422 387418 530186 387654
rect 530422 387418 566186 387654
rect 566422 387418 590102 387654
rect 590338 387418 590520 387654
rect -6596 387334 590520 387418
rect -6596 387098 -6414 387334
rect -6178 387098 26186 387334
rect 26422 387098 62186 387334
rect 62422 387098 98186 387334
rect 98422 387098 134186 387334
rect 134422 387098 170186 387334
rect 170422 387098 206186 387334
rect 206422 387098 242186 387334
rect 242422 387098 278186 387334
rect 278422 387098 314186 387334
rect 314422 387098 350186 387334
rect 350422 387098 386186 387334
rect 386422 387098 422186 387334
rect 422422 387098 458186 387334
rect 458422 387098 494186 387334
rect 494422 387098 530186 387334
rect 530422 387098 566186 387334
rect 566422 387098 590102 387334
rect 590338 387098 590520 387334
rect -6596 387076 590520 387098
rect -6596 387074 -5996 387076
rect 26004 387074 26604 387076
rect 62004 387074 62604 387076
rect 98004 387074 98604 387076
rect 134004 387074 134604 387076
rect 170004 387074 170604 387076
rect 206004 387074 206604 387076
rect 242004 387074 242604 387076
rect 278004 387074 278604 387076
rect 314004 387074 314604 387076
rect 350004 387074 350604 387076
rect 386004 387074 386604 387076
rect 422004 387074 422604 387076
rect 458004 387074 458604 387076
rect 494004 387074 494604 387076
rect 530004 387074 530604 387076
rect 566004 387074 566604 387076
rect 589920 387074 590520 387076
rect -4756 384076 -4156 384078
rect 22404 384076 23004 384078
rect 58404 384076 59004 384078
rect 94404 384076 95004 384078
rect 130404 384076 131004 384078
rect 166404 384076 167004 384078
rect 202404 384076 203004 384078
rect 238404 384076 239004 384078
rect 274404 384076 275004 384078
rect 310404 384076 311004 384078
rect 346404 384076 347004 384078
rect 382404 384076 383004 384078
rect 418404 384076 419004 384078
rect 454404 384076 455004 384078
rect 490404 384076 491004 384078
rect 526404 384076 527004 384078
rect 562404 384076 563004 384078
rect 588080 384076 588680 384078
rect -4756 384054 588680 384076
rect -4756 383818 -4574 384054
rect -4338 383818 22586 384054
rect 22822 383818 58586 384054
rect 58822 383818 94586 384054
rect 94822 383818 130586 384054
rect 130822 383818 166586 384054
rect 166822 383818 202586 384054
rect 202822 383818 238586 384054
rect 238822 383818 274586 384054
rect 274822 383818 310586 384054
rect 310822 383818 346586 384054
rect 346822 383818 382586 384054
rect 382822 383818 418586 384054
rect 418822 383818 454586 384054
rect 454822 383818 490586 384054
rect 490822 383818 526586 384054
rect 526822 383818 562586 384054
rect 562822 383818 588262 384054
rect 588498 383818 588680 384054
rect -4756 383734 588680 383818
rect -4756 383498 -4574 383734
rect -4338 383498 22586 383734
rect 22822 383498 58586 383734
rect 58822 383498 94586 383734
rect 94822 383498 130586 383734
rect 130822 383498 166586 383734
rect 166822 383498 202586 383734
rect 202822 383498 238586 383734
rect 238822 383498 274586 383734
rect 274822 383498 310586 383734
rect 310822 383498 346586 383734
rect 346822 383498 382586 383734
rect 382822 383498 418586 383734
rect 418822 383498 454586 383734
rect 454822 383498 490586 383734
rect 490822 383498 526586 383734
rect 526822 383498 562586 383734
rect 562822 383498 588262 383734
rect 588498 383498 588680 383734
rect -4756 383476 588680 383498
rect -4756 383474 -4156 383476
rect 22404 383474 23004 383476
rect 58404 383474 59004 383476
rect 94404 383474 95004 383476
rect 130404 383474 131004 383476
rect 166404 383474 167004 383476
rect 202404 383474 203004 383476
rect 238404 383474 239004 383476
rect 274404 383474 275004 383476
rect 310404 383474 311004 383476
rect 346404 383474 347004 383476
rect 382404 383474 383004 383476
rect 418404 383474 419004 383476
rect 454404 383474 455004 383476
rect 490404 383474 491004 383476
rect 526404 383474 527004 383476
rect 562404 383474 563004 383476
rect 588080 383474 588680 383476
rect -2916 380476 -2316 380478
rect 18804 380476 19404 380478
rect 54804 380476 55404 380478
rect 90804 380476 91404 380478
rect 126804 380476 127404 380478
rect 162804 380476 163404 380478
rect 198804 380476 199404 380478
rect 234804 380476 235404 380478
rect 270804 380476 271404 380478
rect 306804 380476 307404 380478
rect 342804 380476 343404 380478
rect 378804 380476 379404 380478
rect 414804 380476 415404 380478
rect 450804 380476 451404 380478
rect 486804 380476 487404 380478
rect 522804 380476 523404 380478
rect 558804 380476 559404 380478
rect 586240 380476 586840 380478
rect -2916 380454 586840 380476
rect -2916 380218 -2734 380454
rect -2498 380218 18986 380454
rect 19222 380218 54986 380454
rect 55222 380218 90986 380454
rect 91222 380218 126986 380454
rect 127222 380218 162986 380454
rect 163222 380218 198986 380454
rect 199222 380218 234986 380454
rect 235222 380218 270986 380454
rect 271222 380218 306986 380454
rect 307222 380218 342986 380454
rect 343222 380218 378986 380454
rect 379222 380218 414986 380454
rect 415222 380218 450986 380454
rect 451222 380218 486986 380454
rect 487222 380218 522986 380454
rect 523222 380218 558986 380454
rect 559222 380218 586422 380454
rect 586658 380218 586840 380454
rect -2916 380134 586840 380218
rect -2916 379898 -2734 380134
rect -2498 379898 18986 380134
rect 19222 379898 54986 380134
rect 55222 379898 90986 380134
rect 91222 379898 126986 380134
rect 127222 379898 162986 380134
rect 163222 379898 198986 380134
rect 199222 379898 234986 380134
rect 235222 379898 270986 380134
rect 271222 379898 306986 380134
rect 307222 379898 342986 380134
rect 343222 379898 378986 380134
rect 379222 379898 414986 380134
rect 415222 379898 450986 380134
rect 451222 379898 486986 380134
rect 487222 379898 522986 380134
rect 523222 379898 558986 380134
rect 559222 379898 586422 380134
rect 586658 379898 586840 380134
rect -2916 379876 586840 379898
rect -2916 379874 -2316 379876
rect 18804 379874 19404 379876
rect 54804 379874 55404 379876
rect 90804 379874 91404 379876
rect 126804 379874 127404 379876
rect 162804 379874 163404 379876
rect 198804 379874 199404 379876
rect 234804 379874 235404 379876
rect 270804 379874 271404 379876
rect 306804 379874 307404 379876
rect 342804 379874 343404 379876
rect 378804 379874 379404 379876
rect 414804 379874 415404 379876
rect 450804 379874 451404 379876
rect 486804 379874 487404 379876
rect 522804 379874 523404 379876
rect 558804 379874 559404 379876
rect 586240 379874 586840 379876
rect -7516 373276 -6916 373278
rect 11604 373276 12204 373278
rect 47604 373276 48204 373278
rect 83604 373276 84204 373278
rect 119604 373276 120204 373278
rect 155604 373276 156204 373278
rect 191604 373276 192204 373278
rect 227604 373276 228204 373278
rect 263604 373276 264204 373278
rect 299604 373276 300204 373278
rect 335604 373276 336204 373278
rect 371604 373276 372204 373278
rect 407604 373276 408204 373278
rect 443604 373276 444204 373278
rect 479604 373276 480204 373278
rect 515604 373276 516204 373278
rect 551604 373276 552204 373278
rect 590840 373276 591440 373278
rect -8436 373254 592360 373276
rect -8436 373018 -7334 373254
rect -7098 373018 11786 373254
rect 12022 373018 47786 373254
rect 48022 373018 83786 373254
rect 84022 373018 119786 373254
rect 120022 373018 155786 373254
rect 156022 373018 191786 373254
rect 192022 373018 227786 373254
rect 228022 373018 263786 373254
rect 264022 373018 299786 373254
rect 300022 373018 335786 373254
rect 336022 373018 371786 373254
rect 372022 373018 407786 373254
rect 408022 373018 443786 373254
rect 444022 373018 479786 373254
rect 480022 373018 515786 373254
rect 516022 373018 551786 373254
rect 552022 373018 591022 373254
rect 591258 373018 592360 373254
rect -8436 372934 592360 373018
rect -8436 372698 -7334 372934
rect -7098 372698 11786 372934
rect 12022 372698 47786 372934
rect 48022 372698 83786 372934
rect 84022 372698 119786 372934
rect 120022 372698 155786 372934
rect 156022 372698 191786 372934
rect 192022 372698 227786 372934
rect 228022 372698 263786 372934
rect 264022 372698 299786 372934
rect 300022 372698 335786 372934
rect 336022 372698 371786 372934
rect 372022 372698 407786 372934
rect 408022 372698 443786 372934
rect 444022 372698 479786 372934
rect 480022 372698 515786 372934
rect 516022 372698 551786 372934
rect 552022 372698 591022 372934
rect 591258 372698 592360 372934
rect -8436 372676 592360 372698
rect -7516 372674 -6916 372676
rect 11604 372674 12204 372676
rect 47604 372674 48204 372676
rect 83604 372674 84204 372676
rect 119604 372674 120204 372676
rect 155604 372674 156204 372676
rect 191604 372674 192204 372676
rect 227604 372674 228204 372676
rect 263604 372674 264204 372676
rect 299604 372674 300204 372676
rect 335604 372674 336204 372676
rect 371604 372674 372204 372676
rect 407604 372674 408204 372676
rect 443604 372674 444204 372676
rect 479604 372674 480204 372676
rect 515604 372674 516204 372676
rect 551604 372674 552204 372676
rect 590840 372674 591440 372676
rect -5676 369676 -5076 369678
rect 8004 369676 8604 369678
rect 44004 369676 44604 369678
rect 80004 369676 80604 369678
rect 116004 369676 116604 369678
rect 152004 369676 152604 369678
rect 188004 369676 188604 369678
rect 224004 369676 224604 369678
rect 260004 369676 260604 369678
rect 296004 369676 296604 369678
rect 332004 369676 332604 369678
rect 368004 369676 368604 369678
rect 404004 369676 404604 369678
rect 440004 369676 440604 369678
rect 476004 369676 476604 369678
rect 512004 369676 512604 369678
rect 548004 369676 548604 369678
rect 589000 369676 589600 369678
rect -6596 369654 590520 369676
rect -6596 369418 -5494 369654
rect -5258 369418 8186 369654
rect 8422 369418 44186 369654
rect 44422 369418 80186 369654
rect 80422 369418 116186 369654
rect 116422 369418 152186 369654
rect 152422 369418 188186 369654
rect 188422 369418 224186 369654
rect 224422 369418 260186 369654
rect 260422 369418 296186 369654
rect 296422 369418 332186 369654
rect 332422 369418 368186 369654
rect 368422 369418 404186 369654
rect 404422 369418 440186 369654
rect 440422 369418 476186 369654
rect 476422 369418 512186 369654
rect 512422 369418 548186 369654
rect 548422 369418 589182 369654
rect 589418 369418 590520 369654
rect -6596 369334 590520 369418
rect -6596 369098 -5494 369334
rect -5258 369098 8186 369334
rect 8422 369098 44186 369334
rect 44422 369098 80186 369334
rect 80422 369098 116186 369334
rect 116422 369098 152186 369334
rect 152422 369098 188186 369334
rect 188422 369098 224186 369334
rect 224422 369098 260186 369334
rect 260422 369098 296186 369334
rect 296422 369098 332186 369334
rect 332422 369098 368186 369334
rect 368422 369098 404186 369334
rect 404422 369098 440186 369334
rect 440422 369098 476186 369334
rect 476422 369098 512186 369334
rect 512422 369098 548186 369334
rect 548422 369098 589182 369334
rect 589418 369098 590520 369334
rect -6596 369076 590520 369098
rect -5676 369074 -5076 369076
rect 8004 369074 8604 369076
rect 44004 369074 44604 369076
rect 80004 369074 80604 369076
rect 116004 369074 116604 369076
rect 152004 369074 152604 369076
rect 188004 369074 188604 369076
rect 224004 369074 224604 369076
rect 260004 369074 260604 369076
rect 296004 369074 296604 369076
rect 332004 369074 332604 369076
rect 368004 369074 368604 369076
rect 404004 369074 404604 369076
rect 440004 369074 440604 369076
rect 476004 369074 476604 369076
rect 512004 369074 512604 369076
rect 548004 369074 548604 369076
rect 589000 369074 589600 369076
rect -3836 366076 -3236 366078
rect 4404 366076 5004 366078
rect 40404 366076 41004 366078
rect 76404 366076 77004 366078
rect 112404 366076 113004 366078
rect 148404 366076 149004 366078
rect 184404 366076 185004 366078
rect 220404 366076 221004 366078
rect 256404 366076 257004 366078
rect 292404 366076 293004 366078
rect 328404 366076 329004 366078
rect 364404 366076 365004 366078
rect 400404 366076 401004 366078
rect 436404 366076 437004 366078
rect 472404 366076 473004 366078
rect 508404 366076 509004 366078
rect 544404 366076 545004 366078
rect 580404 366076 581004 366078
rect 587160 366076 587760 366078
rect -4756 366054 588680 366076
rect -4756 365818 -3654 366054
rect -3418 365818 4586 366054
rect 4822 365818 40586 366054
rect 40822 365818 76586 366054
rect 76822 365818 112586 366054
rect 112822 365818 148586 366054
rect 148822 365818 184586 366054
rect 184822 365818 220586 366054
rect 220822 365818 256586 366054
rect 256822 365818 292586 366054
rect 292822 365818 328586 366054
rect 328822 365818 364586 366054
rect 364822 365818 400586 366054
rect 400822 365818 436586 366054
rect 436822 365818 472586 366054
rect 472822 365818 508586 366054
rect 508822 365818 544586 366054
rect 544822 365818 580586 366054
rect 580822 365818 587342 366054
rect 587578 365818 588680 366054
rect -4756 365734 588680 365818
rect -4756 365498 -3654 365734
rect -3418 365498 4586 365734
rect 4822 365498 40586 365734
rect 40822 365498 76586 365734
rect 76822 365498 112586 365734
rect 112822 365498 148586 365734
rect 148822 365498 184586 365734
rect 184822 365498 220586 365734
rect 220822 365498 256586 365734
rect 256822 365498 292586 365734
rect 292822 365498 328586 365734
rect 328822 365498 364586 365734
rect 364822 365498 400586 365734
rect 400822 365498 436586 365734
rect 436822 365498 472586 365734
rect 472822 365498 508586 365734
rect 508822 365498 544586 365734
rect 544822 365498 580586 365734
rect 580822 365498 587342 365734
rect 587578 365498 588680 365734
rect -4756 365476 588680 365498
rect -3836 365474 -3236 365476
rect 4404 365474 5004 365476
rect 40404 365474 41004 365476
rect 76404 365474 77004 365476
rect 112404 365474 113004 365476
rect 148404 365474 149004 365476
rect 184404 365474 185004 365476
rect 220404 365474 221004 365476
rect 256404 365474 257004 365476
rect 292404 365474 293004 365476
rect 328404 365474 329004 365476
rect 364404 365474 365004 365476
rect 400404 365474 401004 365476
rect 436404 365474 437004 365476
rect 472404 365474 473004 365476
rect 508404 365474 509004 365476
rect 544404 365474 545004 365476
rect 580404 365474 581004 365476
rect 587160 365474 587760 365476
rect -1996 362476 -1396 362478
rect 804 362476 1404 362478
rect 36804 362476 37404 362478
rect 72804 362476 73404 362478
rect 108804 362476 109404 362478
rect 144804 362476 145404 362478
rect 180804 362476 181404 362478
rect 216804 362476 217404 362478
rect 252804 362476 253404 362478
rect 288804 362476 289404 362478
rect 324804 362476 325404 362478
rect 360804 362476 361404 362478
rect 396804 362476 397404 362478
rect 432804 362476 433404 362478
rect 468804 362476 469404 362478
rect 504804 362476 505404 362478
rect 540804 362476 541404 362478
rect 576804 362476 577404 362478
rect 585320 362476 585920 362478
rect -2916 362454 586840 362476
rect -2916 362218 -1814 362454
rect -1578 362218 986 362454
rect 1222 362218 36986 362454
rect 37222 362218 72986 362454
rect 73222 362218 108986 362454
rect 109222 362218 144986 362454
rect 145222 362218 180986 362454
rect 181222 362218 216986 362454
rect 217222 362218 252986 362454
rect 253222 362218 288986 362454
rect 289222 362218 324986 362454
rect 325222 362218 360986 362454
rect 361222 362218 396986 362454
rect 397222 362218 432986 362454
rect 433222 362218 468986 362454
rect 469222 362218 504986 362454
rect 505222 362218 540986 362454
rect 541222 362218 576986 362454
rect 577222 362218 585502 362454
rect 585738 362218 586840 362454
rect -2916 362134 586840 362218
rect -2916 361898 -1814 362134
rect -1578 361898 986 362134
rect 1222 361898 36986 362134
rect 37222 361898 72986 362134
rect 73222 361898 108986 362134
rect 109222 361898 144986 362134
rect 145222 361898 180986 362134
rect 181222 361898 216986 362134
rect 217222 361898 252986 362134
rect 253222 361898 288986 362134
rect 289222 361898 324986 362134
rect 325222 361898 360986 362134
rect 361222 361898 396986 362134
rect 397222 361898 432986 362134
rect 433222 361898 468986 362134
rect 469222 361898 504986 362134
rect 505222 361898 540986 362134
rect 541222 361898 576986 362134
rect 577222 361898 585502 362134
rect 585738 361898 586840 362134
rect -2916 361876 586840 361898
rect -1996 361874 -1396 361876
rect 804 361874 1404 361876
rect 36804 361874 37404 361876
rect 72804 361874 73404 361876
rect 108804 361874 109404 361876
rect 144804 361874 145404 361876
rect 180804 361874 181404 361876
rect 216804 361874 217404 361876
rect 252804 361874 253404 361876
rect 288804 361874 289404 361876
rect 324804 361874 325404 361876
rect 360804 361874 361404 361876
rect 396804 361874 397404 361876
rect 432804 361874 433404 361876
rect 468804 361874 469404 361876
rect 504804 361874 505404 361876
rect 540804 361874 541404 361876
rect 576804 361874 577404 361876
rect 585320 361874 585920 361876
rect -8436 355276 -7836 355278
rect 29604 355276 30204 355278
rect 65604 355276 66204 355278
rect 101604 355276 102204 355278
rect 137604 355276 138204 355278
rect 173604 355276 174204 355278
rect 209604 355276 210204 355278
rect 245604 355276 246204 355278
rect 281604 355276 282204 355278
rect 317604 355276 318204 355278
rect 353604 355276 354204 355278
rect 389604 355276 390204 355278
rect 425604 355276 426204 355278
rect 461604 355276 462204 355278
rect 497604 355276 498204 355278
rect 533604 355276 534204 355278
rect 569604 355276 570204 355278
rect 591760 355276 592360 355278
rect -8436 355254 592360 355276
rect -8436 355018 -8254 355254
rect -8018 355018 29786 355254
rect 30022 355018 65786 355254
rect 66022 355018 101786 355254
rect 102022 355018 137786 355254
rect 138022 355018 173786 355254
rect 174022 355018 209786 355254
rect 210022 355018 245786 355254
rect 246022 355018 281786 355254
rect 282022 355018 317786 355254
rect 318022 355018 353786 355254
rect 354022 355018 389786 355254
rect 390022 355018 425786 355254
rect 426022 355018 461786 355254
rect 462022 355018 497786 355254
rect 498022 355018 533786 355254
rect 534022 355018 569786 355254
rect 570022 355018 591942 355254
rect 592178 355018 592360 355254
rect -8436 354934 592360 355018
rect -8436 354698 -8254 354934
rect -8018 354698 29786 354934
rect 30022 354698 65786 354934
rect 66022 354698 101786 354934
rect 102022 354698 137786 354934
rect 138022 354698 173786 354934
rect 174022 354698 209786 354934
rect 210022 354698 245786 354934
rect 246022 354698 281786 354934
rect 282022 354698 317786 354934
rect 318022 354698 353786 354934
rect 354022 354698 389786 354934
rect 390022 354698 425786 354934
rect 426022 354698 461786 354934
rect 462022 354698 497786 354934
rect 498022 354698 533786 354934
rect 534022 354698 569786 354934
rect 570022 354698 591942 354934
rect 592178 354698 592360 354934
rect -8436 354676 592360 354698
rect -8436 354674 -7836 354676
rect 29604 354674 30204 354676
rect 65604 354674 66204 354676
rect 101604 354674 102204 354676
rect 137604 354674 138204 354676
rect 173604 354674 174204 354676
rect 209604 354674 210204 354676
rect 245604 354674 246204 354676
rect 281604 354674 282204 354676
rect 317604 354674 318204 354676
rect 353604 354674 354204 354676
rect 389604 354674 390204 354676
rect 425604 354674 426204 354676
rect 461604 354674 462204 354676
rect 497604 354674 498204 354676
rect 533604 354674 534204 354676
rect 569604 354674 570204 354676
rect 591760 354674 592360 354676
rect -6596 351676 -5996 351678
rect 26004 351676 26604 351678
rect 62004 351676 62604 351678
rect 98004 351676 98604 351678
rect 134004 351676 134604 351678
rect 170004 351676 170604 351678
rect 206004 351676 206604 351678
rect 242004 351676 242604 351678
rect 278004 351676 278604 351678
rect 314004 351676 314604 351678
rect 350004 351676 350604 351678
rect 386004 351676 386604 351678
rect 422004 351676 422604 351678
rect 458004 351676 458604 351678
rect 494004 351676 494604 351678
rect 530004 351676 530604 351678
rect 566004 351676 566604 351678
rect 589920 351676 590520 351678
rect -6596 351654 590520 351676
rect -6596 351418 -6414 351654
rect -6178 351418 26186 351654
rect 26422 351418 62186 351654
rect 62422 351418 98186 351654
rect 98422 351418 134186 351654
rect 134422 351418 170186 351654
rect 170422 351418 206186 351654
rect 206422 351418 242186 351654
rect 242422 351418 278186 351654
rect 278422 351418 314186 351654
rect 314422 351418 350186 351654
rect 350422 351418 386186 351654
rect 386422 351418 422186 351654
rect 422422 351418 458186 351654
rect 458422 351418 494186 351654
rect 494422 351418 530186 351654
rect 530422 351418 566186 351654
rect 566422 351418 590102 351654
rect 590338 351418 590520 351654
rect -6596 351334 590520 351418
rect -6596 351098 -6414 351334
rect -6178 351098 26186 351334
rect 26422 351098 62186 351334
rect 62422 351098 98186 351334
rect 98422 351098 134186 351334
rect 134422 351098 170186 351334
rect 170422 351098 206186 351334
rect 206422 351098 242186 351334
rect 242422 351098 278186 351334
rect 278422 351098 314186 351334
rect 314422 351098 350186 351334
rect 350422 351098 386186 351334
rect 386422 351098 422186 351334
rect 422422 351098 458186 351334
rect 458422 351098 494186 351334
rect 494422 351098 530186 351334
rect 530422 351098 566186 351334
rect 566422 351098 590102 351334
rect 590338 351098 590520 351334
rect -6596 351076 590520 351098
rect -6596 351074 -5996 351076
rect 26004 351074 26604 351076
rect 62004 351074 62604 351076
rect 98004 351074 98604 351076
rect 134004 351074 134604 351076
rect 170004 351074 170604 351076
rect 206004 351074 206604 351076
rect 242004 351074 242604 351076
rect 278004 351074 278604 351076
rect 314004 351074 314604 351076
rect 350004 351074 350604 351076
rect 386004 351074 386604 351076
rect 422004 351074 422604 351076
rect 458004 351074 458604 351076
rect 494004 351074 494604 351076
rect 530004 351074 530604 351076
rect 566004 351074 566604 351076
rect 589920 351074 590520 351076
rect -4756 348076 -4156 348078
rect 22404 348076 23004 348078
rect 58404 348076 59004 348078
rect 94404 348076 95004 348078
rect 130404 348076 131004 348078
rect 166404 348076 167004 348078
rect 202404 348076 203004 348078
rect 238404 348076 239004 348078
rect 274404 348076 275004 348078
rect 310404 348076 311004 348078
rect 346404 348076 347004 348078
rect 382404 348076 383004 348078
rect 418404 348076 419004 348078
rect 454404 348076 455004 348078
rect 490404 348076 491004 348078
rect 526404 348076 527004 348078
rect 562404 348076 563004 348078
rect 588080 348076 588680 348078
rect -4756 348054 588680 348076
rect -4756 347818 -4574 348054
rect -4338 347818 22586 348054
rect 22822 347818 58586 348054
rect 58822 347818 94586 348054
rect 94822 347818 130586 348054
rect 130822 347818 166586 348054
rect 166822 347818 202586 348054
rect 202822 347818 238586 348054
rect 238822 347818 274586 348054
rect 274822 347818 310586 348054
rect 310822 347818 346586 348054
rect 346822 347818 382586 348054
rect 382822 347818 418586 348054
rect 418822 347818 454586 348054
rect 454822 347818 490586 348054
rect 490822 347818 526586 348054
rect 526822 347818 562586 348054
rect 562822 347818 588262 348054
rect 588498 347818 588680 348054
rect -4756 347734 588680 347818
rect -4756 347498 -4574 347734
rect -4338 347498 22586 347734
rect 22822 347498 58586 347734
rect 58822 347498 94586 347734
rect 94822 347498 130586 347734
rect 130822 347498 166586 347734
rect 166822 347498 202586 347734
rect 202822 347498 238586 347734
rect 238822 347498 274586 347734
rect 274822 347498 310586 347734
rect 310822 347498 346586 347734
rect 346822 347498 382586 347734
rect 382822 347498 418586 347734
rect 418822 347498 454586 347734
rect 454822 347498 490586 347734
rect 490822 347498 526586 347734
rect 526822 347498 562586 347734
rect 562822 347498 588262 347734
rect 588498 347498 588680 347734
rect -4756 347476 588680 347498
rect -4756 347474 -4156 347476
rect 22404 347474 23004 347476
rect 58404 347474 59004 347476
rect 94404 347474 95004 347476
rect 130404 347474 131004 347476
rect 166404 347474 167004 347476
rect 202404 347474 203004 347476
rect 238404 347474 239004 347476
rect 274404 347474 275004 347476
rect 310404 347474 311004 347476
rect 346404 347474 347004 347476
rect 382404 347474 383004 347476
rect 418404 347474 419004 347476
rect 454404 347474 455004 347476
rect 490404 347474 491004 347476
rect 526404 347474 527004 347476
rect 562404 347474 563004 347476
rect 588080 347474 588680 347476
rect -2916 344476 -2316 344478
rect 18804 344476 19404 344478
rect 54804 344476 55404 344478
rect 90804 344476 91404 344478
rect 126804 344476 127404 344478
rect 162804 344476 163404 344478
rect 198804 344476 199404 344478
rect 234804 344476 235404 344478
rect 270804 344476 271404 344478
rect 306804 344476 307404 344478
rect 342804 344476 343404 344478
rect 378804 344476 379404 344478
rect 414804 344476 415404 344478
rect 450804 344476 451404 344478
rect 486804 344476 487404 344478
rect 522804 344476 523404 344478
rect 558804 344476 559404 344478
rect 586240 344476 586840 344478
rect -2916 344454 586840 344476
rect -2916 344218 -2734 344454
rect -2498 344218 18986 344454
rect 19222 344218 54986 344454
rect 55222 344218 90986 344454
rect 91222 344218 126986 344454
rect 127222 344218 162986 344454
rect 163222 344218 198986 344454
rect 199222 344218 234986 344454
rect 235222 344218 270986 344454
rect 271222 344218 306986 344454
rect 307222 344218 342986 344454
rect 343222 344218 378986 344454
rect 379222 344218 414986 344454
rect 415222 344218 450986 344454
rect 451222 344218 486986 344454
rect 487222 344218 522986 344454
rect 523222 344218 558986 344454
rect 559222 344218 586422 344454
rect 586658 344218 586840 344454
rect -2916 344134 586840 344218
rect -2916 343898 -2734 344134
rect -2498 343898 18986 344134
rect 19222 343898 54986 344134
rect 55222 343898 90986 344134
rect 91222 343898 126986 344134
rect 127222 343898 162986 344134
rect 163222 343898 198986 344134
rect 199222 343898 234986 344134
rect 235222 343898 270986 344134
rect 271222 343898 306986 344134
rect 307222 343898 342986 344134
rect 343222 343898 378986 344134
rect 379222 343898 414986 344134
rect 415222 343898 450986 344134
rect 451222 343898 486986 344134
rect 487222 343898 522986 344134
rect 523222 343898 558986 344134
rect 559222 343898 586422 344134
rect 586658 343898 586840 344134
rect -2916 343876 586840 343898
rect -2916 343874 -2316 343876
rect 18804 343874 19404 343876
rect 54804 343874 55404 343876
rect 90804 343874 91404 343876
rect 126804 343874 127404 343876
rect 162804 343874 163404 343876
rect 198804 343874 199404 343876
rect 234804 343874 235404 343876
rect 270804 343874 271404 343876
rect 306804 343874 307404 343876
rect 342804 343874 343404 343876
rect 378804 343874 379404 343876
rect 414804 343874 415404 343876
rect 450804 343874 451404 343876
rect 486804 343874 487404 343876
rect 522804 343874 523404 343876
rect 558804 343874 559404 343876
rect 586240 343874 586840 343876
rect -7516 337276 -6916 337278
rect 11604 337276 12204 337278
rect 47604 337276 48204 337278
rect 83604 337276 84204 337278
rect 119604 337276 120204 337278
rect 155604 337276 156204 337278
rect 191604 337276 192204 337278
rect 227604 337276 228204 337278
rect 263604 337276 264204 337278
rect 299604 337276 300204 337278
rect 335604 337276 336204 337278
rect 371604 337276 372204 337278
rect 407604 337276 408204 337278
rect 443604 337276 444204 337278
rect 479604 337276 480204 337278
rect 515604 337276 516204 337278
rect 551604 337276 552204 337278
rect 590840 337276 591440 337278
rect -8436 337254 592360 337276
rect -8436 337018 -7334 337254
rect -7098 337018 11786 337254
rect 12022 337018 47786 337254
rect 48022 337018 83786 337254
rect 84022 337018 119786 337254
rect 120022 337018 155786 337254
rect 156022 337018 191786 337254
rect 192022 337018 227786 337254
rect 228022 337018 263786 337254
rect 264022 337018 299786 337254
rect 300022 337018 335786 337254
rect 336022 337018 371786 337254
rect 372022 337018 407786 337254
rect 408022 337018 443786 337254
rect 444022 337018 479786 337254
rect 480022 337018 515786 337254
rect 516022 337018 551786 337254
rect 552022 337018 591022 337254
rect 591258 337018 592360 337254
rect -8436 336934 592360 337018
rect -8436 336698 -7334 336934
rect -7098 336698 11786 336934
rect 12022 336698 47786 336934
rect 48022 336698 83786 336934
rect 84022 336698 119786 336934
rect 120022 336698 155786 336934
rect 156022 336698 191786 336934
rect 192022 336698 227786 336934
rect 228022 336698 263786 336934
rect 264022 336698 299786 336934
rect 300022 336698 335786 336934
rect 336022 336698 371786 336934
rect 372022 336698 407786 336934
rect 408022 336698 443786 336934
rect 444022 336698 479786 336934
rect 480022 336698 515786 336934
rect 516022 336698 551786 336934
rect 552022 336698 591022 336934
rect 591258 336698 592360 336934
rect -8436 336676 592360 336698
rect -7516 336674 -6916 336676
rect 11604 336674 12204 336676
rect 47604 336674 48204 336676
rect 83604 336674 84204 336676
rect 119604 336674 120204 336676
rect 155604 336674 156204 336676
rect 191604 336674 192204 336676
rect 227604 336674 228204 336676
rect 263604 336674 264204 336676
rect 299604 336674 300204 336676
rect 335604 336674 336204 336676
rect 371604 336674 372204 336676
rect 407604 336674 408204 336676
rect 443604 336674 444204 336676
rect 479604 336674 480204 336676
rect 515604 336674 516204 336676
rect 551604 336674 552204 336676
rect 590840 336674 591440 336676
rect -5676 333676 -5076 333678
rect 8004 333676 8604 333678
rect 44004 333676 44604 333678
rect 80004 333676 80604 333678
rect 116004 333676 116604 333678
rect 152004 333676 152604 333678
rect 188004 333676 188604 333678
rect 224004 333676 224604 333678
rect 260004 333676 260604 333678
rect 296004 333676 296604 333678
rect 332004 333676 332604 333678
rect 368004 333676 368604 333678
rect 404004 333676 404604 333678
rect 440004 333676 440604 333678
rect 476004 333676 476604 333678
rect 512004 333676 512604 333678
rect 548004 333676 548604 333678
rect 589000 333676 589600 333678
rect -6596 333654 590520 333676
rect -6596 333418 -5494 333654
rect -5258 333418 8186 333654
rect 8422 333418 44186 333654
rect 44422 333418 80186 333654
rect 80422 333418 116186 333654
rect 116422 333418 152186 333654
rect 152422 333418 188186 333654
rect 188422 333418 224186 333654
rect 224422 333418 260186 333654
rect 260422 333418 296186 333654
rect 296422 333418 332186 333654
rect 332422 333418 368186 333654
rect 368422 333418 404186 333654
rect 404422 333418 440186 333654
rect 440422 333418 476186 333654
rect 476422 333418 512186 333654
rect 512422 333418 548186 333654
rect 548422 333418 589182 333654
rect 589418 333418 590520 333654
rect -6596 333334 590520 333418
rect -6596 333098 -5494 333334
rect -5258 333098 8186 333334
rect 8422 333098 44186 333334
rect 44422 333098 80186 333334
rect 80422 333098 116186 333334
rect 116422 333098 152186 333334
rect 152422 333098 188186 333334
rect 188422 333098 224186 333334
rect 224422 333098 260186 333334
rect 260422 333098 296186 333334
rect 296422 333098 332186 333334
rect 332422 333098 368186 333334
rect 368422 333098 404186 333334
rect 404422 333098 440186 333334
rect 440422 333098 476186 333334
rect 476422 333098 512186 333334
rect 512422 333098 548186 333334
rect 548422 333098 589182 333334
rect 589418 333098 590520 333334
rect -6596 333076 590520 333098
rect -5676 333074 -5076 333076
rect 8004 333074 8604 333076
rect 44004 333074 44604 333076
rect 80004 333074 80604 333076
rect 116004 333074 116604 333076
rect 152004 333074 152604 333076
rect 188004 333074 188604 333076
rect 224004 333074 224604 333076
rect 260004 333074 260604 333076
rect 296004 333074 296604 333076
rect 332004 333074 332604 333076
rect 368004 333074 368604 333076
rect 404004 333074 404604 333076
rect 440004 333074 440604 333076
rect 476004 333074 476604 333076
rect 512004 333074 512604 333076
rect 548004 333074 548604 333076
rect 589000 333074 589600 333076
rect -3836 330076 -3236 330078
rect 4404 330076 5004 330078
rect 40404 330076 41004 330078
rect 76404 330076 77004 330078
rect 112404 330076 113004 330078
rect 148404 330076 149004 330078
rect 184404 330076 185004 330078
rect 220404 330076 221004 330078
rect 256404 330076 257004 330078
rect 292404 330076 293004 330078
rect 328404 330076 329004 330078
rect 364404 330076 365004 330078
rect 400404 330076 401004 330078
rect 436404 330076 437004 330078
rect 472404 330076 473004 330078
rect 508404 330076 509004 330078
rect 544404 330076 545004 330078
rect 580404 330076 581004 330078
rect 587160 330076 587760 330078
rect -4756 330054 588680 330076
rect -4756 329818 -3654 330054
rect -3418 329818 4586 330054
rect 4822 329818 40586 330054
rect 40822 329818 76586 330054
rect 76822 329818 112586 330054
rect 112822 329818 148586 330054
rect 148822 329818 184586 330054
rect 184822 329818 220586 330054
rect 220822 329818 256586 330054
rect 256822 329818 292586 330054
rect 292822 329818 328586 330054
rect 328822 329818 364586 330054
rect 364822 329818 400586 330054
rect 400822 329818 436586 330054
rect 436822 329818 472586 330054
rect 472822 329818 508586 330054
rect 508822 329818 544586 330054
rect 544822 329818 580586 330054
rect 580822 329818 587342 330054
rect 587578 329818 588680 330054
rect -4756 329734 588680 329818
rect -4756 329498 -3654 329734
rect -3418 329498 4586 329734
rect 4822 329498 40586 329734
rect 40822 329498 76586 329734
rect 76822 329498 112586 329734
rect 112822 329498 148586 329734
rect 148822 329498 184586 329734
rect 184822 329498 220586 329734
rect 220822 329498 256586 329734
rect 256822 329498 292586 329734
rect 292822 329498 328586 329734
rect 328822 329498 364586 329734
rect 364822 329498 400586 329734
rect 400822 329498 436586 329734
rect 436822 329498 472586 329734
rect 472822 329498 508586 329734
rect 508822 329498 544586 329734
rect 544822 329498 580586 329734
rect 580822 329498 587342 329734
rect 587578 329498 588680 329734
rect -4756 329476 588680 329498
rect -3836 329474 -3236 329476
rect 4404 329474 5004 329476
rect 40404 329474 41004 329476
rect 76404 329474 77004 329476
rect 112404 329474 113004 329476
rect 148404 329474 149004 329476
rect 184404 329474 185004 329476
rect 220404 329474 221004 329476
rect 256404 329474 257004 329476
rect 292404 329474 293004 329476
rect 328404 329474 329004 329476
rect 364404 329474 365004 329476
rect 400404 329474 401004 329476
rect 436404 329474 437004 329476
rect 472404 329474 473004 329476
rect 508404 329474 509004 329476
rect 544404 329474 545004 329476
rect 580404 329474 581004 329476
rect 587160 329474 587760 329476
rect -1996 326476 -1396 326478
rect 804 326476 1404 326478
rect 36804 326476 37404 326478
rect 72804 326476 73404 326478
rect 108804 326476 109404 326478
rect 144804 326476 145404 326478
rect 180804 326476 181404 326478
rect 216804 326476 217404 326478
rect 252804 326476 253404 326478
rect 288804 326476 289404 326478
rect 324804 326476 325404 326478
rect 360804 326476 361404 326478
rect 396804 326476 397404 326478
rect 432804 326476 433404 326478
rect 468804 326476 469404 326478
rect 504804 326476 505404 326478
rect 540804 326476 541404 326478
rect 576804 326476 577404 326478
rect 585320 326476 585920 326478
rect -2916 326454 586840 326476
rect -2916 326218 -1814 326454
rect -1578 326218 986 326454
rect 1222 326218 36986 326454
rect 37222 326218 72986 326454
rect 73222 326218 108986 326454
rect 109222 326218 144986 326454
rect 145222 326218 180986 326454
rect 181222 326218 216986 326454
rect 217222 326218 252986 326454
rect 253222 326218 288986 326454
rect 289222 326218 324986 326454
rect 325222 326218 360986 326454
rect 361222 326218 396986 326454
rect 397222 326218 432986 326454
rect 433222 326218 468986 326454
rect 469222 326218 504986 326454
rect 505222 326218 540986 326454
rect 541222 326218 576986 326454
rect 577222 326218 585502 326454
rect 585738 326218 586840 326454
rect -2916 326134 586840 326218
rect -2916 325898 -1814 326134
rect -1578 325898 986 326134
rect 1222 325898 36986 326134
rect 37222 325898 72986 326134
rect 73222 325898 108986 326134
rect 109222 325898 144986 326134
rect 145222 325898 180986 326134
rect 181222 325898 216986 326134
rect 217222 325898 252986 326134
rect 253222 325898 288986 326134
rect 289222 325898 324986 326134
rect 325222 325898 360986 326134
rect 361222 325898 396986 326134
rect 397222 325898 432986 326134
rect 433222 325898 468986 326134
rect 469222 325898 504986 326134
rect 505222 325898 540986 326134
rect 541222 325898 576986 326134
rect 577222 325898 585502 326134
rect 585738 325898 586840 326134
rect -2916 325876 586840 325898
rect -1996 325874 -1396 325876
rect 804 325874 1404 325876
rect 36804 325874 37404 325876
rect 72804 325874 73404 325876
rect 108804 325874 109404 325876
rect 144804 325874 145404 325876
rect 180804 325874 181404 325876
rect 216804 325874 217404 325876
rect 252804 325874 253404 325876
rect 288804 325874 289404 325876
rect 324804 325874 325404 325876
rect 360804 325874 361404 325876
rect 396804 325874 397404 325876
rect 432804 325874 433404 325876
rect 468804 325874 469404 325876
rect 504804 325874 505404 325876
rect 540804 325874 541404 325876
rect 576804 325874 577404 325876
rect 585320 325874 585920 325876
rect -8436 319276 -7836 319278
rect 29604 319276 30204 319278
rect 65604 319276 66204 319278
rect 101604 319276 102204 319278
rect 137604 319276 138204 319278
rect 173604 319276 174204 319278
rect 209604 319276 210204 319278
rect 245604 319276 246204 319278
rect 281604 319276 282204 319278
rect 317604 319276 318204 319278
rect 353604 319276 354204 319278
rect 389604 319276 390204 319278
rect 425604 319276 426204 319278
rect 461604 319276 462204 319278
rect 497604 319276 498204 319278
rect 533604 319276 534204 319278
rect 569604 319276 570204 319278
rect 591760 319276 592360 319278
rect -8436 319254 592360 319276
rect -8436 319018 -8254 319254
rect -8018 319018 29786 319254
rect 30022 319018 65786 319254
rect 66022 319018 101786 319254
rect 102022 319018 137786 319254
rect 138022 319018 173786 319254
rect 174022 319018 209786 319254
rect 210022 319018 245786 319254
rect 246022 319018 281786 319254
rect 282022 319018 317786 319254
rect 318022 319018 353786 319254
rect 354022 319018 389786 319254
rect 390022 319018 425786 319254
rect 426022 319018 461786 319254
rect 462022 319018 497786 319254
rect 498022 319018 533786 319254
rect 534022 319018 569786 319254
rect 570022 319018 591942 319254
rect 592178 319018 592360 319254
rect -8436 318934 592360 319018
rect -8436 318698 -8254 318934
rect -8018 318698 29786 318934
rect 30022 318698 65786 318934
rect 66022 318698 101786 318934
rect 102022 318698 137786 318934
rect 138022 318698 173786 318934
rect 174022 318698 209786 318934
rect 210022 318698 245786 318934
rect 246022 318698 281786 318934
rect 282022 318698 317786 318934
rect 318022 318698 353786 318934
rect 354022 318698 389786 318934
rect 390022 318698 425786 318934
rect 426022 318698 461786 318934
rect 462022 318698 497786 318934
rect 498022 318698 533786 318934
rect 534022 318698 569786 318934
rect 570022 318698 591942 318934
rect 592178 318698 592360 318934
rect -8436 318676 592360 318698
rect -8436 318674 -7836 318676
rect 29604 318674 30204 318676
rect 65604 318674 66204 318676
rect 101604 318674 102204 318676
rect 137604 318674 138204 318676
rect 173604 318674 174204 318676
rect 209604 318674 210204 318676
rect 245604 318674 246204 318676
rect 281604 318674 282204 318676
rect 317604 318674 318204 318676
rect 353604 318674 354204 318676
rect 389604 318674 390204 318676
rect 425604 318674 426204 318676
rect 461604 318674 462204 318676
rect 497604 318674 498204 318676
rect 533604 318674 534204 318676
rect 569604 318674 570204 318676
rect 591760 318674 592360 318676
rect -6596 315676 -5996 315678
rect 26004 315676 26604 315678
rect 62004 315676 62604 315678
rect 98004 315676 98604 315678
rect 134004 315676 134604 315678
rect 170004 315676 170604 315678
rect 206004 315676 206604 315678
rect 242004 315676 242604 315678
rect 278004 315676 278604 315678
rect 314004 315676 314604 315678
rect 350004 315676 350604 315678
rect 386004 315676 386604 315678
rect 422004 315676 422604 315678
rect 458004 315676 458604 315678
rect 494004 315676 494604 315678
rect 530004 315676 530604 315678
rect 566004 315676 566604 315678
rect 589920 315676 590520 315678
rect -6596 315654 590520 315676
rect -6596 315418 -6414 315654
rect -6178 315418 26186 315654
rect 26422 315418 62186 315654
rect 62422 315418 98186 315654
rect 98422 315418 134186 315654
rect 134422 315418 170186 315654
rect 170422 315418 206186 315654
rect 206422 315418 242186 315654
rect 242422 315418 278186 315654
rect 278422 315418 314186 315654
rect 314422 315418 350186 315654
rect 350422 315418 386186 315654
rect 386422 315418 422186 315654
rect 422422 315418 458186 315654
rect 458422 315418 494186 315654
rect 494422 315418 530186 315654
rect 530422 315418 566186 315654
rect 566422 315418 590102 315654
rect 590338 315418 590520 315654
rect -6596 315334 590520 315418
rect -6596 315098 -6414 315334
rect -6178 315098 26186 315334
rect 26422 315098 62186 315334
rect 62422 315098 98186 315334
rect 98422 315098 134186 315334
rect 134422 315098 170186 315334
rect 170422 315098 206186 315334
rect 206422 315098 242186 315334
rect 242422 315098 278186 315334
rect 278422 315098 314186 315334
rect 314422 315098 350186 315334
rect 350422 315098 386186 315334
rect 386422 315098 422186 315334
rect 422422 315098 458186 315334
rect 458422 315098 494186 315334
rect 494422 315098 530186 315334
rect 530422 315098 566186 315334
rect 566422 315098 590102 315334
rect 590338 315098 590520 315334
rect -6596 315076 590520 315098
rect -6596 315074 -5996 315076
rect 26004 315074 26604 315076
rect 62004 315074 62604 315076
rect 98004 315074 98604 315076
rect 134004 315074 134604 315076
rect 170004 315074 170604 315076
rect 206004 315074 206604 315076
rect 242004 315074 242604 315076
rect 278004 315074 278604 315076
rect 314004 315074 314604 315076
rect 350004 315074 350604 315076
rect 386004 315074 386604 315076
rect 422004 315074 422604 315076
rect 458004 315074 458604 315076
rect 494004 315074 494604 315076
rect 530004 315074 530604 315076
rect 566004 315074 566604 315076
rect 589920 315074 590520 315076
rect -4756 312076 -4156 312078
rect 22404 312076 23004 312078
rect 58404 312076 59004 312078
rect 94404 312076 95004 312078
rect 130404 312076 131004 312078
rect 166404 312076 167004 312078
rect 202404 312076 203004 312078
rect 238404 312076 239004 312078
rect 274404 312076 275004 312078
rect 310404 312076 311004 312078
rect 346404 312076 347004 312078
rect 382404 312076 383004 312078
rect 418404 312076 419004 312078
rect 454404 312076 455004 312078
rect 490404 312076 491004 312078
rect 526404 312076 527004 312078
rect 562404 312076 563004 312078
rect 588080 312076 588680 312078
rect -4756 312054 588680 312076
rect -4756 311818 -4574 312054
rect -4338 311818 22586 312054
rect 22822 311818 58586 312054
rect 58822 311818 94586 312054
rect 94822 311818 130586 312054
rect 130822 311818 166586 312054
rect 166822 311818 202586 312054
rect 202822 311818 238586 312054
rect 238822 311818 274586 312054
rect 274822 311818 310586 312054
rect 310822 311818 346586 312054
rect 346822 311818 382586 312054
rect 382822 311818 418586 312054
rect 418822 311818 454586 312054
rect 454822 311818 490586 312054
rect 490822 311818 526586 312054
rect 526822 311818 562586 312054
rect 562822 311818 588262 312054
rect 588498 311818 588680 312054
rect -4756 311734 588680 311818
rect -4756 311498 -4574 311734
rect -4338 311498 22586 311734
rect 22822 311498 58586 311734
rect 58822 311498 94586 311734
rect 94822 311498 130586 311734
rect 130822 311498 166586 311734
rect 166822 311498 202586 311734
rect 202822 311498 238586 311734
rect 238822 311498 274586 311734
rect 274822 311498 310586 311734
rect 310822 311498 346586 311734
rect 346822 311498 382586 311734
rect 382822 311498 418586 311734
rect 418822 311498 454586 311734
rect 454822 311498 490586 311734
rect 490822 311498 526586 311734
rect 526822 311498 562586 311734
rect 562822 311498 588262 311734
rect 588498 311498 588680 311734
rect -4756 311476 588680 311498
rect -4756 311474 -4156 311476
rect 22404 311474 23004 311476
rect 58404 311474 59004 311476
rect 94404 311474 95004 311476
rect 130404 311474 131004 311476
rect 166404 311474 167004 311476
rect 202404 311474 203004 311476
rect 238404 311474 239004 311476
rect 274404 311474 275004 311476
rect 310404 311474 311004 311476
rect 346404 311474 347004 311476
rect 382404 311474 383004 311476
rect 418404 311474 419004 311476
rect 454404 311474 455004 311476
rect 490404 311474 491004 311476
rect 526404 311474 527004 311476
rect 562404 311474 563004 311476
rect 588080 311474 588680 311476
rect -2916 308476 -2316 308478
rect 18804 308476 19404 308478
rect 54804 308476 55404 308478
rect 90804 308476 91404 308478
rect 126804 308476 127404 308478
rect 162804 308476 163404 308478
rect 198804 308476 199404 308478
rect 234804 308476 235404 308478
rect 270804 308476 271404 308478
rect 306804 308476 307404 308478
rect 342804 308476 343404 308478
rect 378804 308476 379404 308478
rect 414804 308476 415404 308478
rect 450804 308476 451404 308478
rect 486804 308476 487404 308478
rect 522804 308476 523404 308478
rect 558804 308476 559404 308478
rect 586240 308476 586840 308478
rect -2916 308454 586840 308476
rect -2916 308218 -2734 308454
rect -2498 308218 18986 308454
rect 19222 308218 54986 308454
rect 55222 308218 90986 308454
rect 91222 308218 126986 308454
rect 127222 308218 162986 308454
rect 163222 308218 198986 308454
rect 199222 308218 234986 308454
rect 235222 308218 270986 308454
rect 271222 308218 306986 308454
rect 307222 308218 342986 308454
rect 343222 308218 378986 308454
rect 379222 308218 414986 308454
rect 415222 308218 450986 308454
rect 451222 308218 486986 308454
rect 487222 308218 522986 308454
rect 523222 308218 558986 308454
rect 559222 308218 586422 308454
rect 586658 308218 586840 308454
rect -2916 308134 586840 308218
rect -2916 307898 -2734 308134
rect -2498 307898 18986 308134
rect 19222 307898 54986 308134
rect 55222 307898 90986 308134
rect 91222 307898 126986 308134
rect 127222 307898 162986 308134
rect 163222 307898 198986 308134
rect 199222 307898 234986 308134
rect 235222 307898 270986 308134
rect 271222 307898 306986 308134
rect 307222 307898 342986 308134
rect 343222 307898 378986 308134
rect 379222 307898 414986 308134
rect 415222 307898 450986 308134
rect 451222 307898 486986 308134
rect 487222 307898 522986 308134
rect 523222 307898 558986 308134
rect 559222 307898 586422 308134
rect 586658 307898 586840 308134
rect -2916 307876 586840 307898
rect -2916 307874 -2316 307876
rect 18804 307874 19404 307876
rect 54804 307874 55404 307876
rect 90804 307874 91404 307876
rect 126804 307874 127404 307876
rect 162804 307874 163404 307876
rect 198804 307874 199404 307876
rect 234804 307874 235404 307876
rect 270804 307874 271404 307876
rect 306804 307874 307404 307876
rect 342804 307874 343404 307876
rect 378804 307874 379404 307876
rect 414804 307874 415404 307876
rect 450804 307874 451404 307876
rect 486804 307874 487404 307876
rect 522804 307874 523404 307876
rect 558804 307874 559404 307876
rect 586240 307874 586840 307876
rect -7516 301276 -6916 301278
rect 11604 301276 12204 301278
rect 47604 301276 48204 301278
rect 83604 301276 84204 301278
rect 119604 301276 120204 301278
rect 155604 301276 156204 301278
rect 191604 301276 192204 301278
rect 227604 301276 228204 301278
rect 263604 301276 264204 301278
rect 299604 301276 300204 301278
rect 335604 301276 336204 301278
rect 371604 301276 372204 301278
rect 407604 301276 408204 301278
rect 443604 301276 444204 301278
rect 479604 301276 480204 301278
rect 515604 301276 516204 301278
rect 551604 301276 552204 301278
rect 590840 301276 591440 301278
rect -8436 301254 592360 301276
rect -8436 301018 -7334 301254
rect -7098 301018 11786 301254
rect 12022 301018 47786 301254
rect 48022 301018 83786 301254
rect 84022 301018 119786 301254
rect 120022 301018 155786 301254
rect 156022 301018 191786 301254
rect 192022 301018 227786 301254
rect 228022 301018 263786 301254
rect 264022 301018 299786 301254
rect 300022 301018 335786 301254
rect 336022 301018 371786 301254
rect 372022 301018 407786 301254
rect 408022 301018 443786 301254
rect 444022 301018 479786 301254
rect 480022 301018 515786 301254
rect 516022 301018 551786 301254
rect 552022 301018 591022 301254
rect 591258 301018 592360 301254
rect -8436 300934 592360 301018
rect -8436 300698 -7334 300934
rect -7098 300698 11786 300934
rect 12022 300698 47786 300934
rect 48022 300698 83786 300934
rect 84022 300698 119786 300934
rect 120022 300698 155786 300934
rect 156022 300698 191786 300934
rect 192022 300698 227786 300934
rect 228022 300698 263786 300934
rect 264022 300698 299786 300934
rect 300022 300698 335786 300934
rect 336022 300698 371786 300934
rect 372022 300698 407786 300934
rect 408022 300698 443786 300934
rect 444022 300698 479786 300934
rect 480022 300698 515786 300934
rect 516022 300698 551786 300934
rect 552022 300698 591022 300934
rect 591258 300698 592360 300934
rect -8436 300676 592360 300698
rect -7516 300674 -6916 300676
rect 11604 300674 12204 300676
rect 47604 300674 48204 300676
rect 83604 300674 84204 300676
rect 119604 300674 120204 300676
rect 155604 300674 156204 300676
rect 191604 300674 192204 300676
rect 227604 300674 228204 300676
rect 263604 300674 264204 300676
rect 299604 300674 300204 300676
rect 335604 300674 336204 300676
rect 371604 300674 372204 300676
rect 407604 300674 408204 300676
rect 443604 300674 444204 300676
rect 479604 300674 480204 300676
rect 515604 300674 516204 300676
rect 551604 300674 552204 300676
rect 590840 300674 591440 300676
rect -5676 297676 -5076 297678
rect 8004 297676 8604 297678
rect 44004 297676 44604 297678
rect 80004 297676 80604 297678
rect 116004 297676 116604 297678
rect 152004 297676 152604 297678
rect 188004 297676 188604 297678
rect 224004 297676 224604 297678
rect 260004 297676 260604 297678
rect 296004 297676 296604 297678
rect 332004 297676 332604 297678
rect 368004 297676 368604 297678
rect 404004 297676 404604 297678
rect 440004 297676 440604 297678
rect 476004 297676 476604 297678
rect 512004 297676 512604 297678
rect 548004 297676 548604 297678
rect 589000 297676 589600 297678
rect -6596 297654 590520 297676
rect -6596 297418 -5494 297654
rect -5258 297418 8186 297654
rect 8422 297418 44186 297654
rect 44422 297418 80186 297654
rect 80422 297418 116186 297654
rect 116422 297418 152186 297654
rect 152422 297418 188186 297654
rect 188422 297418 224186 297654
rect 224422 297418 260186 297654
rect 260422 297418 296186 297654
rect 296422 297418 332186 297654
rect 332422 297418 368186 297654
rect 368422 297418 404186 297654
rect 404422 297418 440186 297654
rect 440422 297418 476186 297654
rect 476422 297418 512186 297654
rect 512422 297418 548186 297654
rect 548422 297418 589182 297654
rect 589418 297418 590520 297654
rect -6596 297334 590520 297418
rect -6596 297098 -5494 297334
rect -5258 297098 8186 297334
rect 8422 297098 44186 297334
rect 44422 297098 80186 297334
rect 80422 297098 116186 297334
rect 116422 297098 152186 297334
rect 152422 297098 188186 297334
rect 188422 297098 224186 297334
rect 224422 297098 260186 297334
rect 260422 297098 296186 297334
rect 296422 297098 332186 297334
rect 332422 297098 368186 297334
rect 368422 297098 404186 297334
rect 404422 297098 440186 297334
rect 440422 297098 476186 297334
rect 476422 297098 512186 297334
rect 512422 297098 548186 297334
rect 548422 297098 589182 297334
rect 589418 297098 590520 297334
rect -6596 297076 590520 297098
rect -5676 297074 -5076 297076
rect 8004 297074 8604 297076
rect 44004 297074 44604 297076
rect 80004 297074 80604 297076
rect 116004 297074 116604 297076
rect 152004 297074 152604 297076
rect 188004 297074 188604 297076
rect 224004 297074 224604 297076
rect 260004 297074 260604 297076
rect 296004 297074 296604 297076
rect 332004 297074 332604 297076
rect 368004 297074 368604 297076
rect 404004 297074 404604 297076
rect 440004 297074 440604 297076
rect 476004 297074 476604 297076
rect 512004 297074 512604 297076
rect 548004 297074 548604 297076
rect 589000 297074 589600 297076
rect -3836 294076 -3236 294078
rect 4404 294076 5004 294078
rect 40404 294076 41004 294078
rect 76404 294076 77004 294078
rect 112404 294076 113004 294078
rect 148404 294076 149004 294078
rect 184404 294076 185004 294078
rect 220404 294076 221004 294078
rect 256404 294076 257004 294078
rect 292404 294076 293004 294078
rect 328404 294076 329004 294078
rect 364404 294076 365004 294078
rect 400404 294076 401004 294078
rect 436404 294076 437004 294078
rect 472404 294076 473004 294078
rect 508404 294076 509004 294078
rect 544404 294076 545004 294078
rect 580404 294076 581004 294078
rect 587160 294076 587760 294078
rect -4756 294054 588680 294076
rect -4756 293818 -3654 294054
rect -3418 293818 4586 294054
rect 4822 293818 40586 294054
rect 40822 293818 76586 294054
rect 76822 293818 112586 294054
rect 112822 293818 148586 294054
rect 148822 293818 184586 294054
rect 184822 293818 220586 294054
rect 220822 293818 256586 294054
rect 256822 293818 292586 294054
rect 292822 293818 328586 294054
rect 328822 293818 364586 294054
rect 364822 293818 400586 294054
rect 400822 293818 436586 294054
rect 436822 293818 472586 294054
rect 472822 293818 508586 294054
rect 508822 293818 544586 294054
rect 544822 293818 580586 294054
rect 580822 293818 587342 294054
rect 587578 293818 588680 294054
rect -4756 293734 588680 293818
rect -4756 293498 -3654 293734
rect -3418 293498 4586 293734
rect 4822 293498 40586 293734
rect 40822 293498 76586 293734
rect 76822 293498 112586 293734
rect 112822 293498 148586 293734
rect 148822 293498 184586 293734
rect 184822 293498 220586 293734
rect 220822 293498 256586 293734
rect 256822 293498 292586 293734
rect 292822 293498 328586 293734
rect 328822 293498 364586 293734
rect 364822 293498 400586 293734
rect 400822 293498 436586 293734
rect 436822 293498 472586 293734
rect 472822 293498 508586 293734
rect 508822 293498 544586 293734
rect 544822 293498 580586 293734
rect 580822 293498 587342 293734
rect 587578 293498 588680 293734
rect -4756 293476 588680 293498
rect -3836 293474 -3236 293476
rect 4404 293474 5004 293476
rect 40404 293474 41004 293476
rect 76404 293474 77004 293476
rect 112404 293474 113004 293476
rect 148404 293474 149004 293476
rect 184404 293474 185004 293476
rect 220404 293474 221004 293476
rect 256404 293474 257004 293476
rect 292404 293474 293004 293476
rect 328404 293474 329004 293476
rect 364404 293474 365004 293476
rect 400404 293474 401004 293476
rect 436404 293474 437004 293476
rect 472404 293474 473004 293476
rect 508404 293474 509004 293476
rect 544404 293474 545004 293476
rect 580404 293474 581004 293476
rect 587160 293474 587760 293476
rect -1996 290476 -1396 290478
rect 804 290476 1404 290478
rect 36804 290476 37404 290478
rect 72804 290476 73404 290478
rect 108804 290476 109404 290478
rect 144804 290476 145404 290478
rect 180804 290476 181404 290478
rect 216804 290476 217404 290478
rect 252804 290476 253404 290478
rect 288804 290476 289404 290478
rect 324804 290476 325404 290478
rect 360804 290476 361404 290478
rect 396804 290476 397404 290478
rect 432804 290476 433404 290478
rect 468804 290476 469404 290478
rect 504804 290476 505404 290478
rect 540804 290476 541404 290478
rect 576804 290476 577404 290478
rect 585320 290476 585920 290478
rect -2916 290454 586840 290476
rect -2916 290218 -1814 290454
rect -1578 290218 986 290454
rect 1222 290218 36986 290454
rect 37222 290218 72986 290454
rect 73222 290218 108986 290454
rect 109222 290218 144986 290454
rect 145222 290218 180986 290454
rect 181222 290218 216986 290454
rect 217222 290218 252986 290454
rect 253222 290218 288986 290454
rect 289222 290218 324986 290454
rect 325222 290218 360986 290454
rect 361222 290218 396986 290454
rect 397222 290218 432986 290454
rect 433222 290218 468986 290454
rect 469222 290218 504986 290454
rect 505222 290218 540986 290454
rect 541222 290218 576986 290454
rect 577222 290218 585502 290454
rect 585738 290218 586840 290454
rect -2916 290134 586840 290218
rect -2916 289898 -1814 290134
rect -1578 289898 986 290134
rect 1222 289898 36986 290134
rect 37222 289898 72986 290134
rect 73222 289898 108986 290134
rect 109222 289898 144986 290134
rect 145222 289898 180986 290134
rect 181222 289898 216986 290134
rect 217222 289898 252986 290134
rect 253222 289898 288986 290134
rect 289222 289898 324986 290134
rect 325222 289898 360986 290134
rect 361222 289898 396986 290134
rect 397222 289898 432986 290134
rect 433222 289898 468986 290134
rect 469222 289898 504986 290134
rect 505222 289898 540986 290134
rect 541222 289898 576986 290134
rect 577222 289898 585502 290134
rect 585738 289898 586840 290134
rect -2916 289876 586840 289898
rect -1996 289874 -1396 289876
rect 804 289874 1404 289876
rect 36804 289874 37404 289876
rect 72804 289874 73404 289876
rect 108804 289874 109404 289876
rect 144804 289874 145404 289876
rect 180804 289874 181404 289876
rect 216804 289874 217404 289876
rect 252804 289874 253404 289876
rect 288804 289874 289404 289876
rect 324804 289874 325404 289876
rect 360804 289874 361404 289876
rect 396804 289874 397404 289876
rect 432804 289874 433404 289876
rect 468804 289874 469404 289876
rect 504804 289874 505404 289876
rect 540804 289874 541404 289876
rect 576804 289874 577404 289876
rect 585320 289874 585920 289876
rect -8436 283276 -7836 283278
rect 29604 283276 30204 283278
rect 65604 283276 66204 283278
rect 101604 283276 102204 283278
rect 137604 283276 138204 283278
rect 173604 283276 174204 283278
rect 209604 283276 210204 283278
rect 245604 283276 246204 283278
rect 281604 283276 282204 283278
rect 317604 283276 318204 283278
rect 353604 283276 354204 283278
rect 389604 283276 390204 283278
rect 425604 283276 426204 283278
rect 461604 283276 462204 283278
rect 497604 283276 498204 283278
rect 533604 283276 534204 283278
rect 569604 283276 570204 283278
rect 591760 283276 592360 283278
rect -8436 283254 592360 283276
rect -8436 283018 -8254 283254
rect -8018 283018 29786 283254
rect 30022 283018 65786 283254
rect 66022 283018 101786 283254
rect 102022 283018 137786 283254
rect 138022 283018 173786 283254
rect 174022 283018 209786 283254
rect 210022 283018 245786 283254
rect 246022 283018 281786 283254
rect 282022 283018 317786 283254
rect 318022 283018 353786 283254
rect 354022 283018 389786 283254
rect 390022 283018 425786 283254
rect 426022 283018 461786 283254
rect 462022 283018 497786 283254
rect 498022 283018 533786 283254
rect 534022 283018 569786 283254
rect 570022 283018 591942 283254
rect 592178 283018 592360 283254
rect -8436 282934 592360 283018
rect -8436 282698 -8254 282934
rect -8018 282698 29786 282934
rect 30022 282698 65786 282934
rect 66022 282698 101786 282934
rect 102022 282698 137786 282934
rect 138022 282698 173786 282934
rect 174022 282698 209786 282934
rect 210022 282698 245786 282934
rect 246022 282698 281786 282934
rect 282022 282698 317786 282934
rect 318022 282698 353786 282934
rect 354022 282698 389786 282934
rect 390022 282698 425786 282934
rect 426022 282698 461786 282934
rect 462022 282698 497786 282934
rect 498022 282698 533786 282934
rect 534022 282698 569786 282934
rect 570022 282698 591942 282934
rect 592178 282698 592360 282934
rect -8436 282676 592360 282698
rect -8436 282674 -7836 282676
rect 29604 282674 30204 282676
rect 65604 282674 66204 282676
rect 101604 282674 102204 282676
rect 137604 282674 138204 282676
rect 173604 282674 174204 282676
rect 209604 282674 210204 282676
rect 245604 282674 246204 282676
rect 281604 282674 282204 282676
rect 317604 282674 318204 282676
rect 353604 282674 354204 282676
rect 389604 282674 390204 282676
rect 425604 282674 426204 282676
rect 461604 282674 462204 282676
rect 497604 282674 498204 282676
rect 533604 282674 534204 282676
rect 569604 282674 570204 282676
rect 591760 282674 592360 282676
rect -6596 279676 -5996 279678
rect 26004 279676 26604 279678
rect 62004 279676 62604 279678
rect 98004 279676 98604 279678
rect 134004 279676 134604 279678
rect 170004 279676 170604 279678
rect 206004 279676 206604 279678
rect 242004 279676 242604 279678
rect 278004 279676 278604 279678
rect 314004 279676 314604 279678
rect 350004 279676 350604 279678
rect 386004 279676 386604 279678
rect 422004 279676 422604 279678
rect 458004 279676 458604 279678
rect 494004 279676 494604 279678
rect 530004 279676 530604 279678
rect 566004 279676 566604 279678
rect 589920 279676 590520 279678
rect -6596 279654 590520 279676
rect -6596 279418 -6414 279654
rect -6178 279418 26186 279654
rect 26422 279418 62186 279654
rect 62422 279418 98186 279654
rect 98422 279418 134186 279654
rect 134422 279418 170186 279654
rect 170422 279418 206186 279654
rect 206422 279418 242186 279654
rect 242422 279418 278186 279654
rect 278422 279418 314186 279654
rect 314422 279418 350186 279654
rect 350422 279418 386186 279654
rect 386422 279418 422186 279654
rect 422422 279418 458186 279654
rect 458422 279418 494186 279654
rect 494422 279418 530186 279654
rect 530422 279418 566186 279654
rect 566422 279418 590102 279654
rect 590338 279418 590520 279654
rect -6596 279334 590520 279418
rect -6596 279098 -6414 279334
rect -6178 279098 26186 279334
rect 26422 279098 62186 279334
rect 62422 279098 98186 279334
rect 98422 279098 134186 279334
rect 134422 279098 170186 279334
rect 170422 279098 206186 279334
rect 206422 279098 242186 279334
rect 242422 279098 278186 279334
rect 278422 279098 314186 279334
rect 314422 279098 350186 279334
rect 350422 279098 386186 279334
rect 386422 279098 422186 279334
rect 422422 279098 458186 279334
rect 458422 279098 494186 279334
rect 494422 279098 530186 279334
rect 530422 279098 566186 279334
rect 566422 279098 590102 279334
rect 590338 279098 590520 279334
rect -6596 279076 590520 279098
rect -6596 279074 -5996 279076
rect 26004 279074 26604 279076
rect 62004 279074 62604 279076
rect 98004 279074 98604 279076
rect 134004 279074 134604 279076
rect 170004 279074 170604 279076
rect 206004 279074 206604 279076
rect 242004 279074 242604 279076
rect 278004 279074 278604 279076
rect 314004 279074 314604 279076
rect 350004 279074 350604 279076
rect 386004 279074 386604 279076
rect 422004 279074 422604 279076
rect 458004 279074 458604 279076
rect 494004 279074 494604 279076
rect 530004 279074 530604 279076
rect 566004 279074 566604 279076
rect 589920 279074 590520 279076
rect -4756 276076 -4156 276078
rect 22404 276076 23004 276078
rect 58404 276076 59004 276078
rect 94404 276076 95004 276078
rect 130404 276076 131004 276078
rect 166404 276076 167004 276078
rect 202404 276076 203004 276078
rect 238404 276076 239004 276078
rect 274404 276076 275004 276078
rect 310404 276076 311004 276078
rect 346404 276076 347004 276078
rect 382404 276076 383004 276078
rect 418404 276076 419004 276078
rect 454404 276076 455004 276078
rect 490404 276076 491004 276078
rect 526404 276076 527004 276078
rect 562404 276076 563004 276078
rect 588080 276076 588680 276078
rect -4756 276054 588680 276076
rect -4756 275818 -4574 276054
rect -4338 275818 22586 276054
rect 22822 275818 58586 276054
rect 58822 275818 94586 276054
rect 94822 275818 130586 276054
rect 130822 275818 166586 276054
rect 166822 275818 202586 276054
rect 202822 275818 238586 276054
rect 238822 275818 274586 276054
rect 274822 275818 310586 276054
rect 310822 275818 346586 276054
rect 346822 275818 382586 276054
rect 382822 275818 418586 276054
rect 418822 275818 454586 276054
rect 454822 275818 490586 276054
rect 490822 275818 526586 276054
rect 526822 275818 562586 276054
rect 562822 275818 588262 276054
rect 588498 275818 588680 276054
rect -4756 275734 588680 275818
rect -4756 275498 -4574 275734
rect -4338 275498 22586 275734
rect 22822 275498 58586 275734
rect 58822 275498 94586 275734
rect 94822 275498 130586 275734
rect 130822 275498 166586 275734
rect 166822 275498 202586 275734
rect 202822 275498 238586 275734
rect 238822 275498 274586 275734
rect 274822 275498 310586 275734
rect 310822 275498 346586 275734
rect 346822 275498 382586 275734
rect 382822 275498 418586 275734
rect 418822 275498 454586 275734
rect 454822 275498 490586 275734
rect 490822 275498 526586 275734
rect 526822 275498 562586 275734
rect 562822 275498 588262 275734
rect 588498 275498 588680 275734
rect -4756 275476 588680 275498
rect -4756 275474 -4156 275476
rect 22404 275474 23004 275476
rect 58404 275474 59004 275476
rect 94404 275474 95004 275476
rect 130404 275474 131004 275476
rect 166404 275474 167004 275476
rect 202404 275474 203004 275476
rect 238404 275474 239004 275476
rect 274404 275474 275004 275476
rect 310404 275474 311004 275476
rect 346404 275474 347004 275476
rect 382404 275474 383004 275476
rect 418404 275474 419004 275476
rect 454404 275474 455004 275476
rect 490404 275474 491004 275476
rect 526404 275474 527004 275476
rect 562404 275474 563004 275476
rect 588080 275474 588680 275476
rect -2916 272476 -2316 272478
rect 18804 272476 19404 272478
rect 54804 272476 55404 272478
rect 90804 272476 91404 272478
rect 126804 272476 127404 272478
rect 162804 272476 163404 272478
rect 198804 272476 199404 272478
rect 234804 272476 235404 272478
rect 270804 272476 271404 272478
rect 306804 272476 307404 272478
rect 342804 272476 343404 272478
rect 378804 272476 379404 272478
rect 414804 272476 415404 272478
rect 450804 272476 451404 272478
rect 486804 272476 487404 272478
rect 522804 272476 523404 272478
rect 558804 272476 559404 272478
rect 586240 272476 586840 272478
rect -2916 272454 586840 272476
rect -2916 272218 -2734 272454
rect -2498 272218 18986 272454
rect 19222 272218 54986 272454
rect 55222 272218 90986 272454
rect 91222 272218 126986 272454
rect 127222 272218 162986 272454
rect 163222 272218 198986 272454
rect 199222 272218 234986 272454
rect 235222 272218 270986 272454
rect 271222 272218 306986 272454
rect 307222 272218 342986 272454
rect 343222 272218 378986 272454
rect 379222 272218 414986 272454
rect 415222 272218 450986 272454
rect 451222 272218 486986 272454
rect 487222 272218 522986 272454
rect 523222 272218 558986 272454
rect 559222 272218 586422 272454
rect 586658 272218 586840 272454
rect -2916 272134 586840 272218
rect -2916 271898 -2734 272134
rect -2498 271898 18986 272134
rect 19222 271898 54986 272134
rect 55222 271898 90986 272134
rect 91222 271898 126986 272134
rect 127222 271898 162986 272134
rect 163222 271898 198986 272134
rect 199222 271898 234986 272134
rect 235222 271898 270986 272134
rect 271222 271898 306986 272134
rect 307222 271898 342986 272134
rect 343222 271898 378986 272134
rect 379222 271898 414986 272134
rect 415222 271898 450986 272134
rect 451222 271898 486986 272134
rect 487222 271898 522986 272134
rect 523222 271898 558986 272134
rect 559222 271898 586422 272134
rect 586658 271898 586840 272134
rect -2916 271876 586840 271898
rect -2916 271874 -2316 271876
rect 18804 271874 19404 271876
rect 54804 271874 55404 271876
rect 90804 271874 91404 271876
rect 126804 271874 127404 271876
rect 162804 271874 163404 271876
rect 198804 271874 199404 271876
rect 234804 271874 235404 271876
rect 270804 271874 271404 271876
rect 306804 271874 307404 271876
rect 342804 271874 343404 271876
rect 378804 271874 379404 271876
rect 414804 271874 415404 271876
rect 450804 271874 451404 271876
rect 486804 271874 487404 271876
rect 522804 271874 523404 271876
rect 558804 271874 559404 271876
rect 586240 271874 586840 271876
rect -7516 265276 -6916 265278
rect 11604 265276 12204 265278
rect 47604 265276 48204 265278
rect 83604 265276 84204 265278
rect 119604 265276 120204 265278
rect 155604 265276 156204 265278
rect 191604 265276 192204 265278
rect 227604 265276 228204 265278
rect 263604 265276 264204 265278
rect 299604 265276 300204 265278
rect 335604 265276 336204 265278
rect 371604 265276 372204 265278
rect 407604 265276 408204 265278
rect 443604 265276 444204 265278
rect 479604 265276 480204 265278
rect 515604 265276 516204 265278
rect 551604 265276 552204 265278
rect 590840 265276 591440 265278
rect -8436 265254 592360 265276
rect -8436 265018 -7334 265254
rect -7098 265018 11786 265254
rect 12022 265018 47786 265254
rect 48022 265018 83786 265254
rect 84022 265018 119786 265254
rect 120022 265018 155786 265254
rect 156022 265018 191786 265254
rect 192022 265018 227786 265254
rect 228022 265018 263786 265254
rect 264022 265018 299786 265254
rect 300022 265018 335786 265254
rect 336022 265018 371786 265254
rect 372022 265018 407786 265254
rect 408022 265018 443786 265254
rect 444022 265018 479786 265254
rect 480022 265018 515786 265254
rect 516022 265018 551786 265254
rect 552022 265018 591022 265254
rect 591258 265018 592360 265254
rect -8436 264934 592360 265018
rect -8436 264698 -7334 264934
rect -7098 264698 11786 264934
rect 12022 264698 47786 264934
rect 48022 264698 83786 264934
rect 84022 264698 119786 264934
rect 120022 264698 155786 264934
rect 156022 264698 191786 264934
rect 192022 264698 227786 264934
rect 228022 264698 263786 264934
rect 264022 264698 299786 264934
rect 300022 264698 335786 264934
rect 336022 264698 371786 264934
rect 372022 264698 407786 264934
rect 408022 264698 443786 264934
rect 444022 264698 479786 264934
rect 480022 264698 515786 264934
rect 516022 264698 551786 264934
rect 552022 264698 591022 264934
rect 591258 264698 592360 264934
rect -8436 264676 592360 264698
rect -7516 264674 -6916 264676
rect 11604 264674 12204 264676
rect 47604 264674 48204 264676
rect 83604 264674 84204 264676
rect 119604 264674 120204 264676
rect 155604 264674 156204 264676
rect 191604 264674 192204 264676
rect 227604 264674 228204 264676
rect 263604 264674 264204 264676
rect 299604 264674 300204 264676
rect 335604 264674 336204 264676
rect 371604 264674 372204 264676
rect 407604 264674 408204 264676
rect 443604 264674 444204 264676
rect 479604 264674 480204 264676
rect 515604 264674 516204 264676
rect 551604 264674 552204 264676
rect 590840 264674 591440 264676
rect -5676 261676 -5076 261678
rect 8004 261676 8604 261678
rect 44004 261676 44604 261678
rect 80004 261676 80604 261678
rect 116004 261676 116604 261678
rect 152004 261676 152604 261678
rect 188004 261676 188604 261678
rect 224004 261676 224604 261678
rect 260004 261676 260604 261678
rect 296004 261676 296604 261678
rect 332004 261676 332604 261678
rect 368004 261676 368604 261678
rect 404004 261676 404604 261678
rect 440004 261676 440604 261678
rect 476004 261676 476604 261678
rect 512004 261676 512604 261678
rect 548004 261676 548604 261678
rect 589000 261676 589600 261678
rect -6596 261654 590520 261676
rect -6596 261418 -5494 261654
rect -5258 261418 8186 261654
rect 8422 261418 44186 261654
rect 44422 261418 80186 261654
rect 80422 261418 116186 261654
rect 116422 261418 152186 261654
rect 152422 261418 188186 261654
rect 188422 261418 224186 261654
rect 224422 261418 260186 261654
rect 260422 261418 296186 261654
rect 296422 261418 332186 261654
rect 332422 261418 368186 261654
rect 368422 261418 404186 261654
rect 404422 261418 440186 261654
rect 440422 261418 476186 261654
rect 476422 261418 512186 261654
rect 512422 261418 548186 261654
rect 548422 261418 589182 261654
rect 589418 261418 590520 261654
rect -6596 261334 590520 261418
rect -6596 261098 -5494 261334
rect -5258 261098 8186 261334
rect 8422 261098 44186 261334
rect 44422 261098 80186 261334
rect 80422 261098 116186 261334
rect 116422 261098 152186 261334
rect 152422 261098 188186 261334
rect 188422 261098 224186 261334
rect 224422 261098 260186 261334
rect 260422 261098 296186 261334
rect 296422 261098 332186 261334
rect 332422 261098 368186 261334
rect 368422 261098 404186 261334
rect 404422 261098 440186 261334
rect 440422 261098 476186 261334
rect 476422 261098 512186 261334
rect 512422 261098 548186 261334
rect 548422 261098 589182 261334
rect 589418 261098 590520 261334
rect -6596 261076 590520 261098
rect -5676 261074 -5076 261076
rect 8004 261074 8604 261076
rect 44004 261074 44604 261076
rect 80004 261074 80604 261076
rect 116004 261074 116604 261076
rect 152004 261074 152604 261076
rect 188004 261074 188604 261076
rect 224004 261074 224604 261076
rect 260004 261074 260604 261076
rect 296004 261074 296604 261076
rect 332004 261074 332604 261076
rect 368004 261074 368604 261076
rect 404004 261074 404604 261076
rect 440004 261074 440604 261076
rect 476004 261074 476604 261076
rect 512004 261074 512604 261076
rect 548004 261074 548604 261076
rect 589000 261074 589600 261076
rect -3836 258076 -3236 258078
rect 4404 258076 5004 258078
rect 40404 258076 41004 258078
rect 76404 258076 77004 258078
rect 112404 258076 113004 258078
rect 148404 258076 149004 258078
rect 184404 258076 185004 258078
rect 220404 258076 221004 258078
rect 256404 258076 257004 258078
rect 292404 258076 293004 258078
rect 328404 258076 329004 258078
rect 364404 258076 365004 258078
rect 400404 258076 401004 258078
rect 436404 258076 437004 258078
rect 472404 258076 473004 258078
rect 508404 258076 509004 258078
rect 544404 258076 545004 258078
rect 580404 258076 581004 258078
rect 587160 258076 587760 258078
rect -4756 258054 588680 258076
rect -4756 257818 -3654 258054
rect -3418 257818 4586 258054
rect 4822 257818 40586 258054
rect 40822 257818 76586 258054
rect 76822 257818 112586 258054
rect 112822 257818 148586 258054
rect 148822 257818 184586 258054
rect 184822 257818 220586 258054
rect 220822 257818 256586 258054
rect 256822 257818 292586 258054
rect 292822 257818 328586 258054
rect 328822 257818 364586 258054
rect 364822 257818 400586 258054
rect 400822 257818 436586 258054
rect 436822 257818 472586 258054
rect 472822 257818 508586 258054
rect 508822 257818 544586 258054
rect 544822 257818 580586 258054
rect 580822 257818 587342 258054
rect 587578 257818 588680 258054
rect -4756 257734 588680 257818
rect -4756 257498 -3654 257734
rect -3418 257498 4586 257734
rect 4822 257498 40586 257734
rect 40822 257498 76586 257734
rect 76822 257498 112586 257734
rect 112822 257498 148586 257734
rect 148822 257498 184586 257734
rect 184822 257498 220586 257734
rect 220822 257498 256586 257734
rect 256822 257498 292586 257734
rect 292822 257498 328586 257734
rect 328822 257498 364586 257734
rect 364822 257498 400586 257734
rect 400822 257498 436586 257734
rect 436822 257498 472586 257734
rect 472822 257498 508586 257734
rect 508822 257498 544586 257734
rect 544822 257498 580586 257734
rect 580822 257498 587342 257734
rect 587578 257498 588680 257734
rect -4756 257476 588680 257498
rect -3836 257474 -3236 257476
rect 4404 257474 5004 257476
rect 40404 257474 41004 257476
rect 76404 257474 77004 257476
rect 112404 257474 113004 257476
rect 148404 257474 149004 257476
rect 184404 257474 185004 257476
rect 220404 257474 221004 257476
rect 256404 257474 257004 257476
rect 292404 257474 293004 257476
rect 328404 257474 329004 257476
rect 364404 257474 365004 257476
rect 400404 257474 401004 257476
rect 436404 257474 437004 257476
rect 472404 257474 473004 257476
rect 508404 257474 509004 257476
rect 544404 257474 545004 257476
rect 580404 257474 581004 257476
rect 587160 257474 587760 257476
rect -1996 254476 -1396 254478
rect 804 254476 1404 254478
rect 36804 254476 37404 254478
rect 72804 254476 73404 254478
rect 108804 254476 109404 254478
rect 144804 254476 145404 254478
rect 180804 254476 181404 254478
rect 216804 254476 217404 254478
rect 252804 254476 253404 254478
rect 288804 254476 289404 254478
rect 324804 254476 325404 254478
rect 360804 254476 361404 254478
rect 396804 254476 397404 254478
rect 432804 254476 433404 254478
rect 468804 254476 469404 254478
rect 504804 254476 505404 254478
rect 540804 254476 541404 254478
rect 576804 254476 577404 254478
rect 585320 254476 585920 254478
rect -2916 254454 586840 254476
rect -2916 254218 -1814 254454
rect -1578 254218 986 254454
rect 1222 254218 36986 254454
rect 37222 254218 72986 254454
rect 73222 254218 108986 254454
rect 109222 254218 144986 254454
rect 145222 254218 180986 254454
rect 181222 254218 216986 254454
rect 217222 254218 252986 254454
rect 253222 254218 288986 254454
rect 289222 254218 324986 254454
rect 325222 254218 360986 254454
rect 361222 254218 396986 254454
rect 397222 254218 432986 254454
rect 433222 254218 468986 254454
rect 469222 254218 504986 254454
rect 505222 254218 540986 254454
rect 541222 254218 576986 254454
rect 577222 254218 585502 254454
rect 585738 254218 586840 254454
rect -2916 254134 586840 254218
rect -2916 253898 -1814 254134
rect -1578 253898 986 254134
rect 1222 253898 36986 254134
rect 37222 253898 72986 254134
rect 73222 253898 108986 254134
rect 109222 253898 144986 254134
rect 145222 253898 180986 254134
rect 181222 253898 216986 254134
rect 217222 253898 252986 254134
rect 253222 253898 288986 254134
rect 289222 253898 324986 254134
rect 325222 253898 360986 254134
rect 361222 253898 396986 254134
rect 397222 253898 432986 254134
rect 433222 253898 468986 254134
rect 469222 253898 504986 254134
rect 505222 253898 540986 254134
rect 541222 253898 576986 254134
rect 577222 253898 585502 254134
rect 585738 253898 586840 254134
rect -2916 253876 586840 253898
rect -1996 253874 -1396 253876
rect 804 253874 1404 253876
rect 36804 253874 37404 253876
rect 72804 253874 73404 253876
rect 108804 253874 109404 253876
rect 144804 253874 145404 253876
rect 180804 253874 181404 253876
rect 216804 253874 217404 253876
rect 252804 253874 253404 253876
rect 288804 253874 289404 253876
rect 324804 253874 325404 253876
rect 360804 253874 361404 253876
rect 396804 253874 397404 253876
rect 432804 253874 433404 253876
rect 468804 253874 469404 253876
rect 504804 253874 505404 253876
rect 540804 253874 541404 253876
rect 576804 253874 577404 253876
rect 585320 253874 585920 253876
rect -8436 247276 -7836 247278
rect 29604 247276 30204 247278
rect 65604 247276 66204 247278
rect 101604 247276 102204 247278
rect 137604 247276 138204 247278
rect 173604 247276 174204 247278
rect 209604 247276 210204 247278
rect 245604 247276 246204 247278
rect 281604 247276 282204 247278
rect 317604 247276 318204 247278
rect 353604 247276 354204 247278
rect 389604 247276 390204 247278
rect 425604 247276 426204 247278
rect 461604 247276 462204 247278
rect 497604 247276 498204 247278
rect 533604 247276 534204 247278
rect 569604 247276 570204 247278
rect 591760 247276 592360 247278
rect -8436 247254 592360 247276
rect -8436 247018 -8254 247254
rect -8018 247018 29786 247254
rect 30022 247018 65786 247254
rect 66022 247018 101786 247254
rect 102022 247018 137786 247254
rect 138022 247018 173786 247254
rect 174022 247018 209786 247254
rect 210022 247018 245786 247254
rect 246022 247018 281786 247254
rect 282022 247018 317786 247254
rect 318022 247018 353786 247254
rect 354022 247018 389786 247254
rect 390022 247018 425786 247254
rect 426022 247018 461786 247254
rect 462022 247018 497786 247254
rect 498022 247018 533786 247254
rect 534022 247018 569786 247254
rect 570022 247018 591942 247254
rect 592178 247018 592360 247254
rect -8436 246934 592360 247018
rect -8436 246698 -8254 246934
rect -8018 246698 29786 246934
rect 30022 246698 65786 246934
rect 66022 246698 101786 246934
rect 102022 246698 137786 246934
rect 138022 246698 173786 246934
rect 174022 246698 209786 246934
rect 210022 246698 245786 246934
rect 246022 246698 281786 246934
rect 282022 246698 317786 246934
rect 318022 246698 353786 246934
rect 354022 246698 389786 246934
rect 390022 246698 425786 246934
rect 426022 246698 461786 246934
rect 462022 246698 497786 246934
rect 498022 246698 533786 246934
rect 534022 246698 569786 246934
rect 570022 246698 591942 246934
rect 592178 246698 592360 246934
rect -8436 246676 592360 246698
rect -8436 246674 -7836 246676
rect 29604 246674 30204 246676
rect 65604 246674 66204 246676
rect 101604 246674 102204 246676
rect 137604 246674 138204 246676
rect 173604 246674 174204 246676
rect 209604 246674 210204 246676
rect 245604 246674 246204 246676
rect 281604 246674 282204 246676
rect 317604 246674 318204 246676
rect 353604 246674 354204 246676
rect 389604 246674 390204 246676
rect 425604 246674 426204 246676
rect 461604 246674 462204 246676
rect 497604 246674 498204 246676
rect 533604 246674 534204 246676
rect 569604 246674 570204 246676
rect 591760 246674 592360 246676
rect -6596 243676 -5996 243678
rect 26004 243676 26604 243678
rect 62004 243676 62604 243678
rect 98004 243676 98604 243678
rect 134004 243676 134604 243678
rect 170004 243676 170604 243678
rect 206004 243676 206604 243678
rect 242004 243676 242604 243678
rect 278004 243676 278604 243678
rect 314004 243676 314604 243678
rect 350004 243676 350604 243678
rect 386004 243676 386604 243678
rect 422004 243676 422604 243678
rect 458004 243676 458604 243678
rect 494004 243676 494604 243678
rect 530004 243676 530604 243678
rect 566004 243676 566604 243678
rect 589920 243676 590520 243678
rect -6596 243654 590520 243676
rect -6596 243418 -6414 243654
rect -6178 243418 26186 243654
rect 26422 243418 62186 243654
rect 62422 243418 98186 243654
rect 98422 243418 134186 243654
rect 134422 243418 170186 243654
rect 170422 243418 206186 243654
rect 206422 243418 242186 243654
rect 242422 243418 278186 243654
rect 278422 243418 314186 243654
rect 314422 243418 350186 243654
rect 350422 243418 386186 243654
rect 386422 243418 422186 243654
rect 422422 243418 458186 243654
rect 458422 243418 494186 243654
rect 494422 243418 530186 243654
rect 530422 243418 566186 243654
rect 566422 243418 590102 243654
rect 590338 243418 590520 243654
rect -6596 243334 590520 243418
rect -6596 243098 -6414 243334
rect -6178 243098 26186 243334
rect 26422 243098 62186 243334
rect 62422 243098 98186 243334
rect 98422 243098 134186 243334
rect 134422 243098 170186 243334
rect 170422 243098 206186 243334
rect 206422 243098 242186 243334
rect 242422 243098 278186 243334
rect 278422 243098 314186 243334
rect 314422 243098 350186 243334
rect 350422 243098 386186 243334
rect 386422 243098 422186 243334
rect 422422 243098 458186 243334
rect 458422 243098 494186 243334
rect 494422 243098 530186 243334
rect 530422 243098 566186 243334
rect 566422 243098 590102 243334
rect 590338 243098 590520 243334
rect -6596 243076 590520 243098
rect -6596 243074 -5996 243076
rect 26004 243074 26604 243076
rect 62004 243074 62604 243076
rect 98004 243074 98604 243076
rect 134004 243074 134604 243076
rect 170004 243074 170604 243076
rect 206004 243074 206604 243076
rect 242004 243074 242604 243076
rect 278004 243074 278604 243076
rect 314004 243074 314604 243076
rect 350004 243074 350604 243076
rect 386004 243074 386604 243076
rect 422004 243074 422604 243076
rect 458004 243074 458604 243076
rect 494004 243074 494604 243076
rect 530004 243074 530604 243076
rect 566004 243074 566604 243076
rect 589920 243074 590520 243076
rect -4756 240076 -4156 240078
rect 22404 240076 23004 240078
rect 58404 240076 59004 240078
rect 94404 240076 95004 240078
rect 130404 240076 131004 240078
rect 166404 240076 167004 240078
rect 202404 240076 203004 240078
rect 238404 240076 239004 240078
rect 274404 240076 275004 240078
rect 310404 240076 311004 240078
rect 346404 240076 347004 240078
rect 382404 240076 383004 240078
rect 418404 240076 419004 240078
rect 454404 240076 455004 240078
rect 490404 240076 491004 240078
rect 526404 240076 527004 240078
rect 562404 240076 563004 240078
rect 588080 240076 588680 240078
rect -4756 240054 588680 240076
rect -4756 239818 -4574 240054
rect -4338 239818 22586 240054
rect 22822 239818 58586 240054
rect 58822 239818 94586 240054
rect 94822 239818 130586 240054
rect 130822 239818 166586 240054
rect 166822 239818 202586 240054
rect 202822 239818 238586 240054
rect 238822 239818 274586 240054
rect 274822 239818 310586 240054
rect 310822 239818 346586 240054
rect 346822 239818 382586 240054
rect 382822 239818 418586 240054
rect 418822 239818 454586 240054
rect 454822 239818 490586 240054
rect 490822 239818 526586 240054
rect 526822 239818 562586 240054
rect 562822 239818 588262 240054
rect 588498 239818 588680 240054
rect -4756 239734 588680 239818
rect -4756 239498 -4574 239734
rect -4338 239498 22586 239734
rect 22822 239498 58586 239734
rect 58822 239498 94586 239734
rect 94822 239498 130586 239734
rect 130822 239498 166586 239734
rect 166822 239498 202586 239734
rect 202822 239498 238586 239734
rect 238822 239498 274586 239734
rect 274822 239498 310586 239734
rect 310822 239498 346586 239734
rect 346822 239498 382586 239734
rect 382822 239498 418586 239734
rect 418822 239498 454586 239734
rect 454822 239498 490586 239734
rect 490822 239498 526586 239734
rect 526822 239498 562586 239734
rect 562822 239498 588262 239734
rect 588498 239498 588680 239734
rect -4756 239476 588680 239498
rect -4756 239474 -4156 239476
rect 22404 239474 23004 239476
rect 58404 239474 59004 239476
rect 94404 239474 95004 239476
rect 130404 239474 131004 239476
rect 166404 239474 167004 239476
rect 202404 239474 203004 239476
rect 238404 239474 239004 239476
rect 274404 239474 275004 239476
rect 310404 239474 311004 239476
rect 346404 239474 347004 239476
rect 382404 239474 383004 239476
rect 418404 239474 419004 239476
rect 454404 239474 455004 239476
rect 490404 239474 491004 239476
rect 526404 239474 527004 239476
rect 562404 239474 563004 239476
rect 588080 239474 588680 239476
rect -2916 236476 -2316 236478
rect 18804 236476 19404 236478
rect 54804 236476 55404 236478
rect 90804 236476 91404 236478
rect 126804 236476 127404 236478
rect 162804 236476 163404 236478
rect 198804 236476 199404 236478
rect 234804 236476 235404 236478
rect 270804 236476 271404 236478
rect 306804 236476 307404 236478
rect 342804 236476 343404 236478
rect 378804 236476 379404 236478
rect 414804 236476 415404 236478
rect 450804 236476 451404 236478
rect 486804 236476 487404 236478
rect 522804 236476 523404 236478
rect 558804 236476 559404 236478
rect 586240 236476 586840 236478
rect -2916 236454 586840 236476
rect -2916 236218 -2734 236454
rect -2498 236218 18986 236454
rect 19222 236218 54986 236454
rect 55222 236218 90986 236454
rect 91222 236218 126986 236454
rect 127222 236218 162986 236454
rect 163222 236218 198986 236454
rect 199222 236218 234986 236454
rect 235222 236218 270986 236454
rect 271222 236218 306986 236454
rect 307222 236218 342986 236454
rect 343222 236218 378986 236454
rect 379222 236218 414986 236454
rect 415222 236218 450986 236454
rect 451222 236218 486986 236454
rect 487222 236218 522986 236454
rect 523222 236218 558986 236454
rect 559222 236218 586422 236454
rect 586658 236218 586840 236454
rect -2916 236134 586840 236218
rect -2916 235898 -2734 236134
rect -2498 235898 18986 236134
rect 19222 235898 54986 236134
rect 55222 235898 90986 236134
rect 91222 235898 126986 236134
rect 127222 235898 162986 236134
rect 163222 235898 198986 236134
rect 199222 235898 234986 236134
rect 235222 235898 270986 236134
rect 271222 235898 306986 236134
rect 307222 235898 342986 236134
rect 343222 235898 378986 236134
rect 379222 235898 414986 236134
rect 415222 235898 450986 236134
rect 451222 235898 486986 236134
rect 487222 235898 522986 236134
rect 523222 235898 558986 236134
rect 559222 235898 586422 236134
rect 586658 235898 586840 236134
rect -2916 235876 586840 235898
rect -2916 235874 -2316 235876
rect 18804 235874 19404 235876
rect 54804 235874 55404 235876
rect 90804 235874 91404 235876
rect 126804 235874 127404 235876
rect 162804 235874 163404 235876
rect 198804 235874 199404 235876
rect 234804 235874 235404 235876
rect 270804 235874 271404 235876
rect 306804 235874 307404 235876
rect 342804 235874 343404 235876
rect 378804 235874 379404 235876
rect 414804 235874 415404 235876
rect 450804 235874 451404 235876
rect 486804 235874 487404 235876
rect 522804 235874 523404 235876
rect 558804 235874 559404 235876
rect 586240 235874 586840 235876
rect -7516 229276 -6916 229278
rect 11604 229276 12204 229278
rect 47604 229276 48204 229278
rect 83604 229276 84204 229278
rect 119604 229276 120204 229278
rect 155604 229276 156204 229278
rect 191604 229276 192204 229278
rect 227604 229276 228204 229278
rect 263604 229276 264204 229278
rect 299604 229276 300204 229278
rect 335604 229276 336204 229278
rect 371604 229276 372204 229278
rect 407604 229276 408204 229278
rect 443604 229276 444204 229278
rect 479604 229276 480204 229278
rect 515604 229276 516204 229278
rect 551604 229276 552204 229278
rect 590840 229276 591440 229278
rect -8436 229254 592360 229276
rect -8436 229018 -7334 229254
rect -7098 229018 11786 229254
rect 12022 229018 47786 229254
rect 48022 229018 83786 229254
rect 84022 229018 119786 229254
rect 120022 229018 155786 229254
rect 156022 229018 191786 229254
rect 192022 229018 227786 229254
rect 228022 229018 263786 229254
rect 264022 229018 299786 229254
rect 300022 229018 335786 229254
rect 336022 229018 371786 229254
rect 372022 229018 407786 229254
rect 408022 229018 443786 229254
rect 444022 229018 479786 229254
rect 480022 229018 515786 229254
rect 516022 229018 551786 229254
rect 552022 229018 591022 229254
rect 591258 229018 592360 229254
rect -8436 228934 592360 229018
rect -8436 228698 -7334 228934
rect -7098 228698 11786 228934
rect 12022 228698 47786 228934
rect 48022 228698 83786 228934
rect 84022 228698 119786 228934
rect 120022 228698 155786 228934
rect 156022 228698 191786 228934
rect 192022 228698 227786 228934
rect 228022 228698 263786 228934
rect 264022 228698 299786 228934
rect 300022 228698 335786 228934
rect 336022 228698 371786 228934
rect 372022 228698 407786 228934
rect 408022 228698 443786 228934
rect 444022 228698 479786 228934
rect 480022 228698 515786 228934
rect 516022 228698 551786 228934
rect 552022 228698 591022 228934
rect 591258 228698 592360 228934
rect -8436 228676 592360 228698
rect -7516 228674 -6916 228676
rect 11604 228674 12204 228676
rect 47604 228674 48204 228676
rect 83604 228674 84204 228676
rect 119604 228674 120204 228676
rect 155604 228674 156204 228676
rect 191604 228674 192204 228676
rect 227604 228674 228204 228676
rect 263604 228674 264204 228676
rect 299604 228674 300204 228676
rect 335604 228674 336204 228676
rect 371604 228674 372204 228676
rect 407604 228674 408204 228676
rect 443604 228674 444204 228676
rect 479604 228674 480204 228676
rect 515604 228674 516204 228676
rect 551604 228674 552204 228676
rect 590840 228674 591440 228676
rect -5676 225676 -5076 225678
rect 8004 225676 8604 225678
rect 44004 225676 44604 225678
rect 80004 225676 80604 225678
rect 116004 225676 116604 225678
rect 152004 225676 152604 225678
rect 188004 225676 188604 225678
rect 224004 225676 224604 225678
rect 260004 225676 260604 225678
rect 296004 225676 296604 225678
rect 332004 225676 332604 225678
rect 368004 225676 368604 225678
rect 404004 225676 404604 225678
rect 440004 225676 440604 225678
rect 476004 225676 476604 225678
rect 512004 225676 512604 225678
rect 548004 225676 548604 225678
rect 589000 225676 589600 225678
rect -6596 225654 590520 225676
rect -6596 225418 -5494 225654
rect -5258 225418 8186 225654
rect 8422 225418 44186 225654
rect 44422 225418 80186 225654
rect 80422 225418 116186 225654
rect 116422 225418 152186 225654
rect 152422 225418 188186 225654
rect 188422 225418 224186 225654
rect 224422 225418 260186 225654
rect 260422 225418 296186 225654
rect 296422 225418 332186 225654
rect 332422 225418 368186 225654
rect 368422 225418 404186 225654
rect 404422 225418 440186 225654
rect 440422 225418 476186 225654
rect 476422 225418 512186 225654
rect 512422 225418 548186 225654
rect 548422 225418 589182 225654
rect 589418 225418 590520 225654
rect -6596 225334 590520 225418
rect -6596 225098 -5494 225334
rect -5258 225098 8186 225334
rect 8422 225098 44186 225334
rect 44422 225098 80186 225334
rect 80422 225098 116186 225334
rect 116422 225098 152186 225334
rect 152422 225098 188186 225334
rect 188422 225098 224186 225334
rect 224422 225098 260186 225334
rect 260422 225098 296186 225334
rect 296422 225098 332186 225334
rect 332422 225098 368186 225334
rect 368422 225098 404186 225334
rect 404422 225098 440186 225334
rect 440422 225098 476186 225334
rect 476422 225098 512186 225334
rect 512422 225098 548186 225334
rect 548422 225098 589182 225334
rect 589418 225098 590520 225334
rect -6596 225076 590520 225098
rect -5676 225074 -5076 225076
rect 8004 225074 8604 225076
rect 44004 225074 44604 225076
rect 80004 225074 80604 225076
rect 116004 225074 116604 225076
rect 152004 225074 152604 225076
rect 188004 225074 188604 225076
rect 224004 225074 224604 225076
rect 260004 225074 260604 225076
rect 296004 225074 296604 225076
rect 332004 225074 332604 225076
rect 368004 225074 368604 225076
rect 404004 225074 404604 225076
rect 440004 225074 440604 225076
rect 476004 225074 476604 225076
rect 512004 225074 512604 225076
rect 548004 225074 548604 225076
rect 589000 225074 589600 225076
rect -3836 222076 -3236 222078
rect 4404 222076 5004 222078
rect 40404 222076 41004 222078
rect 76404 222076 77004 222078
rect 112404 222076 113004 222078
rect 148404 222076 149004 222078
rect 184404 222076 185004 222078
rect 220404 222076 221004 222078
rect 256404 222076 257004 222078
rect 292404 222076 293004 222078
rect 328404 222076 329004 222078
rect 364404 222076 365004 222078
rect 400404 222076 401004 222078
rect 436404 222076 437004 222078
rect 472404 222076 473004 222078
rect 508404 222076 509004 222078
rect 544404 222076 545004 222078
rect 580404 222076 581004 222078
rect 587160 222076 587760 222078
rect -4756 222054 588680 222076
rect -4756 221818 -3654 222054
rect -3418 221818 4586 222054
rect 4822 221818 40586 222054
rect 40822 221818 76586 222054
rect 76822 221818 112586 222054
rect 112822 221818 148586 222054
rect 148822 221818 184586 222054
rect 184822 221818 220586 222054
rect 220822 221818 256586 222054
rect 256822 221818 292586 222054
rect 292822 221818 328586 222054
rect 328822 221818 364586 222054
rect 364822 221818 400586 222054
rect 400822 221818 436586 222054
rect 436822 221818 472586 222054
rect 472822 221818 508586 222054
rect 508822 221818 544586 222054
rect 544822 221818 580586 222054
rect 580822 221818 587342 222054
rect 587578 221818 588680 222054
rect -4756 221734 588680 221818
rect -4756 221498 -3654 221734
rect -3418 221498 4586 221734
rect 4822 221498 40586 221734
rect 40822 221498 76586 221734
rect 76822 221498 112586 221734
rect 112822 221498 148586 221734
rect 148822 221498 184586 221734
rect 184822 221498 220586 221734
rect 220822 221498 256586 221734
rect 256822 221498 292586 221734
rect 292822 221498 328586 221734
rect 328822 221498 364586 221734
rect 364822 221498 400586 221734
rect 400822 221498 436586 221734
rect 436822 221498 472586 221734
rect 472822 221498 508586 221734
rect 508822 221498 544586 221734
rect 544822 221498 580586 221734
rect 580822 221498 587342 221734
rect 587578 221498 588680 221734
rect -4756 221476 588680 221498
rect -3836 221474 -3236 221476
rect 4404 221474 5004 221476
rect 40404 221474 41004 221476
rect 76404 221474 77004 221476
rect 112404 221474 113004 221476
rect 148404 221474 149004 221476
rect 184404 221474 185004 221476
rect 220404 221474 221004 221476
rect 256404 221474 257004 221476
rect 292404 221474 293004 221476
rect 328404 221474 329004 221476
rect 364404 221474 365004 221476
rect 400404 221474 401004 221476
rect 436404 221474 437004 221476
rect 472404 221474 473004 221476
rect 508404 221474 509004 221476
rect 544404 221474 545004 221476
rect 580404 221474 581004 221476
rect 587160 221474 587760 221476
rect -1996 218476 -1396 218478
rect 804 218476 1404 218478
rect 36804 218476 37404 218478
rect 72804 218476 73404 218478
rect 108804 218476 109404 218478
rect 144804 218476 145404 218478
rect 180804 218476 181404 218478
rect 216804 218476 217404 218478
rect 252804 218476 253404 218478
rect 288804 218476 289404 218478
rect 324804 218476 325404 218478
rect 360804 218476 361404 218478
rect 396804 218476 397404 218478
rect 432804 218476 433404 218478
rect 468804 218476 469404 218478
rect 504804 218476 505404 218478
rect 540804 218476 541404 218478
rect 576804 218476 577404 218478
rect 585320 218476 585920 218478
rect -2916 218454 586840 218476
rect -2916 218218 -1814 218454
rect -1578 218218 986 218454
rect 1222 218218 36986 218454
rect 37222 218218 72986 218454
rect 73222 218218 108986 218454
rect 109222 218218 144986 218454
rect 145222 218218 180986 218454
rect 181222 218218 216986 218454
rect 217222 218218 252986 218454
rect 253222 218218 288986 218454
rect 289222 218218 324986 218454
rect 325222 218218 360986 218454
rect 361222 218218 396986 218454
rect 397222 218218 432986 218454
rect 433222 218218 468986 218454
rect 469222 218218 504986 218454
rect 505222 218218 540986 218454
rect 541222 218218 576986 218454
rect 577222 218218 585502 218454
rect 585738 218218 586840 218454
rect -2916 218134 586840 218218
rect -2916 217898 -1814 218134
rect -1578 217898 986 218134
rect 1222 217898 36986 218134
rect 37222 217898 72986 218134
rect 73222 217898 108986 218134
rect 109222 217898 144986 218134
rect 145222 217898 180986 218134
rect 181222 217898 216986 218134
rect 217222 217898 252986 218134
rect 253222 217898 288986 218134
rect 289222 217898 324986 218134
rect 325222 217898 360986 218134
rect 361222 217898 396986 218134
rect 397222 217898 432986 218134
rect 433222 217898 468986 218134
rect 469222 217898 504986 218134
rect 505222 217898 540986 218134
rect 541222 217898 576986 218134
rect 577222 217898 585502 218134
rect 585738 217898 586840 218134
rect -2916 217876 586840 217898
rect -1996 217874 -1396 217876
rect 804 217874 1404 217876
rect 36804 217874 37404 217876
rect 72804 217874 73404 217876
rect 108804 217874 109404 217876
rect 144804 217874 145404 217876
rect 180804 217874 181404 217876
rect 216804 217874 217404 217876
rect 252804 217874 253404 217876
rect 288804 217874 289404 217876
rect 324804 217874 325404 217876
rect 360804 217874 361404 217876
rect 396804 217874 397404 217876
rect 432804 217874 433404 217876
rect 468804 217874 469404 217876
rect 504804 217874 505404 217876
rect 540804 217874 541404 217876
rect 576804 217874 577404 217876
rect 585320 217874 585920 217876
rect -8436 211276 -7836 211278
rect 29604 211276 30204 211278
rect 65604 211276 66204 211278
rect 101604 211276 102204 211278
rect 137604 211276 138204 211278
rect 173604 211276 174204 211278
rect 209604 211276 210204 211278
rect 245604 211276 246204 211278
rect 281604 211276 282204 211278
rect 317604 211276 318204 211278
rect 353604 211276 354204 211278
rect 389604 211276 390204 211278
rect 425604 211276 426204 211278
rect 461604 211276 462204 211278
rect 497604 211276 498204 211278
rect 533604 211276 534204 211278
rect 569604 211276 570204 211278
rect 591760 211276 592360 211278
rect -8436 211254 592360 211276
rect -8436 211018 -8254 211254
rect -8018 211018 29786 211254
rect 30022 211018 65786 211254
rect 66022 211018 101786 211254
rect 102022 211018 137786 211254
rect 138022 211018 173786 211254
rect 174022 211018 209786 211254
rect 210022 211018 245786 211254
rect 246022 211018 281786 211254
rect 282022 211018 317786 211254
rect 318022 211018 353786 211254
rect 354022 211018 389786 211254
rect 390022 211018 425786 211254
rect 426022 211018 461786 211254
rect 462022 211018 497786 211254
rect 498022 211018 533786 211254
rect 534022 211018 569786 211254
rect 570022 211018 591942 211254
rect 592178 211018 592360 211254
rect -8436 210934 592360 211018
rect -8436 210698 -8254 210934
rect -8018 210698 29786 210934
rect 30022 210698 65786 210934
rect 66022 210698 101786 210934
rect 102022 210698 137786 210934
rect 138022 210698 173786 210934
rect 174022 210698 209786 210934
rect 210022 210698 245786 210934
rect 246022 210698 281786 210934
rect 282022 210698 317786 210934
rect 318022 210698 353786 210934
rect 354022 210698 389786 210934
rect 390022 210698 425786 210934
rect 426022 210698 461786 210934
rect 462022 210698 497786 210934
rect 498022 210698 533786 210934
rect 534022 210698 569786 210934
rect 570022 210698 591942 210934
rect 592178 210698 592360 210934
rect -8436 210676 592360 210698
rect -8436 210674 -7836 210676
rect 29604 210674 30204 210676
rect 65604 210674 66204 210676
rect 101604 210674 102204 210676
rect 137604 210674 138204 210676
rect 173604 210674 174204 210676
rect 209604 210674 210204 210676
rect 245604 210674 246204 210676
rect 281604 210674 282204 210676
rect 317604 210674 318204 210676
rect 353604 210674 354204 210676
rect 389604 210674 390204 210676
rect 425604 210674 426204 210676
rect 461604 210674 462204 210676
rect 497604 210674 498204 210676
rect 533604 210674 534204 210676
rect 569604 210674 570204 210676
rect 591760 210674 592360 210676
rect -6596 207676 -5996 207678
rect 26004 207676 26604 207678
rect 62004 207676 62604 207678
rect 98004 207676 98604 207678
rect 134004 207676 134604 207678
rect 170004 207676 170604 207678
rect 206004 207676 206604 207678
rect 242004 207676 242604 207678
rect 278004 207676 278604 207678
rect 314004 207676 314604 207678
rect 350004 207676 350604 207678
rect 386004 207676 386604 207678
rect 422004 207676 422604 207678
rect 458004 207676 458604 207678
rect 494004 207676 494604 207678
rect 530004 207676 530604 207678
rect 566004 207676 566604 207678
rect 589920 207676 590520 207678
rect -6596 207654 590520 207676
rect -6596 207418 -6414 207654
rect -6178 207418 26186 207654
rect 26422 207418 62186 207654
rect 62422 207418 98186 207654
rect 98422 207418 134186 207654
rect 134422 207418 170186 207654
rect 170422 207418 206186 207654
rect 206422 207418 242186 207654
rect 242422 207418 278186 207654
rect 278422 207418 314186 207654
rect 314422 207418 350186 207654
rect 350422 207418 386186 207654
rect 386422 207418 422186 207654
rect 422422 207418 458186 207654
rect 458422 207418 494186 207654
rect 494422 207418 530186 207654
rect 530422 207418 566186 207654
rect 566422 207418 590102 207654
rect 590338 207418 590520 207654
rect -6596 207334 590520 207418
rect -6596 207098 -6414 207334
rect -6178 207098 26186 207334
rect 26422 207098 62186 207334
rect 62422 207098 98186 207334
rect 98422 207098 134186 207334
rect 134422 207098 170186 207334
rect 170422 207098 206186 207334
rect 206422 207098 242186 207334
rect 242422 207098 278186 207334
rect 278422 207098 314186 207334
rect 314422 207098 350186 207334
rect 350422 207098 386186 207334
rect 386422 207098 422186 207334
rect 422422 207098 458186 207334
rect 458422 207098 494186 207334
rect 494422 207098 530186 207334
rect 530422 207098 566186 207334
rect 566422 207098 590102 207334
rect 590338 207098 590520 207334
rect -6596 207076 590520 207098
rect -6596 207074 -5996 207076
rect 26004 207074 26604 207076
rect 62004 207074 62604 207076
rect 98004 207074 98604 207076
rect 134004 207074 134604 207076
rect 170004 207074 170604 207076
rect 206004 207074 206604 207076
rect 242004 207074 242604 207076
rect 278004 207074 278604 207076
rect 314004 207074 314604 207076
rect 350004 207074 350604 207076
rect 386004 207074 386604 207076
rect 422004 207074 422604 207076
rect 458004 207074 458604 207076
rect 494004 207074 494604 207076
rect 530004 207074 530604 207076
rect 566004 207074 566604 207076
rect 589920 207074 590520 207076
rect -4756 204076 -4156 204078
rect 22404 204076 23004 204078
rect 58404 204076 59004 204078
rect 94404 204076 95004 204078
rect 130404 204076 131004 204078
rect 166404 204076 167004 204078
rect 202404 204076 203004 204078
rect 238404 204076 239004 204078
rect 274404 204076 275004 204078
rect 310404 204076 311004 204078
rect 346404 204076 347004 204078
rect 382404 204076 383004 204078
rect 418404 204076 419004 204078
rect 454404 204076 455004 204078
rect 490404 204076 491004 204078
rect 526404 204076 527004 204078
rect 562404 204076 563004 204078
rect 588080 204076 588680 204078
rect -4756 204054 588680 204076
rect -4756 203818 -4574 204054
rect -4338 203818 22586 204054
rect 22822 203818 58586 204054
rect 58822 203818 94586 204054
rect 94822 203818 130586 204054
rect 130822 203818 166586 204054
rect 166822 203818 202586 204054
rect 202822 203818 238586 204054
rect 238822 203818 274586 204054
rect 274822 203818 310586 204054
rect 310822 203818 346586 204054
rect 346822 203818 382586 204054
rect 382822 203818 418586 204054
rect 418822 203818 454586 204054
rect 454822 203818 490586 204054
rect 490822 203818 526586 204054
rect 526822 203818 562586 204054
rect 562822 203818 588262 204054
rect 588498 203818 588680 204054
rect -4756 203734 588680 203818
rect -4756 203498 -4574 203734
rect -4338 203498 22586 203734
rect 22822 203498 58586 203734
rect 58822 203498 94586 203734
rect 94822 203498 130586 203734
rect 130822 203498 166586 203734
rect 166822 203498 202586 203734
rect 202822 203498 238586 203734
rect 238822 203498 274586 203734
rect 274822 203498 310586 203734
rect 310822 203498 346586 203734
rect 346822 203498 382586 203734
rect 382822 203498 418586 203734
rect 418822 203498 454586 203734
rect 454822 203498 490586 203734
rect 490822 203498 526586 203734
rect 526822 203498 562586 203734
rect 562822 203498 588262 203734
rect 588498 203498 588680 203734
rect -4756 203476 588680 203498
rect -4756 203474 -4156 203476
rect 22404 203474 23004 203476
rect 58404 203474 59004 203476
rect 94404 203474 95004 203476
rect 130404 203474 131004 203476
rect 166404 203474 167004 203476
rect 202404 203474 203004 203476
rect 238404 203474 239004 203476
rect 274404 203474 275004 203476
rect 310404 203474 311004 203476
rect 346404 203474 347004 203476
rect 382404 203474 383004 203476
rect 418404 203474 419004 203476
rect 454404 203474 455004 203476
rect 490404 203474 491004 203476
rect 526404 203474 527004 203476
rect 562404 203474 563004 203476
rect 588080 203474 588680 203476
rect -2916 200476 -2316 200478
rect 18804 200476 19404 200478
rect 54804 200476 55404 200478
rect 90804 200476 91404 200478
rect 126804 200476 127404 200478
rect 162804 200476 163404 200478
rect 198804 200476 199404 200478
rect 234804 200476 235404 200478
rect 270804 200476 271404 200478
rect 306804 200476 307404 200478
rect 342804 200476 343404 200478
rect 378804 200476 379404 200478
rect 414804 200476 415404 200478
rect 450804 200476 451404 200478
rect 486804 200476 487404 200478
rect 522804 200476 523404 200478
rect 558804 200476 559404 200478
rect 586240 200476 586840 200478
rect -2916 200454 586840 200476
rect -2916 200218 -2734 200454
rect -2498 200218 18986 200454
rect 19222 200218 54986 200454
rect 55222 200218 90986 200454
rect 91222 200218 126986 200454
rect 127222 200218 162986 200454
rect 163222 200218 198986 200454
rect 199222 200218 234986 200454
rect 235222 200218 270986 200454
rect 271222 200218 306986 200454
rect 307222 200218 342986 200454
rect 343222 200218 378986 200454
rect 379222 200218 414986 200454
rect 415222 200218 450986 200454
rect 451222 200218 486986 200454
rect 487222 200218 522986 200454
rect 523222 200218 558986 200454
rect 559222 200218 586422 200454
rect 586658 200218 586840 200454
rect -2916 200134 586840 200218
rect -2916 199898 -2734 200134
rect -2498 199898 18986 200134
rect 19222 199898 54986 200134
rect 55222 199898 90986 200134
rect 91222 199898 126986 200134
rect 127222 199898 162986 200134
rect 163222 199898 198986 200134
rect 199222 199898 234986 200134
rect 235222 199898 270986 200134
rect 271222 199898 306986 200134
rect 307222 199898 342986 200134
rect 343222 199898 378986 200134
rect 379222 199898 414986 200134
rect 415222 199898 450986 200134
rect 451222 199898 486986 200134
rect 487222 199898 522986 200134
rect 523222 199898 558986 200134
rect 559222 199898 586422 200134
rect 586658 199898 586840 200134
rect -2916 199876 586840 199898
rect -2916 199874 -2316 199876
rect 18804 199874 19404 199876
rect 54804 199874 55404 199876
rect 90804 199874 91404 199876
rect 126804 199874 127404 199876
rect 162804 199874 163404 199876
rect 198804 199874 199404 199876
rect 234804 199874 235404 199876
rect 270804 199874 271404 199876
rect 306804 199874 307404 199876
rect 342804 199874 343404 199876
rect 378804 199874 379404 199876
rect 414804 199874 415404 199876
rect 450804 199874 451404 199876
rect 486804 199874 487404 199876
rect 522804 199874 523404 199876
rect 558804 199874 559404 199876
rect 586240 199874 586840 199876
rect -7516 193276 -6916 193278
rect 11604 193276 12204 193278
rect 47604 193276 48204 193278
rect 83604 193276 84204 193278
rect 119604 193276 120204 193278
rect 155604 193276 156204 193278
rect 191604 193276 192204 193278
rect 227604 193276 228204 193278
rect 263604 193276 264204 193278
rect 299604 193276 300204 193278
rect 335604 193276 336204 193278
rect 371604 193276 372204 193278
rect 407604 193276 408204 193278
rect 443604 193276 444204 193278
rect 479604 193276 480204 193278
rect 515604 193276 516204 193278
rect 551604 193276 552204 193278
rect 590840 193276 591440 193278
rect -8436 193254 592360 193276
rect -8436 193018 -7334 193254
rect -7098 193018 11786 193254
rect 12022 193018 47786 193254
rect 48022 193018 83786 193254
rect 84022 193018 119786 193254
rect 120022 193018 155786 193254
rect 156022 193018 191786 193254
rect 192022 193018 227786 193254
rect 228022 193018 263786 193254
rect 264022 193018 299786 193254
rect 300022 193018 335786 193254
rect 336022 193018 371786 193254
rect 372022 193018 407786 193254
rect 408022 193018 443786 193254
rect 444022 193018 479786 193254
rect 480022 193018 515786 193254
rect 516022 193018 551786 193254
rect 552022 193018 591022 193254
rect 591258 193018 592360 193254
rect -8436 192934 592360 193018
rect -8436 192698 -7334 192934
rect -7098 192698 11786 192934
rect 12022 192698 47786 192934
rect 48022 192698 83786 192934
rect 84022 192698 119786 192934
rect 120022 192698 155786 192934
rect 156022 192698 191786 192934
rect 192022 192698 227786 192934
rect 228022 192698 263786 192934
rect 264022 192698 299786 192934
rect 300022 192698 335786 192934
rect 336022 192698 371786 192934
rect 372022 192698 407786 192934
rect 408022 192698 443786 192934
rect 444022 192698 479786 192934
rect 480022 192698 515786 192934
rect 516022 192698 551786 192934
rect 552022 192698 591022 192934
rect 591258 192698 592360 192934
rect -8436 192676 592360 192698
rect -7516 192674 -6916 192676
rect 11604 192674 12204 192676
rect 47604 192674 48204 192676
rect 83604 192674 84204 192676
rect 119604 192674 120204 192676
rect 155604 192674 156204 192676
rect 191604 192674 192204 192676
rect 227604 192674 228204 192676
rect 263604 192674 264204 192676
rect 299604 192674 300204 192676
rect 335604 192674 336204 192676
rect 371604 192674 372204 192676
rect 407604 192674 408204 192676
rect 443604 192674 444204 192676
rect 479604 192674 480204 192676
rect 515604 192674 516204 192676
rect 551604 192674 552204 192676
rect 590840 192674 591440 192676
rect -5676 189676 -5076 189678
rect 8004 189676 8604 189678
rect 44004 189676 44604 189678
rect 80004 189676 80604 189678
rect 116004 189676 116604 189678
rect 152004 189676 152604 189678
rect 188004 189676 188604 189678
rect 224004 189676 224604 189678
rect 260004 189676 260604 189678
rect 296004 189676 296604 189678
rect 332004 189676 332604 189678
rect 368004 189676 368604 189678
rect 404004 189676 404604 189678
rect 440004 189676 440604 189678
rect 476004 189676 476604 189678
rect 512004 189676 512604 189678
rect 548004 189676 548604 189678
rect 589000 189676 589600 189678
rect -6596 189654 590520 189676
rect -6596 189418 -5494 189654
rect -5258 189418 8186 189654
rect 8422 189418 44186 189654
rect 44422 189418 80186 189654
rect 80422 189418 116186 189654
rect 116422 189418 152186 189654
rect 152422 189418 188186 189654
rect 188422 189418 224186 189654
rect 224422 189418 260186 189654
rect 260422 189418 296186 189654
rect 296422 189418 332186 189654
rect 332422 189418 368186 189654
rect 368422 189418 404186 189654
rect 404422 189418 440186 189654
rect 440422 189418 476186 189654
rect 476422 189418 512186 189654
rect 512422 189418 548186 189654
rect 548422 189418 589182 189654
rect 589418 189418 590520 189654
rect -6596 189334 590520 189418
rect -6596 189098 -5494 189334
rect -5258 189098 8186 189334
rect 8422 189098 44186 189334
rect 44422 189098 80186 189334
rect 80422 189098 116186 189334
rect 116422 189098 152186 189334
rect 152422 189098 188186 189334
rect 188422 189098 224186 189334
rect 224422 189098 260186 189334
rect 260422 189098 296186 189334
rect 296422 189098 332186 189334
rect 332422 189098 368186 189334
rect 368422 189098 404186 189334
rect 404422 189098 440186 189334
rect 440422 189098 476186 189334
rect 476422 189098 512186 189334
rect 512422 189098 548186 189334
rect 548422 189098 589182 189334
rect 589418 189098 590520 189334
rect -6596 189076 590520 189098
rect -5676 189074 -5076 189076
rect 8004 189074 8604 189076
rect 44004 189074 44604 189076
rect 80004 189074 80604 189076
rect 116004 189074 116604 189076
rect 152004 189074 152604 189076
rect 188004 189074 188604 189076
rect 224004 189074 224604 189076
rect 260004 189074 260604 189076
rect 296004 189074 296604 189076
rect 332004 189074 332604 189076
rect 368004 189074 368604 189076
rect 404004 189074 404604 189076
rect 440004 189074 440604 189076
rect 476004 189074 476604 189076
rect 512004 189074 512604 189076
rect 548004 189074 548604 189076
rect 589000 189074 589600 189076
rect -3836 186076 -3236 186078
rect 4404 186076 5004 186078
rect 40404 186076 41004 186078
rect 76404 186076 77004 186078
rect 112404 186076 113004 186078
rect 148404 186076 149004 186078
rect 184404 186076 185004 186078
rect 220404 186076 221004 186078
rect 256404 186076 257004 186078
rect 292404 186076 293004 186078
rect 328404 186076 329004 186078
rect 364404 186076 365004 186078
rect 400404 186076 401004 186078
rect 436404 186076 437004 186078
rect 472404 186076 473004 186078
rect 508404 186076 509004 186078
rect 544404 186076 545004 186078
rect 580404 186076 581004 186078
rect 587160 186076 587760 186078
rect -4756 186054 588680 186076
rect -4756 185818 -3654 186054
rect -3418 185818 4586 186054
rect 4822 185818 40586 186054
rect 40822 185818 76586 186054
rect 76822 185818 112586 186054
rect 112822 185818 148586 186054
rect 148822 185818 184586 186054
rect 184822 185818 220586 186054
rect 220822 185818 256586 186054
rect 256822 185818 292586 186054
rect 292822 185818 328586 186054
rect 328822 185818 364586 186054
rect 364822 185818 400586 186054
rect 400822 185818 436586 186054
rect 436822 185818 472586 186054
rect 472822 185818 508586 186054
rect 508822 185818 544586 186054
rect 544822 185818 580586 186054
rect 580822 185818 587342 186054
rect 587578 185818 588680 186054
rect -4756 185734 588680 185818
rect -4756 185498 -3654 185734
rect -3418 185498 4586 185734
rect 4822 185498 40586 185734
rect 40822 185498 76586 185734
rect 76822 185498 112586 185734
rect 112822 185498 148586 185734
rect 148822 185498 184586 185734
rect 184822 185498 220586 185734
rect 220822 185498 256586 185734
rect 256822 185498 292586 185734
rect 292822 185498 328586 185734
rect 328822 185498 364586 185734
rect 364822 185498 400586 185734
rect 400822 185498 436586 185734
rect 436822 185498 472586 185734
rect 472822 185498 508586 185734
rect 508822 185498 544586 185734
rect 544822 185498 580586 185734
rect 580822 185498 587342 185734
rect 587578 185498 588680 185734
rect -4756 185476 588680 185498
rect -3836 185474 -3236 185476
rect 4404 185474 5004 185476
rect 40404 185474 41004 185476
rect 76404 185474 77004 185476
rect 112404 185474 113004 185476
rect 148404 185474 149004 185476
rect 184404 185474 185004 185476
rect 220404 185474 221004 185476
rect 256404 185474 257004 185476
rect 292404 185474 293004 185476
rect 328404 185474 329004 185476
rect 364404 185474 365004 185476
rect 400404 185474 401004 185476
rect 436404 185474 437004 185476
rect 472404 185474 473004 185476
rect 508404 185474 509004 185476
rect 544404 185474 545004 185476
rect 580404 185474 581004 185476
rect 587160 185474 587760 185476
rect -1996 182476 -1396 182478
rect 804 182476 1404 182478
rect 36804 182476 37404 182478
rect 72804 182476 73404 182478
rect 108804 182476 109404 182478
rect 144804 182476 145404 182478
rect 180804 182476 181404 182478
rect 216804 182476 217404 182478
rect 252804 182476 253404 182478
rect 288804 182476 289404 182478
rect 324804 182476 325404 182478
rect 360804 182476 361404 182478
rect 396804 182476 397404 182478
rect 432804 182476 433404 182478
rect 468804 182476 469404 182478
rect 504804 182476 505404 182478
rect 540804 182476 541404 182478
rect 576804 182476 577404 182478
rect 585320 182476 585920 182478
rect -2916 182454 586840 182476
rect -2916 182218 -1814 182454
rect -1578 182218 986 182454
rect 1222 182218 36986 182454
rect 37222 182218 72986 182454
rect 73222 182218 108986 182454
rect 109222 182218 144986 182454
rect 145222 182218 180986 182454
rect 181222 182218 216986 182454
rect 217222 182218 252986 182454
rect 253222 182218 288986 182454
rect 289222 182218 324986 182454
rect 325222 182218 360986 182454
rect 361222 182218 396986 182454
rect 397222 182218 432986 182454
rect 433222 182218 468986 182454
rect 469222 182218 504986 182454
rect 505222 182218 540986 182454
rect 541222 182218 576986 182454
rect 577222 182218 585502 182454
rect 585738 182218 586840 182454
rect -2916 182134 586840 182218
rect -2916 181898 -1814 182134
rect -1578 181898 986 182134
rect 1222 181898 36986 182134
rect 37222 181898 72986 182134
rect 73222 181898 108986 182134
rect 109222 181898 144986 182134
rect 145222 181898 180986 182134
rect 181222 181898 216986 182134
rect 217222 181898 252986 182134
rect 253222 181898 288986 182134
rect 289222 181898 324986 182134
rect 325222 181898 360986 182134
rect 361222 181898 396986 182134
rect 397222 181898 432986 182134
rect 433222 181898 468986 182134
rect 469222 181898 504986 182134
rect 505222 181898 540986 182134
rect 541222 181898 576986 182134
rect 577222 181898 585502 182134
rect 585738 181898 586840 182134
rect -2916 181876 586840 181898
rect -1996 181874 -1396 181876
rect 804 181874 1404 181876
rect 36804 181874 37404 181876
rect 72804 181874 73404 181876
rect 108804 181874 109404 181876
rect 144804 181874 145404 181876
rect 180804 181874 181404 181876
rect 216804 181874 217404 181876
rect 252804 181874 253404 181876
rect 288804 181874 289404 181876
rect 324804 181874 325404 181876
rect 360804 181874 361404 181876
rect 396804 181874 397404 181876
rect 432804 181874 433404 181876
rect 468804 181874 469404 181876
rect 504804 181874 505404 181876
rect 540804 181874 541404 181876
rect 576804 181874 577404 181876
rect 585320 181874 585920 181876
rect -8436 175276 -7836 175278
rect 29604 175276 30204 175278
rect 65604 175276 66204 175278
rect 101604 175276 102204 175278
rect 137604 175276 138204 175278
rect 173604 175276 174204 175278
rect 209604 175276 210204 175278
rect 245604 175276 246204 175278
rect 281604 175276 282204 175278
rect 317604 175276 318204 175278
rect 353604 175276 354204 175278
rect 389604 175276 390204 175278
rect 425604 175276 426204 175278
rect 461604 175276 462204 175278
rect 497604 175276 498204 175278
rect 533604 175276 534204 175278
rect 569604 175276 570204 175278
rect 591760 175276 592360 175278
rect -8436 175254 592360 175276
rect -8436 175018 -8254 175254
rect -8018 175018 29786 175254
rect 30022 175018 65786 175254
rect 66022 175018 101786 175254
rect 102022 175018 137786 175254
rect 138022 175018 173786 175254
rect 174022 175018 209786 175254
rect 210022 175018 245786 175254
rect 246022 175018 281786 175254
rect 282022 175018 317786 175254
rect 318022 175018 353786 175254
rect 354022 175018 389786 175254
rect 390022 175018 425786 175254
rect 426022 175018 461786 175254
rect 462022 175018 497786 175254
rect 498022 175018 533786 175254
rect 534022 175018 569786 175254
rect 570022 175018 591942 175254
rect 592178 175018 592360 175254
rect -8436 174934 592360 175018
rect -8436 174698 -8254 174934
rect -8018 174698 29786 174934
rect 30022 174698 65786 174934
rect 66022 174698 101786 174934
rect 102022 174698 137786 174934
rect 138022 174698 173786 174934
rect 174022 174698 209786 174934
rect 210022 174698 245786 174934
rect 246022 174698 281786 174934
rect 282022 174698 317786 174934
rect 318022 174698 353786 174934
rect 354022 174698 389786 174934
rect 390022 174698 425786 174934
rect 426022 174698 461786 174934
rect 462022 174698 497786 174934
rect 498022 174698 533786 174934
rect 534022 174698 569786 174934
rect 570022 174698 591942 174934
rect 592178 174698 592360 174934
rect -8436 174676 592360 174698
rect -8436 174674 -7836 174676
rect 29604 174674 30204 174676
rect 65604 174674 66204 174676
rect 101604 174674 102204 174676
rect 137604 174674 138204 174676
rect 173604 174674 174204 174676
rect 209604 174674 210204 174676
rect 245604 174674 246204 174676
rect 281604 174674 282204 174676
rect 317604 174674 318204 174676
rect 353604 174674 354204 174676
rect 389604 174674 390204 174676
rect 425604 174674 426204 174676
rect 461604 174674 462204 174676
rect 497604 174674 498204 174676
rect 533604 174674 534204 174676
rect 569604 174674 570204 174676
rect 591760 174674 592360 174676
rect -6596 171676 -5996 171678
rect 26004 171676 26604 171678
rect 62004 171676 62604 171678
rect 98004 171676 98604 171678
rect 134004 171676 134604 171678
rect 170004 171676 170604 171678
rect 206004 171676 206604 171678
rect 242004 171676 242604 171678
rect 278004 171676 278604 171678
rect 314004 171676 314604 171678
rect 350004 171676 350604 171678
rect 386004 171676 386604 171678
rect 422004 171676 422604 171678
rect 458004 171676 458604 171678
rect 494004 171676 494604 171678
rect 530004 171676 530604 171678
rect 566004 171676 566604 171678
rect 589920 171676 590520 171678
rect -6596 171654 590520 171676
rect -6596 171418 -6414 171654
rect -6178 171418 26186 171654
rect 26422 171418 62186 171654
rect 62422 171418 98186 171654
rect 98422 171418 134186 171654
rect 134422 171418 170186 171654
rect 170422 171418 206186 171654
rect 206422 171418 242186 171654
rect 242422 171418 278186 171654
rect 278422 171418 314186 171654
rect 314422 171418 350186 171654
rect 350422 171418 386186 171654
rect 386422 171418 422186 171654
rect 422422 171418 458186 171654
rect 458422 171418 494186 171654
rect 494422 171418 530186 171654
rect 530422 171418 566186 171654
rect 566422 171418 590102 171654
rect 590338 171418 590520 171654
rect -6596 171334 590520 171418
rect -6596 171098 -6414 171334
rect -6178 171098 26186 171334
rect 26422 171098 62186 171334
rect 62422 171098 98186 171334
rect 98422 171098 134186 171334
rect 134422 171098 170186 171334
rect 170422 171098 206186 171334
rect 206422 171098 242186 171334
rect 242422 171098 278186 171334
rect 278422 171098 314186 171334
rect 314422 171098 350186 171334
rect 350422 171098 386186 171334
rect 386422 171098 422186 171334
rect 422422 171098 458186 171334
rect 458422 171098 494186 171334
rect 494422 171098 530186 171334
rect 530422 171098 566186 171334
rect 566422 171098 590102 171334
rect 590338 171098 590520 171334
rect -6596 171076 590520 171098
rect -6596 171074 -5996 171076
rect 26004 171074 26604 171076
rect 62004 171074 62604 171076
rect 98004 171074 98604 171076
rect 134004 171074 134604 171076
rect 170004 171074 170604 171076
rect 206004 171074 206604 171076
rect 242004 171074 242604 171076
rect 278004 171074 278604 171076
rect 314004 171074 314604 171076
rect 350004 171074 350604 171076
rect 386004 171074 386604 171076
rect 422004 171074 422604 171076
rect 458004 171074 458604 171076
rect 494004 171074 494604 171076
rect 530004 171074 530604 171076
rect 566004 171074 566604 171076
rect 589920 171074 590520 171076
rect -4756 168076 -4156 168078
rect 22404 168076 23004 168078
rect 58404 168076 59004 168078
rect 94404 168076 95004 168078
rect 130404 168076 131004 168078
rect 166404 168076 167004 168078
rect 202404 168076 203004 168078
rect 238404 168076 239004 168078
rect 274404 168076 275004 168078
rect 310404 168076 311004 168078
rect 346404 168076 347004 168078
rect 382404 168076 383004 168078
rect 418404 168076 419004 168078
rect 454404 168076 455004 168078
rect 490404 168076 491004 168078
rect 526404 168076 527004 168078
rect 562404 168076 563004 168078
rect 588080 168076 588680 168078
rect -4756 168054 588680 168076
rect -4756 167818 -4574 168054
rect -4338 167818 22586 168054
rect 22822 167818 58586 168054
rect 58822 167818 94586 168054
rect 94822 167818 130586 168054
rect 130822 167818 166586 168054
rect 166822 167818 202586 168054
rect 202822 167818 238586 168054
rect 238822 167818 274586 168054
rect 274822 167818 310586 168054
rect 310822 167818 346586 168054
rect 346822 167818 382586 168054
rect 382822 167818 418586 168054
rect 418822 167818 454586 168054
rect 454822 167818 490586 168054
rect 490822 167818 526586 168054
rect 526822 167818 562586 168054
rect 562822 167818 588262 168054
rect 588498 167818 588680 168054
rect -4756 167734 588680 167818
rect -4756 167498 -4574 167734
rect -4338 167498 22586 167734
rect 22822 167498 58586 167734
rect 58822 167498 94586 167734
rect 94822 167498 130586 167734
rect 130822 167498 166586 167734
rect 166822 167498 202586 167734
rect 202822 167498 238586 167734
rect 238822 167498 274586 167734
rect 274822 167498 310586 167734
rect 310822 167498 346586 167734
rect 346822 167498 382586 167734
rect 382822 167498 418586 167734
rect 418822 167498 454586 167734
rect 454822 167498 490586 167734
rect 490822 167498 526586 167734
rect 526822 167498 562586 167734
rect 562822 167498 588262 167734
rect 588498 167498 588680 167734
rect -4756 167476 588680 167498
rect -4756 167474 -4156 167476
rect 22404 167474 23004 167476
rect 58404 167474 59004 167476
rect 94404 167474 95004 167476
rect 130404 167474 131004 167476
rect 166404 167474 167004 167476
rect 202404 167474 203004 167476
rect 238404 167474 239004 167476
rect 274404 167474 275004 167476
rect 310404 167474 311004 167476
rect 346404 167474 347004 167476
rect 382404 167474 383004 167476
rect 418404 167474 419004 167476
rect 454404 167474 455004 167476
rect 490404 167474 491004 167476
rect 526404 167474 527004 167476
rect 562404 167474 563004 167476
rect 588080 167474 588680 167476
rect -2916 164476 -2316 164478
rect 18804 164476 19404 164478
rect 54804 164476 55404 164478
rect 90804 164476 91404 164478
rect 126804 164476 127404 164478
rect 162804 164476 163404 164478
rect 198804 164476 199404 164478
rect 234804 164476 235404 164478
rect 270804 164476 271404 164478
rect 306804 164476 307404 164478
rect 342804 164476 343404 164478
rect 378804 164476 379404 164478
rect 414804 164476 415404 164478
rect 450804 164476 451404 164478
rect 486804 164476 487404 164478
rect 522804 164476 523404 164478
rect 558804 164476 559404 164478
rect 586240 164476 586840 164478
rect -2916 164454 586840 164476
rect -2916 164218 -2734 164454
rect -2498 164218 18986 164454
rect 19222 164218 54986 164454
rect 55222 164218 90986 164454
rect 91222 164218 126986 164454
rect 127222 164218 162986 164454
rect 163222 164218 198986 164454
rect 199222 164218 234986 164454
rect 235222 164218 270986 164454
rect 271222 164218 306986 164454
rect 307222 164218 342986 164454
rect 343222 164218 378986 164454
rect 379222 164218 414986 164454
rect 415222 164218 450986 164454
rect 451222 164218 486986 164454
rect 487222 164218 522986 164454
rect 523222 164218 558986 164454
rect 559222 164218 586422 164454
rect 586658 164218 586840 164454
rect -2916 164134 586840 164218
rect -2916 163898 -2734 164134
rect -2498 163898 18986 164134
rect 19222 163898 54986 164134
rect 55222 163898 90986 164134
rect 91222 163898 126986 164134
rect 127222 163898 162986 164134
rect 163222 163898 198986 164134
rect 199222 163898 234986 164134
rect 235222 163898 270986 164134
rect 271222 163898 306986 164134
rect 307222 163898 342986 164134
rect 343222 163898 378986 164134
rect 379222 163898 414986 164134
rect 415222 163898 450986 164134
rect 451222 163898 486986 164134
rect 487222 163898 522986 164134
rect 523222 163898 558986 164134
rect 559222 163898 586422 164134
rect 586658 163898 586840 164134
rect -2916 163876 586840 163898
rect -2916 163874 -2316 163876
rect 18804 163874 19404 163876
rect 54804 163874 55404 163876
rect 90804 163874 91404 163876
rect 126804 163874 127404 163876
rect 162804 163874 163404 163876
rect 198804 163874 199404 163876
rect 234804 163874 235404 163876
rect 270804 163874 271404 163876
rect 306804 163874 307404 163876
rect 342804 163874 343404 163876
rect 378804 163874 379404 163876
rect 414804 163874 415404 163876
rect 450804 163874 451404 163876
rect 486804 163874 487404 163876
rect 522804 163874 523404 163876
rect 558804 163874 559404 163876
rect 586240 163874 586840 163876
rect -7516 157276 -6916 157278
rect 11604 157276 12204 157278
rect 47604 157276 48204 157278
rect 83604 157276 84204 157278
rect 119604 157276 120204 157278
rect 155604 157276 156204 157278
rect 191604 157276 192204 157278
rect 227604 157276 228204 157278
rect 263604 157276 264204 157278
rect 299604 157276 300204 157278
rect 335604 157276 336204 157278
rect 371604 157276 372204 157278
rect 407604 157276 408204 157278
rect 443604 157276 444204 157278
rect 479604 157276 480204 157278
rect 515604 157276 516204 157278
rect 551604 157276 552204 157278
rect 590840 157276 591440 157278
rect -8436 157254 592360 157276
rect -8436 157018 -7334 157254
rect -7098 157018 11786 157254
rect 12022 157018 47786 157254
rect 48022 157018 83786 157254
rect 84022 157018 119786 157254
rect 120022 157018 155786 157254
rect 156022 157018 191786 157254
rect 192022 157018 227786 157254
rect 228022 157018 263786 157254
rect 264022 157018 299786 157254
rect 300022 157018 335786 157254
rect 336022 157018 371786 157254
rect 372022 157018 407786 157254
rect 408022 157018 443786 157254
rect 444022 157018 479786 157254
rect 480022 157018 515786 157254
rect 516022 157018 551786 157254
rect 552022 157018 591022 157254
rect 591258 157018 592360 157254
rect -8436 156934 592360 157018
rect -8436 156698 -7334 156934
rect -7098 156698 11786 156934
rect 12022 156698 47786 156934
rect 48022 156698 83786 156934
rect 84022 156698 119786 156934
rect 120022 156698 155786 156934
rect 156022 156698 191786 156934
rect 192022 156698 227786 156934
rect 228022 156698 263786 156934
rect 264022 156698 299786 156934
rect 300022 156698 335786 156934
rect 336022 156698 371786 156934
rect 372022 156698 407786 156934
rect 408022 156698 443786 156934
rect 444022 156698 479786 156934
rect 480022 156698 515786 156934
rect 516022 156698 551786 156934
rect 552022 156698 591022 156934
rect 591258 156698 592360 156934
rect -8436 156676 592360 156698
rect -7516 156674 -6916 156676
rect 11604 156674 12204 156676
rect 47604 156674 48204 156676
rect 83604 156674 84204 156676
rect 119604 156674 120204 156676
rect 155604 156674 156204 156676
rect 191604 156674 192204 156676
rect 227604 156674 228204 156676
rect 263604 156674 264204 156676
rect 299604 156674 300204 156676
rect 335604 156674 336204 156676
rect 371604 156674 372204 156676
rect 407604 156674 408204 156676
rect 443604 156674 444204 156676
rect 479604 156674 480204 156676
rect 515604 156674 516204 156676
rect 551604 156674 552204 156676
rect 590840 156674 591440 156676
rect -5676 153676 -5076 153678
rect 8004 153676 8604 153678
rect 44004 153676 44604 153678
rect 80004 153676 80604 153678
rect 116004 153676 116604 153678
rect 152004 153676 152604 153678
rect 188004 153676 188604 153678
rect 224004 153676 224604 153678
rect 260004 153676 260604 153678
rect 296004 153676 296604 153678
rect 332004 153676 332604 153678
rect 368004 153676 368604 153678
rect 404004 153676 404604 153678
rect 440004 153676 440604 153678
rect 476004 153676 476604 153678
rect 512004 153676 512604 153678
rect 548004 153676 548604 153678
rect 589000 153676 589600 153678
rect -6596 153654 590520 153676
rect -6596 153418 -5494 153654
rect -5258 153418 8186 153654
rect 8422 153418 44186 153654
rect 44422 153418 80186 153654
rect 80422 153418 116186 153654
rect 116422 153418 152186 153654
rect 152422 153418 188186 153654
rect 188422 153418 224186 153654
rect 224422 153418 260186 153654
rect 260422 153418 296186 153654
rect 296422 153418 332186 153654
rect 332422 153418 368186 153654
rect 368422 153418 404186 153654
rect 404422 153418 440186 153654
rect 440422 153418 476186 153654
rect 476422 153418 512186 153654
rect 512422 153418 548186 153654
rect 548422 153418 589182 153654
rect 589418 153418 590520 153654
rect -6596 153334 590520 153418
rect -6596 153098 -5494 153334
rect -5258 153098 8186 153334
rect 8422 153098 44186 153334
rect 44422 153098 80186 153334
rect 80422 153098 116186 153334
rect 116422 153098 152186 153334
rect 152422 153098 188186 153334
rect 188422 153098 224186 153334
rect 224422 153098 260186 153334
rect 260422 153098 296186 153334
rect 296422 153098 332186 153334
rect 332422 153098 368186 153334
rect 368422 153098 404186 153334
rect 404422 153098 440186 153334
rect 440422 153098 476186 153334
rect 476422 153098 512186 153334
rect 512422 153098 548186 153334
rect 548422 153098 589182 153334
rect 589418 153098 590520 153334
rect -6596 153076 590520 153098
rect -5676 153074 -5076 153076
rect 8004 153074 8604 153076
rect 44004 153074 44604 153076
rect 80004 153074 80604 153076
rect 116004 153074 116604 153076
rect 152004 153074 152604 153076
rect 188004 153074 188604 153076
rect 224004 153074 224604 153076
rect 260004 153074 260604 153076
rect 296004 153074 296604 153076
rect 332004 153074 332604 153076
rect 368004 153074 368604 153076
rect 404004 153074 404604 153076
rect 440004 153074 440604 153076
rect 476004 153074 476604 153076
rect 512004 153074 512604 153076
rect 548004 153074 548604 153076
rect 589000 153074 589600 153076
rect -3836 150076 -3236 150078
rect 4404 150076 5004 150078
rect 40404 150076 41004 150078
rect 76404 150076 77004 150078
rect 112404 150076 113004 150078
rect 148404 150076 149004 150078
rect 184404 150076 185004 150078
rect 220404 150076 221004 150078
rect 256404 150076 257004 150078
rect 292404 150076 293004 150078
rect 328404 150076 329004 150078
rect 364404 150076 365004 150078
rect 400404 150076 401004 150078
rect 436404 150076 437004 150078
rect 472404 150076 473004 150078
rect 508404 150076 509004 150078
rect 544404 150076 545004 150078
rect 580404 150076 581004 150078
rect 587160 150076 587760 150078
rect -4756 150054 588680 150076
rect -4756 149818 -3654 150054
rect -3418 149818 4586 150054
rect 4822 149818 40586 150054
rect 40822 149818 76586 150054
rect 76822 149818 112586 150054
rect 112822 149818 148586 150054
rect 148822 149818 184586 150054
rect 184822 149818 220586 150054
rect 220822 149818 256586 150054
rect 256822 149818 292586 150054
rect 292822 149818 328586 150054
rect 328822 149818 364586 150054
rect 364822 149818 400586 150054
rect 400822 149818 436586 150054
rect 436822 149818 472586 150054
rect 472822 149818 508586 150054
rect 508822 149818 544586 150054
rect 544822 149818 580586 150054
rect 580822 149818 587342 150054
rect 587578 149818 588680 150054
rect -4756 149734 588680 149818
rect -4756 149498 -3654 149734
rect -3418 149498 4586 149734
rect 4822 149498 40586 149734
rect 40822 149498 76586 149734
rect 76822 149498 112586 149734
rect 112822 149498 148586 149734
rect 148822 149498 184586 149734
rect 184822 149498 220586 149734
rect 220822 149498 256586 149734
rect 256822 149498 292586 149734
rect 292822 149498 328586 149734
rect 328822 149498 364586 149734
rect 364822 149498 400586 149734
rect 400822 149498 436586 149734
rect 436822 149498 472586 149734
rect 472822 149498 508586 149734
rect 508822 149498 544586 149734
rect 544822 149498 580586 149734
rect 580822 149498 587342 149734
rect 587578 149498 588680 149734
rect -4756 149476 588680 149498
rect -3836 149474 -3236 149476
rect 4404 149474 5004 149476
rect 40404 149474 41004 149476
rect 76404 149474 77004 149476
rect 112404 149474 113004 149476
rect 148404 149474 149004 149476
rect 184404 149474 185004 149476
rect 220404 149474 221004 149476
rect 256404 149474 257004 149476
rect 292404 149474 293004 149476
rect 328404 149474 329004 149476
rect 364404 149474 365004 149476
rect 400404 149474 401004 149476
rect 436404 149474 437004 149476
rect 472404 149474 473004 149476
rect 508404 149474 509004 149476
rect 544404 149474 545004 149476
rect 580404 149474 581004 149476
rect 587160 149474 587760 149476
rect -1996 146476 -1396 146478
rect 804 146476 1404 146478
rect 36804 146476 37404 146478
rect 72804 146476 73404 146478
rect 108804 146476 109404 146478
rect 144804 146476 145404 146478
rect 180804 146476 181404 146478
rect 216804 146476 217404 146478
rect 252804 146476 253404 146478
rect 288804 146476 289404 146478
rect 324804 146476 325404 146478
rect 360804 146476 361404 146478
rect 396804 146476 397404 146478
rect 432804 146476 433404 146478
rect 468804 146476 469404 146478
rect 504804 146476 505404 146478
rect 540804 146476 541404 146478
rect 576804 146476 577404 146478
rect 585320 146476 585920 146478
rect -2916 146454 586840 146476
rect -2916 146218 -1814 146454
rect -1578 146218 986 146454
rect 1222 146218 36986 146454
rect 37222 146218 72986 146454
rect 73222 146218 108986 146454
rect 109222 146218 144986 146454
rect 145222 146218 180986 146454
rect 181222 146218 216986 146454
rect 217222 146218 252986 146454
rect 253222 146218 288986 146454
rect 289222 146218 324986 146454
rect 325222 146218 360986 146454
rect 361222 146218 396986 146454
rect 397222 146218 432986 146454
rect 433222 146218 468986 146454
rect 469222 146218 504986 146454
rect 505222 146218 540986 146454
rect 541222 146218 576986 146454
rect 577222 146218 585502 146454
rect 585738 146218 586840 146454
rect -2916 146134 586840 146218
rect -2916 145898 -1814 146134
rect -1578 145898 986 146134
rect 1222 145898 36986 146134
rect 37222 145898 72986 146134
rect 73222 145898 108986 146134
rect 109222 145898 144986 146134
rect 145222 145898 180986 146134
rect 181222 145898 216986 146134
rect 217222 145898 252986 146134
rect 253222 145898 288986 146134
rect 289222 145898 324986 146134
rect 325222 145898 360986 146134
rect 361222 145898 396986 146134
rect 397222 145898 432986 146134
rect 433222 145898 468986 146134
rect 469222 145898 504986 146134
rect 505222 145898 540986 146134
rect 541222 145898 576986 146134
rect 577222 145898 585502 146134
rect 585738 145898 586840 146134
rect -2916 145876 586840 145898
rect -1996 145874 -1396 145876
rect 804 145874 1404 145876
rect 36804 145874 37404 145876
rect 72804 145874 73404 145876
rect 108804 145874 109404 145876
rect 144804 145874 145404 145876
rect 180804 145874 181404 145876
rect 216804 145874 217404 145876
rect 252804 145874 253404 145876
rect 288804 145874 289404 145876
rect 324804 145874 325404 145876
rect 360804 145874 361404 145876
rect 396804 145874 397404 145876
rect 432804 145874 433404 145876
rect 468804 145874 469404 145876
rect 504804 145874 505404 145876
rect 540804 145874 541404 145876
rect 576804 145874 577404 145876
rect 585320 145874 585920 145876
rect -8436 139276 -7836 139278
rect 29604 139276 30204 139278
rect 65604 139276 66204 139278
rect 101604 139276 102204 139278
rect 137604 139276 138204 139278
rect 173604 139276 174204 139278
rect 209604 139276 210204 139278
rect 245604 139276 246204 139278
rect 281604 139276 282204 139278
rect 317604 139276 318204 139278
rect 353604 139276 354204 139278
rect 389604 139276 390204 139278
rect 425604 139276 426204 139278
rect 461604 139276 462204 139278
rect 497604 139276 498204 139278
rect 533604 139276 534204 139278
rect 569604 139276 570204 139278
rect 591760 139276 592360 139278
rect -8436 139254 592360 139276
rect -8436 139018 -8254 139254
rect -8018 139018 29786 139254
rect 30022 139018 65786 139254
rect 66022 139018 101786 139254
rect 102022 139018 137786 139254
rect 138022 139018 173786 139254
rect 174022 139018 209786 139254
rect 210022 139018 245786 139254
rect 246022 139018 281786 139254
rect 282022 139018 317786 139254
rect 318022 139018 353786 139254
rect 354022 139018 389786 139254
rect 390022 139018 425786 139254
rect 426022 139018 461786 139254
rect 462022 139018 497786 139254
rect 498022 139018 533786 139254
rect 534022 139018 569786 139254
rect 570022 139018 591942 139254
rect 592178 139018 592360 139254
rect -8436 138934 592360 139018
rect -8436 138698 -8254 138934
rect -8018 138698 29786 138934
rect 30022 138698 65786 138934
rect 66022 138698 101786 138934
rect 102022 138698 137786 138934
rect 138022 138698 173786 138934
rect 174022 138698 209786 138934
rect 210022 138698 245786 138934
rect 246022 138698 281786 138934
rect 282022 138698 317786 138934
rect 318022 138698 353786 138934
rect 354022 138698 389786 138934
rect 390022 138698 425786 138934
rect 426022 138698 461786 138934
rect 462022 138698 497786 138934
rect 498022 138698 533786 138934
rect 534022 138698 569786 138934
rect 570022 138698 591942 138934
rect 592178 138698 592360 138934
rect -8436 138676 592360 138698
rect -8436 138674 -7836 138676
rect 29604 138674 30204 138676
rect 65604 138674 66204 138676
rect 101604 138674 102204 138676
rect 137604 138674 138204 138676
rect 173604 138674 174204 138676
rect 209604 138674 210204 138676
rect 245604 138674 246204 138676
rect 281604 138674 282204 138676
rect 317604 138674 318204 138676
rect 353604 138674 354204 138676
rect 389604 138674 390204 138676
rect 425604 138674 426204 138676
rect 461604 138674 462204 138676
rect 497604 138674 498204 138676
rect 533604 138674 534204 138676
rect 569604 138674 570204 138676
rect 591760 138674 592360 138676
rect -6596 135676 -5996 135678
rect 26004 135676 26604 135678
rect 62004 135676 62604 135678
rect 98004 135676 98604 135678
rect 134004 135676 134604 135678
rect 170004 135676 170604 135678
rect 206004 135676 206604 135678
rect 242004 135676 242604 135678
rect 278004 135676 278604 135678
rect 314004 135676 314604 135678
rect 350004 135676 350604 135678
rect 386004 135676 386604 135678
rect 422004 135676 422604 135678
rect 458004 135676 458604 135678
rect 494004 135676 494604 135678
rect 530004 135676 530604 135678
rect 566004 135676 566604 135678
rect 589920 135676 590520 135678
rect -6596 135654 590520 135676
rect -6596 135418 -6414 135654
rect -6178 135418 26186 135654
rect 26422 135418 62186 135654
rect 62422 135418 98186 135654
rect 98422 135418 134186 135654
rect 134422 135418 170186 135654
rect 170422 135418 206186 135654
rect 206422 135418 242186 135654
rect 242422 135418 278186 135654
rect 278422 135418 314186 135654
rect 314422 135418 350186 135654
rect 350422 135418 386186 135654
rect 386422 135418 422186 135654
rect 422422 135418 458186 135654
rect 458422 135418 494186 135654
rect 494422 135418 530186 135654
rect 530422 135418 566186 135654
rect 566422 135418 590102 135654
rect 590338 135418 590520 135654
rect -6596 135334 590520 135418
rect -6596 135098 -6414 135334
rect -6178 135098 26186 135334
rect 26422 135098 62186 135334
rect 62422 135098 98186 135334
rect 98422 135098 134186 135334
rect 134422 135098 170186 135334
rect 170422 135098 206186 135334
rect 206422 135098 242186 135334
rect 242422 135098 278186 135334
rect 278422 135098 314186 135334
rect 314422 135098 350186 135334
rect 350422 135098 386186 135334
rect 386422 135098 422186 135334
rect 422422 135098 458186 135334
rect 458422 135098 494186 135334
rect 494422 135098 530186 135334
rect 530422 135098 566186 135334
rect 566422 135098 590102 135334
rect 590338 135098 590520 135334
rect -6596 135076 590520 135098
rect -6596 135074 -5996 135076
rect 26004 135074 26604 135076
rect 62004 135074 62604 135076
rect 98004 135074 98604 135076
rect 134004 135074 134604 135076
rect 170004 135074 170604 135076
rect 206004 135074 206604 135076
rect 242004 135074 242604 135076
rect 278004 135074 278604 135076
rect 314004 135074 314604 135076
rect 350004 135074 350604 135076
rect 386004 135074 386604 135076
rect 422004 135074 422604 135076
rect 458004 135074 458604 135076
rect 494004 135074 494604 135076
rect 530004 135074 530604 135076
rect 566004 135074 566604 135076
rect 589920 135074 590520 135076
rect -4756 132076 -4156 132078
rect 22404 132076 23004 132078
rect 58404 132076 59004 132078
rect 94404 132076 95004 132078
rect 130404 132076 131004 132078
rect 166404 132076 167004 132078
rect 202404 132076 203004 132078
rect 238404 132076 239004 132078
rect 274404 132076 275004 132078
rect 310404 132076 311004 132078
rect 346404 132076 347004 132078
rect 382404 132076 383004 132078
rect 418404 132076 419004 132078
rect 454404 132076 455004 132078
rect 490404 132076 491004 132078
rect 526404 132076 527004 132078
rect 562404 132076 563004 132078
rect 588080 132076 588680 132078
rect -4756 132054 588680 132076
rect -4756 131818 -4574 132054
rect -4338 131818 22586 132054
rect 22822 131818 58586 132054
rect 58822 131818 94586 132054
rect 94822 131818 130586 132054
rect 130822 131818 166586 132054
rect 166822 131818 202586 132054
rect 202822 131818 238586 132054
rect 238822 131818 274586 132054
rect 274822 131818 310586 132054
rect 310822 131818 346586 132054
rect 346822 131818 382586 132054
rect 382822 131818 418586 132054
rect 418822 131818 454586 132054
rect 454822 131818 490586 132054
rect 490822 131818 526586 132054
rect 526822 131818 562586 132054
rect 562822 131818 588262 132054
rect 588498 131818 588680 132054
rect -4756 131734 588680 131818
rect -4756 131498 -4574 131734
rect -4338 131498 22586 131734
rect 22822 131498 58586 131734
rect 58822 131498 94586 131734
rect 94822 131498 130586 131734
rect 130822 131498 166586 131734
rect 166822 131498 202586 131734
rect 202822 131498 238586 131734
rect 238822 131498 274586 131734
rect 274822 131498 310586 131734
rect 310822 131498 346586 131734
rect 346822 131498 382586 131734
rect 382822 131498 418586 131734
rect 418822 131498 454586 131734
rect 454822 131498 490586 131734
rect 490822 131498 526586 131734
rect 526822 131498 562586 131734
rect 562822 131498 588262 131734
rect 588498 131498 588680 131734
rect -4756 131476 588680 131498
rect -4756 131474 -4156 131476
rect 22404 131474 23004 131476
rect 58404 131474 59004 131476
rect 94404 131474 95004 131476
rect 130404 131474 131004 131476
rect 166404 131474 167004 131476
rect 202404 131474 203004 131476
rect 238404 131474 239004 131476
rect 274404 131474 275004 131476
rect 310404 131474 311004 131476
rect 346404 131474 347004 131476
rect 382404 131474 383004 131476
rect 418404 131474 419004 131476
rect 454404 131474 455004 131476
rect 490404 131474 491004 131476
rect 526404 131474 527004 131476
rect 562404 131474 563004 131476
rect 588080 131474 588680 131476
rect -2916 128476 -2316 128478
rect 18804 128476 19404 128478
rect 54804 128476 55404 128478
rect 90804 128476 91404 128478
rect 126804 128476 127404 128478
rect 162804 128476 163404 128478
rect 198804 128476 199404 128478
rect 234804 128476 235404 128478
rect 270804 128476 271404 128478
rect 306804 128476 307404 128478
rect 342804 128476 343404 128478
rect 378804 128476 379404 128478
rect 414804 128476 415404 128478
rect 450804 128476 451404 128478
rect 486804 128476 487404 128478
rect 522804 128476 523404 128478
rect 558804 128476 559404 128478
rect 586240 128476 586840 128478
rect -2916 128454 586840 128476
rect -2916 128218 -2734 128454
rect -2498 128218 18986 128454
rect 19222 128218 54986 128454
rect 55222 128218 90986 128454
rect 91222 128218 126986 128454
rect 127222 128218 162986 128454
rect 163222 128218 198986 128454
rect 199222 128218 234986 128454
rect 235222 128218 270986 128454
rect 271222 128218 306986 128454
rect 307222 128218 342986 128454
rect 343222 128218 378986 128454
rect 379222 128218 414986 128454
rect 415222 128218 450986 128454
rect 451222 128218 486986 128454
rect 487222 128218 522986 128454
rect 523222 128218 558986 128454
rect 559222 128218 586422 128454
rect 586658 128218 586840 128454
rect -2916 128134 586840 128218
rect -2916 127898 -2734 128134
rect -2498 127898 18986 128134
rect 19222 127898 54986 128134
rect 55222 127898 90986 128134
rect 91222 127898 126986 128134
rect 127222 127898 162986 128134
rect 163222 127898 198986 128134
rect 199222 127898 234986 128134
rect 235222 127898 270986 128134
rect 271222 127898 306986 128134
rect 307222 127898 342986 128134
rect 343222 127898 378986 128134
rect 379222 127898 414986 128134
rect 415222 127898 450986 128134
rect 451222 127898 486986 128134
rect 487222 127898 522986 128134
rect 523222 127898 558986 128134
rect 559222 127898 586422 128134
rect 586658 127898 586840 128134
rect -2916 127876 586840 127898
rect -2916 127874 -2316 127876
rect 18804 127874 19404 127876
rect 54804 127874 55404 127876
rect 90804 127874 91404 127876
rect 126804 127874 127404 127876
rect 162804 127874 163404 127876
rect 198804 127874 199404 127876
rect 234804 127874 235404 127876
rect 270804 127874 271404 127876
rect 306804 127874 307404 127876
rect 342804 127874 343404 127876
rect 378804 127874 379404 127876
rect 414804 127874 415404 127876
rect 450804 127874 451404 127876
rect 486804 127874 487404 127876
rect 522804 127874 523404 127876
rect 558804 127874 559404 127876
rect 586240 127874 586840 127876
rect -7516 121276 -6916 121278
rect 11604 121276 12204 121278
rect 47604 121276 48204 121278
rect 83604 121276 84204 121278
rect 119604 121276 120204 121278
rect 155604 121276 156204 121278
rect 191604 121276 192204 121278
rect 227604 121276 228204 121278
rect 263604 121276 264204 121278
rect 299604 121276 300204 121278
rect 335604 121276 336204 121278
rect 371604 121276 372204 121278
rect 407604 121276 408204 121278
rect 443604 121276 444204 121278
rect 479604 121276 480204 121278
rect 515604 121276 516204 121278
rect 551604 121276 552204 121278
rect 590840 121276 591440 121278
rect -8436 121254 592360 121276
rect -8436 121018 -7334 121254
rect -7098 121018 11786 121254
rect 12022 121018 47786 121254
rect 48022 121018 83786 121254
rect 84022 121018 119786 121254
rect 120022 121018 155786 121254
rect 156022 121018 191786 121254
rect 192022 121018 227786 121254
rect 228022 121018 263786 121254
rect 264022 121018 299786 121254
rect 300022 121018 335786 121254
rect 336022 121018 371786 121254
rect 372022 121018 407786 121254
rect 408022 121018 443786 121254
rect 444022 121018 479786 121254
rect 480022 121018 515786 121254
rect 516022 121018 551786 121254
rect 552022 121018 591022 121254
rect 591258 121018 592360 121254
rect -8436 120934 592360 121018
rect -8436 120698 -7334 120934
rect -7098 120698 11786 120934
rect 12022 120698 47786 120934
rect 48022 120698 83786 120934
rect 84022 120698 119786 120934
rect 120022 120698 155786 120934
rect 156022 120698 191786 120934
rect 192022 120698 227786 120934
rect 228022 120698 263786 120934
rect 264022 120698 299786 120934
rect 300022 120698 335786 120934
rect 336022 120698 371786 120934
rect 372022 120698 407786 120934
rect 408022 120698 443786 120934
rect 444022 120698 479786 120934
rect 480022 120698 515786 120934
rect 516022 120698 551786 120934
rect 552022 120698 591022 120934
rect 591258 120698 592360 120934
rect -8436 120676 592360 120698
rect -7516 120674 -6916 120676
rect 11604 120674 12204 120676
rect 47604 120674 48204 120676
rect 83604 120674 84204 120676
rect 119604 120674 120204 120676
rect 155604 120674 156204 120676
rect 191604 120674 192204 120676
rect 227604 120674 228204 120676
rect 263604 120674 264204 120676
rect 299604 120674 300204 120676
rect 335604 120674 336204 120676
rect 371604 120674 372204 120676
rect 407604 120674 408204 120676
rect 443604 120674 444204 120676
rect 479604 120674 480204 120676
rect 515604 120674 516204 120676
rect 551604 120674 552204 120676
rect 590840 120674 591440 120676
rect -5676 117676 -5076 117678
rect 8004 117676 8604 117678
rect 44004 117676 44604 117678
rect 80004 117676 80604 117678
rect 116004 117676 116604 117678
rect 152004 117676 152604 117678
rect 188004 117676 188604 117678
rect 224004 117676 224604 117678
rect 260004 117676 260604 117678
rect 296004 117676 296604 117678
rect 332004 117676 332604 117678
rect 368004 117676 368604 117678
rect 404004 117676 404604 117678
rect 440004 117676 440604 117678
rect 476004 117676 476604 117678
rect 512004 117676 512604 117678
rect 548004 117676 548604 117678
rect 589000 117676 589600 117678
rect -6596 117654 590520 117676
rect -6596 117418 -5494 117654
rect -5258 117418 8186 117654
rect 8422 117418 44186 117654
rect 44422 117418 80186 117654
rect 80422 117418 116186 117654
rect 116422 117418 152186 117654
rect 152422 117418 188186 117654
rect 188422 117418 224186 117654
rect 224422 117418 260186 117654
rect 260422 117418 296186 117654
rect 296422 117418 332186 117654
rect 332422 117418 368186 117654
rect 368422 117418 404186 117654
rect 404422 117418 440186 117654
rect 440422 117418 476186 117654
rect 476422 117418 512186 117654
rect 512422 117418 548186 117654
rect 548422 117418 589182 117654
rect 589418 117418 590520 117654
rect -6596 117334 590520 117418
rect -6596 117098 -5494 117334
rect -5258 117098 8186 117334
rect 8422 117098 44186 117334
rect 44422 117098 80186 117334
rect 80422 117098 116186 117334
rect 116422 117098 152186 117334
rect 152422 117098 188186 117334
rect 188422 117098 224186 117334
rect 224422 117098 260186 117334
rect 260422 117098 296186 117334
rect 296422 117098 332186 117334
rect 332422 117098 368186 117334
rect 368422 117098 404186 117334
rect 404422 117098 440186 117334
rect 440422 117098 476186 117334
rect 476422 117098 512186 117334
rect 512422 117098 548186 117334
rect 548422 117098 589182 117334
rect 589418 117098 590520 117334
rect -6596 117076 590520 117098
rect -5676 117074 -5076 117076
rect 8004 117074 8604 117076
rect 44004 117074 44604 117076
rect 80004 117074 80604 117076
rect 116004 117074 116604 117076
rect 152004 117074 152604 117076
rect 188004 117074 188604 117076
rect 224004 117074 224604 117076
rect 260004 117074 260604 117076
rect 296004 117074 296604 117076
rect 332004 117074 332604 117076
rect 368004 117074 368604 117076
rect 404004 117074 404604 117076
rect 440004 117074 440604 117076
rect 476004 117074 476604 117076
rect 512004 117074 512604 117076
rect 548004 117074 548604 117076
rect 589000 117074 589600 117076
rect -3836 114076 -3236 114078
rect 4404 114076 5004 114078
rect 40404 114076 41004 114078
rect 76404 114076 77004 114078
rect 112404 114076 113004 114078
rect 148404 114076 149004 114078
rect 184404 114076 185004 114078
rect 220404 114076 221004 114078
rect 256404 114076 257004 114078
rect 292404 114076 293004 114078
rect 328404 114076 329004 114078
rect 364404 114076 365004 114078
rect 400404 114076 401004 114078
rect 436404 114076 437004 114078
rect 472404 114076 473004 114078
rect 508404 114076 509004 114078
rect 544404 114076 545004 114078
rect 580404 114076 581004 114078
rect 587160 114076 587760 114078
rect -4756 114054 588680 114076
rect -4756 113818 -3654 114054
rect -3418 113818 4586 114054
rect 4822 113818 40586 114054
rect 40822 113818 76586 114054
rect 76822 113818 112586 114054
rect 112822 113818 148586 114054
rect 148822 113818 184586 114054
rect 184822 113818 220586 114054
rect 220822 113818 256586 114054
rect 256822 113818 292586 114054
rect 292822 113818 328586 114054
rect 328822 113818 364586 114054
rect 364822 113818 400586 114054
rect 400822 113818 436586 114054
rect 436822 113818 472586 114054
rect 472822 113818 508586 114054
rect 508822 113818 544586 114054
rect 544822 113818 580586 114054
rect 580822 113818 587342 114054
rect 587578 113818 588680 114054
rect -4756 113734 588680 113818
rect -4756 113498 -3654 113734
rect -3418 113498 4586 113734
rect 4822 113498 40586 113734
rect 40822 113498 76586 113734
rect 76822 113498 112586 113734
rect 112822 113498 148586 113734
rect 148822 113498 184586 113734
rect 184822 113498 220586 113734
rect 220822 113498 256586 113734
rect 256822 113498 292586 113734
rect 292822 113498 328586 113734
rect 328822 113498 364586 113734
rect 364822 113498 400586 113734
rect 400822 113498 436586 113734
rect 436822 113498 472586 113734
rect 472822 113498 508586 113734
rect 508822 113498 544586 113734
rect 544822 113498 580586 113734
rect 580822 113498 587342 113734
rect 587578 113498 588680 113734
rect -4756 113476 588680 113498
rect -3836 113474 -3236 113476
rect 4404 113474 5004 113476
rect 40404 113474 41004 113476
rect 76404 113474 77004 113476
rect 112404 113474 113004 113476
rect 148404 113474 149004 113476
rect 184404 113474 185004 113476
rect 220404 113474 221004 113476
rect 256404 113474 257004 113476
rect 292404 113474 293004 113476
rect 328404 113474 329004 113476
rect 364404 113474 365004 113476
rect 400404 113474 401004 113476
rect 436404 113474 437004 113476
rect 472404 113474 473004 113476
rect 508404 113474 509004 113476
rect 544404 113474 545004 113476
rect 580404 113474 581004 113476
rect 587160 113474 587760 113476
rect -1996 110476 -1396 110478
rect 804 110476 1404 110478
rect 36804 110476 37404 110478
rect 72804 110476 73404 110478
rect 108804 110476 109404 110478
rect 144804 110476 145404 110478
rect 180804 110476 181404 110478
rect 216804 110476 217404 110478
rect 252804 110476 253404 110478
rect 288804 110476 289404 110478
rect 324804 110476 325404 110478
rect 360804 110476 361404 110478
rect 396804 110476 397404 110478
rect 432804 110476 433404 110478
rect 468804 110476 469404 110478
rect 504804 110476 505404 110478
rect 540804 110476 541404 110478
rect 576804 110476 577404 110478
rect 585320 110476 585920 110478
rect -2916 110454 586840 110476
rect -2916 110218 -1814 110454
rect -1578 110218 986 110454
rect 1222 110218 36986 110454
rect 37222 110218 72986 110454
rect 73222 110218 108986 110454
rect 109222 110218 144986 110454
rect 145222 110218 180986 110454
rect 181222 110218 216986 110454
rect 217222 110218 252986 110454
rect 253222 110218 288986 110454
rect 289222 110218 324986 110454
rect 325222 110218 360986 110454
rect 361222 110218 396986 110454
rect 397222 110218 432986 110454
rect 433222 110218 468986 110454
rect 469222 110218 504986 110454
rect 505222 110218 540986 110454
rect 541222 110218 576986 110454
rect 577222 110218 585502 110454
rect 585738 110218 586840 110454
rect -2916 110134 586840 110218
rect -2916 109898 -1814 110134
rect -1578 109898 986 110134
rect 1222 109898 36986 110134
rect 37222 109898 72986 110134
rect 73222 109898 108986 110134
rect 109222 109898 144986 110134
rect 145222 109898 180986 110134
rect 181222 109898 216986 110134
rect 217222 109898 252986 110134
rect 253222 109898 288986 110134
rect 289222 109898 324986 110134
rect 325222 109898 360986 110134
rect 361222 109898 396986 110134
rect 397222 109898 432986 110134
rect 433222 109898 468986 110134
rect 469222 109898 504986 110134
rect 505222 109898 540986 110134
rect 541222 109898 576986 110134
rect 577222 109898 585502 110134
rect 585738 109898 586840 110134
rect -2916 109876 586840 109898
rect -1996 109874 -1396 109876
rect 804 109874 1404 109876
rect 36804 109874 37404 109876
rect 72804 109874 73404 109876
rect 108804 109874 109404 109876
rect 144804 109874 145404 109876
rect 180804 109874 181404 109876
rect 216804 109874 217404 109876
rect 252804 109874 253404 109876
rect 288804 109874 289404 109876
rect 324804 109874 325404 109876
rect 360804 109874 361404 109876
rect 396804 109874 397404 109876
rect 432804 109874 433404 109876
rect 468804 109874 469404 109876
rect 504804 109874 505404 109876
rect 540804 109874 541404 109876
rect 576804 109874 577404 109876
rect 585320 109874 585920 109876
rect -8436 103276 -7836 103278
rect 29604 103276 30204 103278
rect 65604 103276 66204 103278
rect 101604 103276 102204 103278
rect 137604 103276 138204 103278
rect 173604 103276 174204 103278
rect 209604 103276 210204 103278
rect 245604 103276 246204 103278
rect 281604 103276 282204 103278
rect 317604 103276 318204 103278
rect 353604 103276 354204 103278
rect 389604 103276 390204 103278
rect 425604 103276 426204 103278
rect 461604 103276 462204 103278
rect 497604 103276 498204 103278
rect 533604 103276 534204 103278
rect 569604 103276 570204 103278
rect 591760 103276 592360 103278
rect -8436 103254 592360 103276
rect -8436 103018 -8254 103254
rect -8018 103018 29786 103254
rect 30022 103018 65786 103254
rect 66022 103018 101786 103254
rect 102022 103018 137786 103254
rect 138022 103018 173786 103254
rect 174022 103018 209786 103254
rect 210022 103018 245786 103254
rect 246022 103018 281786 103254
rect 282022 103018 317786 103254
rect 318022 103018 353786 103254
rect 354022 103018 389786 103254
rect 390022 103018 425786 103254
rect 426022 103018 461786 103254
rect 462022 103018 497786 103254
rect 498022 103018 533786 103254
rect 534022 103018 569786 103254
rect 570022 103018 591942 103254
rect 592178 103018 592360 103254
rect -8436 102934 592360 103018
rect -8436 102698 -8254 102934
rect -8018 102698 29786 102934
rect 30022 102698 65786 102934
rect 66022 102698 101786 102934
rect 102022 102698 137786 102934
rect 138022 102698 173786 102934
rect 174022 102698 209786 102934
rect 210022 102698 245786 102934
rect 246022 102698 281786 102934
rect 282022 102698 317786 102934
rect 318022 102698 353786 102934
rect 354022 102698 389786 102934
rect 390022 102698 425786 102934
rect 426022 102698 461786 102934
rect 462022 102698 497786 102934
rect 498022 102698 533786 102934
rect 534022 102698 569786 102934
rect 570022 102698 591942 102934
rect 592178 102698 592360 102934
rect -8436 102676 592360 102698
rect -8436 102674 -7836 102676
rect 29604 102674 30204 102676
rect 65604 102674 66204 102676
rect 101604 102674 102204 102676
rect 137604 102674 138204 102676
rect 173604 102674 174204 102676
rect 209604 102674 210204 102676
rect 245604 102674 246204 102676
rect 281604 102674 282204 102676
rect 317604 102674 318204 102676
rect 353604 102674 354204 102676
rect 389604 102674 390204 102676
rect 425604 102674 426204 102676
rect 461604 102674 462204 102676
rect 497604 102674 498204 102676
rect 533604 102674 534204 102676
rect 569604 102674 570204 102676
rect 591760 102674 592360 102676
rect -6596 99676 -5996 99678
rect 26004 99676 26604 99678
rect 62004 99676 62604 99678
rect 98004 99676 98604 99678
rect 134004 99676 134604 99678
rect 170004 99676 170604 99678
rect 206004 99676 206604 99678
rect 242004 99676 242604 99678
rect 278004 99676 278604 99678
rect 314004 99676 314604 99678
rect 350004 99676 350604 99678
rect 386004 99676 386604 99678
rect 422004 99676 422604 99678
rect 458004 99676 458604 99678
rect 494004 99676 494604 99678
rect 530004 99676 530604 99678
rect 566004 99676 566604 99678
rect 589920 99676 590520 99678
rect -6596 99654 590520 99676
rect -6596 99418 -6414 99654
rect -6178 99418 26186 99654
rect 26422 99418 62186 99654
rect 62422 99418 98186 99654
rect 98422 99418 134186 99654
rect 134422 99418 170186 99654
rect 170422 99418 206186 99654
rect 206422 99418 242186 99654
rect 242422 99418 278186 99654
rect 278422 99418 314186 99654
rect 314422 99418 350186 99654
rect 350422 99418 386186 99654
rect 386422 99418 422186 99654
rect 422422 99418 458186 99654
rect 458422 99418 494186 99654
rect 494422 99418 530186 99654
rect 530422 99418 566186 99654
rect 566422 99418 590102 99654
rect 590338 99418 590520 99654
rect -6596 99334 590520 99418
rect -6596 99098 -6414 99334
rect -6178 99098 26186 99334
rect 26422 99098 62186 99334
rect 62422 99098 98186 99334
rect 98422 99098 134186 99334
rect 134422 99098 170186 99334
rect 170422 99098 206186 99334
rect 206422 99098 242186 99334
rect 242422 99098 278186 99334
rect 278422 99098 314186 99334
rect 314422 99098 350186 99334
rect 350422 99098 386186 99334
rect 386422 99098 422186 99334
rect 422422 99098 458186 99334
rect 458422 99098 494186 99334
rect 494422 99098 530186 99334
rect 530422 99098 566186 99334
rect 566422 99098 590102 99334
rect 590338 99098 590520 99334
rect -6596 99076 590520 99098
rect -6596 99074 -5996 99076
rect 26004 99074 26604 99076
rect 62004 99074 62604 99076
rect 98004 99074 98604 99076
rect 134004 99074 134604 99076
rect 170004 99074 170604 99076
rect 206004 99074 206604 99076
rect 242004 99074 242604 99076
rect 278004 99074 278604 99076
rect 314004 99074 314604 99076
rect 350004 99074 350604 99076
rect 386004 99074 386604 99076
rect 422004 99074 422604 99076
rect 458004 99074 458604 99076
rect 494004 99074 494604 99076
rect 530004 99074 530604 99076
rect 566004 99074 566604 99076
rect 589920 99074 590520 99076
rect -4756 96076 -4156 96078
rect 22404 96076 23004 96078
rect 58404 96076 59004 96078
rect 94404 96076 95004 96078
rect 130404 96076 131004 96078
rect 166404 96076 167004 96078
rect 202404 96076 203004 96078
rect 238404 96076 239004 96078
rect 274404 96076 275004 96078
rect 310404 96076 311004 96078
rect 346404 96076 347004 96078
rect 382404 96076 383004 96078
rect 418404 96076 419004 96078
rect 454404 96076 455004 96078
rect 490404 96076 491004 96078
rect 526404 96076 527004 96078
rect 562404 96076 563004 96078
rect 588080 96076 588680 96078
rect -4756 96054 588680 96076
rect -4756 95818 -4574 96054
rect -4338 95818 22586 96054
rect 22822 95818 58586 96054
rect 58822 95818 94586 96054
rect 94822 95818 130586 96054
rect 130822 95818 166586 96054
rect 166822 95818 202586 96054
rect 202822 95818 238586 96054
rect 238822 95818 274586 96054
rect 274822 95818 310586 96054
rect 310822 95818 346586 96054
rect 346822 95818 382586 96054
rect 382822 95818 418586 96054
rect 418822 95818 454586 96054
rect 454822 95818 490586 96054
rect 490822 95818 526586 96054
rect 526822 95818 562586 96054
rect 562822 95818 588262 96054
rect 588498 95818 588680 96054
rect -4756 95734 588680 95818
rect -4756 95498 -4574 95734
rect -4338 95498 22586 95734
rect 22822 95498 58586 95734
rect 58822 95498 94586 95734
rect 94822 95498 130586 95734
rect 130822 95498 166586 95734
rect 166822 95498 202586 95734
rect 202822 95498 238586 95734
rect 238822 95498 274586 95734
rect 274822 95498 310586 95734
rect 310822 95498 346586 95734
rect 346822 95498 382586 95734
rect 382822 95498 418586 95734
rect 418822 95498 454586 95734
rect 454822 95498 490586 95734
rect 490822 95498 526586 95734
rect 526822 95498 562586 95734
rect 562822 95498 588262 95734
rect 588498 95498 588680 95734
rect -4756 95476 588680 95498
rect -4756 95474 -4156 95476
rect 22404 95474 23004 95476
rect 58404 95474 59004 95476
rect 94404 95474 95004 95476
rect 130404 95474 131004 95476
rect 166404 95474 167004 95476
rect 202404 95474 203004 95476
rect 238404 95474 239004 95476
rect 274404 95474 275004 95476
rect 310404 95474 311004 95476
rect 346404 95474 347004 95476
rect 382404 95474 383004 95476
rect 418404 95474 419004 95476
rect 454404 95474 455004 95476
rect 490404 95474 491004 95476
rect 526404 95474 527004 95476
rect 562404 95474 563004 95476
rect 588080 95474 588680 95476
rect -2916 92476 -2316 92478
rect 18804 92476 19404 92478
rect 54804 92476 55404 92478
rect 90804 92476 91404 92478
rect 126804 92476 127404 92478
rect 162804 92476 163404 92478
rect 198804 92476 199404 92478
rect 234804 92476 235404 92478
rect 270804 92476 271404 92478
rect 306804 92476 307404 92478
rect 342804 92476 343404 92478
rect 378804 92476 379404 92478
rect 414804 92476 415404 92478
rect 450804 92476 451404 92478
rect 486804 92476 487404 92478
rect 522804 92476 523404 92478
rect 558804 92476 559404 92478
rect 586240 92476 586840 92478
rect -2916 92454 586840 92476
rect -2916 92218 -2734 92454
rect -2498 92218 18986 92454
rect 19222 92218 54986 92454
rect 55222 92218 90986 92454
rect 91222 92218 126986 92454
rect 127222 92218 162986 92454
rect 163222 92218 198986 92454
rect 199222 92218 234986 92454
rect 235222 92218 270986 92454
rect 271222 92218 306986 92454
rect 307222 92218 342986 92454
rect 343222 92218 378986 92454
rect 379222 92218 414986 92454
rect 415222 92218 450986 92454
rect 451222 92218 486986 92454
rect 487222 92218 522986 92454
rect 523222 92218 558986 92454
rect 559222 92218 586422 92454
rect 586658 92218 586840 92454
rect -2916 92134 586840 92218
rect -2916 91898 -2734 92134
rect -2498 91898 18986 92134
rect 19222 91898 54986 92134
rect 55222 91898 90986 92134
rect 91222 91898 126986 92134
rect 127222 91898 162986 92134
rect 163222 91898 198986 92134
rect 199222 91898 234986 92134
rect 235222 91898 270986 92134
rect 271222 91898 306986 92134
rect 307222 91898 342986 92134
rect 343222 91898 378986 92134
rect 379222 91898 414986 92134
rect 415222 91898 450986 92134
rect 451222 91898 486986 92134
rect 487222 91898 522986 92134
rect 523222 91898 558986 92134
rect 559222 91898 586422 92134
rect 586658 91898 586840 92134
rect -2916 91876 586840 91898
rect -2916 91874 -2316 91876
rect 18804 91874 19404 91876
rect 54804 91874 55404 91876
rect 90804 91874 91404 91876
rect 126804 91874 127404 91876
rect 162804 91874 163404 91876
rect 198804 91874 199404 91876
rect 234804 91874 235404 91876
rect 270804 91874 271404 91876
rect 306804 91874 307404 91876
rect 342804 91874 343404 91876
rect 378804 91874 379404 91876
rect 414804 91874 415404 91876
rect 450804 91874 451404 91876
rect 486804 91874 487404 91876
rect 522804 91874 523404 91876
rect 558804 91874 559404 91876
rect 586240 91874 586840 91876
rect -7516 85276 -6916 85278
rect 11604 85276 12204 85278
rect 47604 85276 48204 85278
rect 83604 85276 84204 85278
rect 119604 85276 120204 85278
rect 155604 85276 156204 85278
rect 191604 85276 192204 85278
rect 227604 85276 228204 85278
rect 263604 85276 264204 85278
rect 299604 85276 300204 85278
rect 335604 85276 336204 85278
rect 371604 85276 372204 85278
rect 407604 85276 408204 85278
rect 443604 85276 444204 85278
rect 479604 85276 480204 85278
rect 515604 85276 516204 85278
rect 551604 85276 552204 85278
rect 590840 85276 591440 85278
rect -8436 85254 592360 85276
rect -8436 85018 -7334 85254
rect -7098 85018 11786 85254
rect 12022 85018 47786 85254
rect 48022 85018 83786 85254
rect 84022 85018 119786 85254
rect 120022 85018 155786 85254
rect 156022 85018 191786 85254
rect 192022 85018 227786 85254
rect 228022 85018 263786 85254
rect 264022 85018 299786 85254
rect 300022 85018 335786 85254
rect 336022 85018 371786 85254
rect 372022 85018 407786 85254
rect 408022 85018 443786 85254
rect 444022 85018 479786 85254
rect 480022 85018 515786 85254
rect 516022 85018 551786 85254
rect 552022 85018 591022 85254
rect 591258 85018 592360 85254
rect -8436 84934 592360 85018
rect -8436 84698 -7334 84934
rect -7098 84698 11786 84934
rect 12022 84698 47786 84934
rect 48022 84698 83786 84934
rect 84022 84698 119786 84934
rect 120022 84698 155786 84934
rect 156022 84698 191786 84934
rect 192022 84698 227786 84934
rect 228022 84698 263786 84934
rect 264022 84698 299786 84934
rect 300022 84698 335786 84934
rect 336022 84698 371786 84934
rect 372022 84698 407786 84934
rect 408022 84698 443786 84934
rect 444022 84698 479786 84934
rect 480022 84698 515786 84934
rect 516022 84698 551786 84934
rect 552022 84698 591022 84934
rect 591258 84698 592360 84934
rect -8436 84676 592360 84698
rect -7516 84674 -6916 84676
rect 11604 84674 12204 84676
rect 47604 84674 48204 84676
rect 83604 84674 84204 84676
rect 119604 84674 120204 84676
rect 155604 84674 156204 84676
rect 191604 84674 192204 84676
rect 227604 84674 228204 84676
rect 263604 84674 264204 84676
rect 299604 84674 300204 84676
rect 335604 84674 336204 84676
rect 371604 84674 372204 84676
rect 407604 84674 408204 84676
rect 443604 84674 444204 84676
rect 479604 84674 480204 84676
rect 515604 84674 516204 84676
rect 551604 84674 552204 84676
rect 590840 84674 591440 84676
rect -5676 81676 -5076 81678
rect 8004 81676 8604 81678
rect 44004 81676 44604 81678
rect 80004 81676 80604 81678
rect 116004 81676 116604 81678
rect 152004 81676 152604 81678
rect 188004 81676 188604 81678
rect 224004 81676 224604 81678
rect 260004 81676 260604 81678
rect 296004 81676 296604 81678
rect 332004 81676 332604 81678
rect 368004 81676 368604 81678
rect 404004 81676 404604 81678
rect 440004 81676 440604 81678
rect 476004 81676 476604 81678
rect 512004 81676 512604 81678
rect 548004 81676 548604 81678
rect 589000 81676 589600 81678
rect -6596 81654 590520 81676
rect -6596 81418 -5494 81654
rect -5258 81418 8186 81654
rect 8422 81418 44186 81654
rect 44422 81418 80186 81654
rect 80422 81418 116186 81654
rect 116422 81418 152186 81654
rect 152422 81418 188186 81654
rect 188422 81418 224186 81654
rect 224422 81418 260186 81654
rect 260422 81418 296186 81654
rect 296422 81418 332186 81654
rect 332422 81418 368186 81654
rect 368422 81418 404186 81654
rect 404422 81418 440186 81654
rect 440422 81418 476186 81654
rect 476422 81418 512186 81654
rect 512422 81418 548186 81654
rect 548422 81418 589182 81654
rect 589418 81418 590520 81654
rect -6596 81334 590520 81418
rect -6596 81098 -5494 81334
rect -5258 81098 8186 81334
rect 8422 81098 44186 81334
rect 44422 81098 80186 81334
rect 80422 81098 116186 81334
rect 116422 81098 152186 81334
rect 152422 81098 188186 81334
rect 188422 81098 224186 81334
rect 224422 81098 260186 81334
rect 260422 81098 296186 81334
rect 296422 81098 332186 81334
rect 332422 81098 368186 81334
rect 368422 81098 404186 81334
rect 404422 81098 440186 81334
rect 440422 81098 476186 81334
rect 476422 81098 512186 81334
rect 512422 81098 548186 81334
rect 548422 81098 589182 81334
rect 589418 81098 590520 81334
rect -6596 81076 590520 81098
rect -5676 81074 -5076 81076
rect 8004 81074 8604 81076
rect 44004 81074 44604 81076
rect 80004 81074 80604 81076
rect 116004 81074 116604 81076
rect 152004 81074 152604 81076
rect 188004 81074 188604 81076
rect 224004 81074 224604 81076
rect 260004 81074 260604 81076
rect 296004 81074 296604 81076
rect 332004 81074 332604 81076
rect 368004 81074 368604 81076
rect 404004 81074 404604 81076
rect 440004 81074 440604 81076
rect 476004 81074 476604 81076
rect 512004 81074 512604 81076
rect 548004 81074 548604 81076
rect 589000 81074 589600 81076
rect -3836 78076 -3236 78078
rect 4404 78076 5004 78078
rect 40404 78076 41004 78078
rect 76404 78076 77004 78078
rect 112404 78076 113004 78078
rect 148404 78076 149004 78078
rect 184404 78076 185004 78078
rect 220404 78076 221004 78078
rect 256404 78076 257004 78078
rect 292404 78076 293004 78078
rect 328404 78076 329004 78078
rect 364404 78076 365004 78078
rect 400404 78076 401004 78078
rect 436404 78076 437004 78078
rect 472404 78076 473004 78078
rect 508404 78076 509004 78078
rect 544404 78076 545004 78078
rect 580404 78076 581004 78078
rect 587160 78076 587760 78078
rect -4756 78054 588680 78076
rect -4756 77818 -3654 78054
rect -3418 77818 4586 78054
rect 4822 77818 40586 78054
rect 40822 77818 76586 78054
rect 76822 77818 112586 78054
rect 112822 77818 148586 78054
rect 148822 77818 184586 78054
rect 184822 77818 220586 78054
rect 220822 77818 256586 78054
rect 256822 77818 292586 78054
rect 292822 77818 328586 78054
rect 328822 77818 364586 78054
rect 364822 77818 400586 78054
rect 400822 77818 436586 78054
rect 436822 77818 472586 78054
rect 472822 77818 508586 78054
rect 508822 77818 544586 78054
rect 544822 77818 580586 78054
rect 580822 77818 587342 78054
rect 587578 77818 588680 78054
rect -4756 77734 588680 77818
rect -4756 77498 -3654 77734
rect -3418 77498 4586 77734
rect 4822 77498 40586 77734
rect 40822 77498 76586 77734
rect 76822 77498 112586 77734
rect 112822 77498 148586 77734
rect 148822 77498 184586 77734
rect 184822 77498 220586 77734
rect 220822 77498 256586 77734
rect 256822 77498 292586 77734
rect 292822 77498 328586 77734
rect 328822 77498 364586 77734
rect 364822 77498 400586 77734
rect 400822 77498 436586 77734
rect 436822 77498 472586 77734
rect 472822 77498 508586 77734
rect 508822 77498 544586 77734
rect 544822 77498 580586 77734
rect 580822 77498 587342 77734
rect 587578 77498 588680 77734
rect -4756 77476 588680 77498
rect -3836 77474 -3236 77476
rect 4404 77474 5004 77476
rect 40404 77474 41004 77476
rect 76404 77474 77004 77476
rect 112404 77474 113004 77476
rect 148404 77474 149004 77476
rect 184404 77474 185004 77476
rect 220404 77474 221004 77476
rect 256404 77474 257004 77476
rect 292404 77474 293004 77476
rect 328404 77474 329004 77476
rect 364404 77474 365004 77476
rect 400404 77474 401004 77476
rect 436404 77474 437004 77476
rect 472404 77474 473004 77476
rect 508404 77474 509004 77476
rect 544404 77474 545004 77476
rect 580404 77474 581004 77476
rect 587160 77474 587760 77476
rect -1996 74476 -1396 74478
rect 804 74476 1404 74478
rect 36804 74476 37404 74478
rect 72804 74476 73404 74478
rect 108804 74476 109404 74478
rect 144804 74476 145404 74478
rect 180804 74476 181404 74478
rect 216804 74476 217404 74478
rect 252804 74476 253404 74478
rect 288804 74476 289404 74478
rect 324804 74476 325404 74478
rect 360804 74476 361404 74478
rect 396804 74476 397404 74478
rect 432804 74476 433404 74478
rect 468804 74476 469404 74478
rect 504804 74476 505404 74478
rect 540804 74476 541404 74478
rect 576804 74476 577404 74478
rect 585320 74476 585920 74478
rect -2916 74454 586840 74476
rect -2916 74218 -1814 74454
rect -1578 74218 986 74454
rect 1222 74218 36986 74454
rect 37222 74218 72986 74454
rect 73222 74218 108986 74454
rect 109222 74218 144986 74454
rect 145222 74218 180986 74454
rect 181222 74218 216986 74454
rect 217222 74218 252986 74454
rect 253222 74218 288986 74454
rect 289222 74218 324986 74454
rect 325222 74218 360986 74454
rect 361222 74218 396986 74454
rect 397222 74218 432986 74454
rect 433222 74218 468986 74454
rect 469222 74218 504986 74454
rect 505222 74218 540986 74454
rect 541222 74218 576986 74454
rect 577222 74218 585502 74454
rect 585738 74218 586840 74454
rect -2916 74134 586840 74218
rect -2916 73898 -1814 74134
rect -1578 73898 986 74134
rect 1222 73898 36986 74134
rect 37222 73898 72986 74134
rect 73222 73898 108986 74134
rect 109222 73898 144986 74134
rect 145222 73898 180986 74134
rect 181222 73898 216986 74134
rect 217222 73898 252986 74134
rect 253222 73898 288986 74134
rect 289222 73898 324986 74134
rect 325222 73898 360986 74134
rect 361222 73898 396986 74134
rect 397222 73898 432986 74134
rect 433222 73898 468986 74134
rect 469222 73898 504986 74134
rect 505222 73898 540986 74134
rect 541222 73898 576986 74134
rect 577222 73898 585502 74134
rect 585738 73898 586840 74134
rect -2916 73876 586840 73898
rect -1996 73874 -1396 73876
rect 804 73874 1404 73876
rect 36804 73874 37404 73876
rect 72804 73874 73404 73876
rect 108804 73874 109404 73876
rect 144804 73874 145404 73876
rect 180804 73874 181404 73876
rect 216804 73874 217404 73876
rect 252804 73874 253404 73876
rect 288804 73874 289404 73876
rect 324804 73874 325404 73876
rect 360804 73874 361404 73876
rect 396804 73874 397404 73876
rect 432804 73874 433404 73876
rect 468804 73874 469404 73876
rect 504804 73874 505404 73876
rect 540804 73874 541404 73876
rect 576804 73874 577404 73876
rect 585320 73874 585920 73876
rect -8436 67276 -7836 67278
rect 29604 67276 30204 67278
rect 65604 67276 66204 67278
rect 101604 67276 102204 67278
rect 137604 67276 138204 67278
rect 173604 67276 174204 67278
rect 209604 67276 210204 67278
rect 245604 67276 246204 67278
rect 281604 67276 282204 67278
rect 317604 67276 318204 67278
rect 353604 67276 354204 67278
rect 389604 67276 390204 67278
rect 425604 67276 426204 67278
rect 461604 67276 462204 67278
rect 497604 67276 498204 67278
rect 533604 67276 534204 67278
rect 569604 67276 570204 67278
rect 591760 67276 592360 67278
rect -8436 67254 592360 67276
rect -8436 67018 -8254 67254
rect -8018 67018 29786 67254
rect 30022 67018 65786 67254
rect 66022 67018 101786 67254
rect 102022 67018 137786 67254
rect 138022 67018 173786 67254
rect 174022 67018 209786 67254
rect 210022 67018 245786 67254
rect 246022 67018 281786 67254
rect 282022 67018 317786 67254
rect 318022 67018 353786 67254
rect 354022 67018 389786 67254
rect 390022 67018 425786 67254
rect 426022 67018 461786 67254
rect 462022 67018 497786 67254
rect 498022 67018 533786 67254
rect 534022 67018 569786 67254
rect 570022 67018 591942 67254
rect 592178 67018 592360 67254
rect -8436 66934 592360 67018
rect -8436 66698 -8254 66934
rect -8018 66698 29786 66934
rect 30022 66698 65786 66934
rect 66022 66698 101786 66934
rect 102022 66698 137786 66934
rect 138022 66698 173786 66934
rect 174022 66698 209786 66934
rect 210022 66698 245786 66934
rect 246022 66698 281786 66934
rect 282022 66698 317786 66934
rect 318022 66698 353786 66934
rect 354022 66698 389786 66934
rect 390022 66698 425786 66934
rect 426022 66698 461786 66934
rect 462022 66698 497786 66934
rect 498022 66698 533786 66934
rect 534022 66698 569786 66934
rect 570022 66698 591942 66934
rect 592178 66698 592360 66934
rect -8436 66676 592360 66698
rect -8436 66674 -7836 66676
rect 29604 66674 30204 66676
rect 65604 66674 66204 66676
rect 101604 66674 102204 66676
rect 137604 66674 138204 66676
rect 173604 66674 174204 66676
rect 209604 66674 210204 66676
rect 245604 66674 246204 66676
rect 281604 66674 282204 66676
rect 317604 66674 318204 66676
rect 353604 66674 354204 66676
rect 389604 66674 390204 66676
rect 425604 66674 426204 66676
rect 461604 66674 462204 66676
rect 497604 66674 498204 66676
rect 533604 66674 534204 66676
rect 569604 66674 570204 66676
rect 591760 66674 592360 66676
rect -6596 63676 -5996 63678
rect 26004 63676 26604 63678
rect 62004 63676 62604 63678
rect 98004 63676 98604 63678
rect 134004 63676 134604 63678
rect 170004 63676 170604 63678
rect 206004 63676 206604 63678
rect 242004 63676 242604 63678
rect 278004 63676 278604 63678
rect 314004 63676 314604 63678
rect 350004 63676 350604 63678
rect 386004 63676 386604 63678
rect 422004 63676 422604 63678
rect 458004 63676 458604 63678
rect 494004 63676 494604 63678
rect 530004 63676 530604 63678
rect 566004 63676 566604 63678
rect 589920 63676 590520 63678
rect -6596 63654 590520 63676
rect -6596 63418 -6414 63654
rect -6178 63418 26186 63654
rect 26422 63418 62186 63654
rect 62422 63418 98186 63654
rect 98422 63418 134186 63654
rect 134422 63418 170186 63654
rect 170422 63418 206186 63654
rect 206422 63418 242186 63654
rect 242422 63418 278186 63654
rect 278422 63418 314186 63654
rect 314422 63418 350186 63654
rect 350422 63418 386186 63654
rect 386422 63418 422186 63654
rect 422422 63418 458186 63654
rect 458422 63418 494186 63654
rect 494422 63418 530186 63654
rect 530422 63418 566186 63654
rect 566422 63418 590102 63654
rect 590338 63418 590520 63654
rect -6596 63334 590520 63418
rect -6596 63098 -6414 63334
rect -6178 63098 26186 63334
rect 26422 63098 62186 63334
rect 62422 63098 98186 63334
rect 98422 63098 134186 63334
rect 134422 63098 170186 63334
rect 170422 63098 206186 63334
rect 206422 63098 242186 63334
rect 242422 63098 278186 63334
rect 278422 63098 314186 63334
rect 314422 63098 350186 63334
rect 350422 63098 386186 63334
rect 386422 63098 422186 63334
rect 422422 63098 458186 63334
rect 458422 63098 494186 63334
rect 494422 63098 530186 63334
rect 530422 63098 566186 63334
rect 566422 63098 590102 63334
rect 590338 63098 590520 63334
rect -6596 63076 590520 63098
rect -6596 63074 -5996 63076
rect 26004 63074 26604 63076
rect 62004 63074 62604 63076
rect 98004 63074 98604 63076
rect 134004 63074 134604 63076
rect 170004 63074 170604 63076
rect 206004 63074 206604 63076
rect 242004 63074 242604 63076
rect 278004 63074 278604 63076
rect 314004 63074 314604 63076
rect 350004 63074 350604 63076
rect 386004 63074 386604 63076
rect 422004 63074 422604 63076
rect 458004 63074 458604 63076
rect 494004 63074 494604 63076
rect 530004 63074 530604 63076
rect 566004 63074 566604 63076
rect 589920 63074 590520 63076
rect -4756 60076 -4156 60078
rect 22404 60076 23004 60078
rect 58404 60076 59004 60078
rect 94404 60076 95004 60078
rect 130404 60076 131004 60078
rect 166404 60076 167004 60078
rect 202404 60076 203004 60078
rect 238404 60076 239004 60078
rect 274404 60076 275004 60078
rect 310404 60076 311004 60078
rect 346404 60076 347004 60078
rect 382404 60076 383004 60078
rect 418404 60076 419004 60078
rect 454404 60076 455004 60078
rect 490404 60076 491004 60078
rect 526404 60076 527004 60078
rect 562404 60076 563004 60078
rect 588080 60076 588680 60078
rect -4756 60054 588680 60076
rect -4756 59818 -4574 60054
rect -4338 59818 22586 60054
rect 22822 59818 58586 60054
rect 58822 59818 94586 60054
rect 94822 59818 130586 60054
rect 130822 59818 166586 60054
rect 166822 59818 202586 60054
rect 202822 59818 238586 60054
rect 238822 59818 274586 60054
rect 274822 59818 310586 60054
rect 310822 59818 346586 60054
rect 346822 59818 382586 60054
rect 382822 59818 418586 60054
rect 418822 59818 454586 60054
rect 454822 59818 490586 60054
rect 490822 59818 526586 60054
rect 526822 59818 562586 60054
rect 562822 59818 588262 60054
rect 588498 59818 588680 60054
rect -4756 59734 588680 59818
rect -4756 59498 -4574 59734
rect -4338 59498 22586 59734
rect 22822 59498 58586 59734
rect 58822 59498 94586 59734
rect 94822 59498 130586 59734
rect 130822 59498 166586 59734
rect 166822 59498 202586 59734
rect 202822 59498 238586 59734
rect 238822 59498 274586 59734
rect 274822 59498 310586 59734
rect 310822 59498 346586 59734
rect 346822 59498 382586 59734
rect 382822 59498 418586 59734
rect 418822 59498 454586 59734
rect 454822 59498 490586 59734
rect 490822 59498 526586 59734
rect 526822 59498 562586 59734
rect 562822 59498 588262 59734
rect 588498 59498 588680 59734
rect -4756 59476 588680 59498
rect -4756 59474 -4156 59476
rect 22404 59474 23004 59476
rect 58404 59474 59004 59476
rect 94404 59474 95004 59476
rect 130404 59474 131004 59476
rect 166404 59474 167004 59476
rect 202404 59474 203004 59476
rect 238404 59474 239004 59476
rect 274404 59474 275004 59476
rect 310404 59474 311004 59476
rect 346404 59474 347004 59476
rect 382404 59474 383004 59476
rect 418404 59474 419004 59476
rect 454404 59474 455004 59476
rect 490404 59474 491004 59476
rect 526404 59474 527004 59476
rect 562404 59474 563004 59476
rect 588080 59474 588680 59476
rect -2916 56476 -2316 56478
rect 18804 56476 19404 56478
rect 54804 56476 55404 56478
rect 90804 56476 91404 56478
rect 126804 56476 127404 56478
rect 162804 56476 163404 56478
rect 198804 56476 199404 56478
rect 234804 56476 235404 56478
rect 270804 56476 271404 56478
rect 306804 56476 307404 56478
rect 342804 56476 343404 56478
rect 378804 56476 379404 56478
rect 414804 56476 415404 56478
rect 450804 56476 451404 56478
rect 486804 56476 487404 56478
rect 522804 56476 523404 56478
rect 558804 56476 559404 56478
rect 586240 56476 586840 56478
rect -2916 56454 586840 56476
rect -2916 56218 -2734 56454
rect -2498 56218 18986 56454
rect 19222 56218 54986 56454
rect 55222 56218 90986 56454
rect 91222 56218 126986 56454
rect 127222 56218 162986 56454
rect 163222 56218 198986 56454
rect 199222 56218 234986 56454
rect 235222 56218 270986 56454
rect 271222 56218 306986 56454
rect 307222 56218 342986 56454
rect 343222 56218 378986 56454
rect 379222 56218 414986 56454
rect 415222 56218 450986 56454
rect 451222 56218 486986 56454
rect 487222 56218 522986 56454
rect 523222 56218 558986 56454
rect 559222 56218 586422 56454
rect 586658 56218 586840 56454
rect -2916 56134 586840 56218
rect -2916 55898 -2734 56134
rect -2498 55898 18986 56134
rect 19222 55898 54986 56134
rect 55222 55898 90986 56134
rect 91222 55898 126986 56134
rect 127222 55898 162986 56134
rect 163222 55898 198986 56134
rect 199222 55898 234986 56134
rect 235222 55898 270986 56134
rect 271222 55898 306986 56134
rect 307222 55898 342986 56134
rect 343222 55898 378986 56134
rect 379222 55898 414986 56134
rect 415222 55898 450986 56134
rect 451222 55898 486986 56134
rect 487222 55898 522986 56134
rect 523222 55898 558986 56134
rect 559222 55898 586422 56134
rect 586658 55898 586840 56134
rect -2916 55876 586840 55898
rect -2916 55874 -2316 55876
rect 18804 55874 19404 55876
rect 54804 55874 55404 55876
rect 90804 55874 91404 55876
rect 126804 55874 127404 55876
rect 162804 55874 163404 55876
rect 198804 55874 199404 55876
rect 234804 55874 235404 55876
rect 270804 55874 271404 55876
rect 306804 55874 307404 55876
rect 342804 55874 343404 55876
rect 378804 55874 379404 55876
rect 414804 55874 415404 55876
rect 450804 55874 451404 55876
rect 486804 55874 487404 55876
rect 522804 55874 523404 55876
rect 558804 55874 559404 55876
rect 586240 55874 586840 55876
rect -7516 49276 -6916 49278
rect 11604 49276 12204 49278
rect 47604 49276 48204 49278
rect 83604 49276 84204 49278
rect 119604 49276 120204 49278
rect 155604 49276 156204 49278
rect 191604 49276 192204 49278
rect 227604 49276 228204 49278
rect 263604 49276 264204 49278
rect 299604 49276 300204 49278
rect 335604 49276 336204 49278
rect 371604 49276 372204 49278
rect 407604 49276 408204 49278
rect 443604 49276 444204 49278
rect 479604 49276 480204 49278
rect 515604 49276 516204 49278
rect 551604 49276 552204 49278
rect 590840 49276 591440 49278
rect -8436 49254 592360 49276
rect -8436 49018 -7334 49254
rect -7098 49018 11786 49254
rect 12022 49018 47786 49254
rect 48022 49018 83786 49254
rect 84022 49018 119786 49254
rect 120022 49018 155786 49254
rect 156022 49018 191786 49254
rect 192022 49018 227786 49254
rect 228022 49018 263786 49254
rect 264022 49018 299786 49254
rect 300022 49018 335786 49254
rect 336022 49018 371786 49254
rect 372022 49018 407786 49254
rect 408022 49018 443786 49254
rect 444022 49018 479786 49254
rect 480022 49018 515786 49254
rect 516022 49018 551786 49254
rect 552022 49018 591022 49254
rect 591258 49018 592360 49254
rect -8436 48934 592360 49018
rect -8436 48698 -7334 48934
rect -7098 48698 11786 48934
rect 12022 48698 47786 48934
rect 48022 48698 83786 48934
rect 84022 48698 119786 48934
rect 120022 48698 155786 48934
rect 156022 48698 191786 48934
rect 192022 48698 227786 48934
rect 228022 48698 263786 48934
rect 264022 48698 299786 48934
rect 300022 48698 335786 48934
rect 336022 48698 371786 48934
rect 372022 48698 407786 48934
rect 408022 48698 443786 48934
rect 444022 48698 479786 48934
rect 480022 48698 515786 48934
rect 516022 48698 551786 48934
rect 552022 48698 591022 48934
rect 591258 48698 592360 48934
rect -8436 48676 592360 48698
rect -7516 48674 -6916 48676
rect 11604 48674 12204 48676
rect 47604 48674 48204 48676
rect 83604 48674 84204 48676
rect 119604 48674 120204 48676
rect 155604 48674 156204 48676
rect 191604 48674 192204 48676
rect 227604 48674 228204 48676
rect 263604 48674 264204 48676
rect 299604 48674 300204 48676
rect 335604 48674 336204 48676
rect 371604 48674 372204 48676
rect 407604 48674 408204 48676
rect 443604 48674 444204 48676
rect 479604 48674 480204 48676
rect 515604 48674 516204 48676
rect 551604 48674 552204 48676
rect 590840 48674 591440 48676
rect -5676 45676 -5076 45678
rect 8004 45676 8604 45678
rect 44004 45676 44604 45678
rect 80004 45676 80604 45678
rect 116004 45676 116604 45678
rect 152004 45676 152604 45678
rect 188004 45676 188604 45678
rect 224004 45676 224604 45678
rect 260004 45676 260604 45678
rect 296004 45676 296604 45678
rect 332004 45676 332604 45678
rect 368004 45676 368604 45678
rect 404004 45676 404604 45678
rect 440004 45676 440604 45678
rect 476004 45676 476604 45678
rect 512004 45676 512604 45678
rect 548004 45676 548604 45678
rect 589000 45676 589600 45678
rect -6596 45654 590520 45676
rect -6596 45418 -5494 45654
rect -5258 45418 8186 45654
rect 8422 45418 44186 45654
rect 44422 45418 80186 45654
rect 80422 45418 116186 45654
rect 116422 45418 152186 45654
rect 152422 45418 188186 45654
rect 188422 45418 224186 45654
rect 224422 45418 260186 45654
rect 260422 45418 296186 45654
rect 296422 45418 332186 45654
rect 332422 45418 368186 45654
rect 368422 45418 404186 45654
rect 404422 45418 440186 45654
rect 440422 45418 476186 45654
rect 476422 45418 512186 45654
rect 512422 45418 548186 45654
rect 548422 45418 589182 45654
rect 589418 45418 590520 45654
rect -6596 45334 590520 45418
rect -6596 45098 -5494 45334
rect -5258 45098 8186 45334
rect 8422 45098 44186 45334
rect 44422 45098 80186 45334
rect 80422 45098 116186 45334
rect 116422 45098 152186 45334
rect 152422 45098 188186 45334
rect 188422 45098 224186 45334
rect 224422 45098 260186 45334
rect 260422 45098 296186 45334
rect 296422 45098 332186 45334
rect 332422 45098 368186 45334
rect 368422 45098 404186 45334
rect 404422 45098 440186 45334
rect 440422 45098 476186 45334
rect 476422 45098 512186 45334
rect 512422 45098 548186 45334
rect 548422 45098 589182 45334
rect 589418 45098 590520 45334
rect -6596 45076 590520 45098
rect -5676 45074 -5076 45076
rect 8004 45074 8604 45076
rect 44004 45074 44604 45076
rect 80004 45074 80604 45076
rect 116004 45074 116604 45076
rect 152004 45074 152604 45076
rect 188004 45074 188604 45076
rect 224004 45074 224604 45076
rect 260004 45074 260604 45076
rect 296004 45074 296604 45076
rect 332004 45074 332604 45076
rect 368004 45074 368604 45076
rect 404004 45074 404604 45076
rect 440004 45074 440604 45076
rect 476004 45074 476604 45076
rect 512004 45074 512604 45076
rect 548004 45074 548604 45076
rect 589000 45074 589600 45076
rect -3836 42076 -3236 42078
rect 4404 42076 5004 42078
rect 40404 42076 41004 42078
rect 76404 42076 77004 42078
rect 112404 42076 113004 42078
rect 148404 42076 149004 42078
rect 184404 42076 185004 42078
rect 220404 42076 221004 42078
rect 256404 42076 257004 42078
rect 292404 42076 293004 42078
rect 328404 42076 329004 42078
rect 364404 42076 365004 42078
rect 400404 42076 401004 42078
rect 436404 42076 437004 42078
rect 472404 42076 473004 42078
rect 508404 42076 509004 42078
rect 544404 42076 545004 42078
rect 580404 42076 581004 42078
rect 587160 42076 587760 42078
rect -4756 42054 588680 42076
rect -4756 41818 -3654 42054
rect -3418 41818 4586 42054
rect 4822 41818 40586 42054
rect 40822 41818 76586 42054
rect 76822 41818 112586 42054
rect 112822 41818 148586 42054
rect 148822 41818 184586 42054
rect 184822 41818 220586 42054
rect 220822 41818 256586 42054
rect 256822 41818 292586 42054
rect 292822 41818 328586 42054
rect 328822 41818 364586 42054
rect 364822 41818 400586 42054
rect 400822 41818 436586 42054
rect 436822 41818 472586 42054
rect 472822 41818 508586 42054
rect 508822 41818 544586 42054
rect 544822 41818 580586 42054
rect 580822 41818 587342 42054
rect 587578 41818 588680 42054
rect -4756 41734 588680 41818
rect -4756 41498 -3654 41734
rect -3418 41498 4586 41734
rect 4822 41498 40586 41734
rect 40822 41498 76586 41734
rect 76822 41498 112586 41734
rect 112822 41498 148586 41734
rect 148822 41498 184586 41734
rect 184822 41498 220586 41734
rect 220822 41498 256586 41734
rect 256822 41498 292586 41734
rect 292822 41498 328586 41734
rect 328822 41498 364586 41734
rect 364822 41498 400586 41734
rect 400822 41498 436586 41734
rect 436822 41498 472586 41734
rect 472822 41498 508586 41734
rect 508822 41498 544586 41734
rect 544822 41498 580586 41734
rect 580822 41498 587342 41734
rect 587578 41498 588680 41734
rect -4756 41476 588680 41498
rect -3836 41474 -3236 41476
rect 4404 41474 5004 41476
rect 40404 41474 41004 41476
rect 76404 41474 77004 41476
rect 112404 41474 113004 41476
rect 148404 41474 149004 41476
rect 184404 41474 185004 41476
rect 220404 41474 221004 41476
rect 256404 41474 257004 41476
rect 292404 41474 293004 41476
rect 328404 41474 329004 41476
rect 364404 41474 365004 41476
rect 400404 41474 401004 41476
rect 436404 41474 437004 41476
rect 472404 41474 473004 41476
rect 508404 41474 509004 41476
rect 544404 41474 545004 41476
rect 580404 41474 581004 41476
rect 587160 41474 587760 41476
rect -1996 38476 -1396 38478
rect 804 38476 1404 38478
rect 36804 38476 37404 38478
rect 72804 38476 73404 38478
rect 108804 38476 109404 38478
rect 144804 38476 145404 38478
rect 180804 38476 181404 38478
rect 216804 38476 217404 38478
rect 252804 38476 253404 38478
rect 288804 38476 289404 38478
rect 324804 38476 325404 38478
rect 360804 38476 361404 38478
rect 396804 38476 397404 38478
rect 432804 38476 433404 38478
rect 468804 38476 469404 38478
rect 504804 38476 505404 38478
rect 540804 38476 541404 38478
rect 576804 38476 577404 38478
rect 585320 38476 585920 38478
rect -2916 38454 586840 38476
rect -2916 38218 -1814 38454
rect -1578 38218 986 38454
rect 1222 38218 36986 38454
rect 37222 38218 72986 38454
rect 73222 38218 108986 38454
rect 109222 38218 144986 38454
rect 145222 38218 180986 38454
rect 181222 38218 216986 38454
rect 217222 38218 252986 38454
rect 253222 38218 288986 38454
rect 289222 38218 324986 38454
rect 325222 38218 360986 38454
rect 361222 38218 396986 38454
rect 397222 38218 432986 38454
rect 433222 38218 468986 38454
rect 469222 38218 504986 38454
rect 505222 38218 540986 38454
rect 541222 38218 576986 38454
rect 577222 38218 585502 38454
rect 585738 38218 586840 38454
rect -2916 38134 586840 38218
rect -2916 37898 -1814 38134
rect -1578 37898 986 38134
rect 1222 37898 36986 38134
rect 37222 37898 72986 38134
rect 73222 37898 108986 38134
rect 109222 37898 144986 38134
rect 145222 37898 180986 38134
rect 181222 37898 216986 38134
rect 217222 37898 252986 38134
rect 253222 37898 288986 38134
rect 289222 37898 324986 38134
rect 325222 37898 360986 38134
rect 361222 37898 396986 38134
rect 397222 37898 432986 38134
rect 433222 37898 468986 38134
rect 469222 37898 504986 38134
rect 505222 37898 540986 38134
rect 541222 37898 576986 38134
rect 577222 37898 585502 38134
rect 585738 37898 586840 38134
rect -2916 37876 586840 37898
rect -1996 37874 -1396 37876
rect 804 37874 1404 37876
rect 36804 37874 37404 37876
rect 72804 37874 73404 37876
rect 108804 37874 109404 37876
rect 144804 37874 145404 37876
rect 180804 37874 181404 37876
rect 216804 37874 217404 37876
rect 252804 37874 253404 37876
rect 288804 37874 289404 37876
rect 324804 37874 325404 37876
rect 360804 37874 361404 37876
rect 396804 37874 397404 37876
rect 432804 37874 433404 37876
rect 468804 37874 469404 37876
rect 504804 37874 505404 37876
rect 540804 37874 541404 37876
rect 576804 37874 577404 37876
rect 585320 37874 585920 37876
rect -8436 31276 -7836 31278
rect 29604 31276 30204 31278
rect 65604 31276 66204 31278
rect 101604 31276 102204 31278
rect 137604 31276 138204 31278
rect 173604 31276 174204 31278
rect 209604 31276 210204 31278
rect 245604 31276 246204 31278
rect 281604 31276 282204 31278
rect 317604 31276 318204 31278
rect 353604 31276 354204 31278
rect 389604 31276 390204 31278
rect 425604 31276 426204 31278
rect 461604 31276 462204 31278
rect 497604 31276 498204 31278
rect 533604 31276 534204 31278
rect 569604 31276 570204 31278
rect 591760 31276 592360 31278
rect -8436 31254 592360 31276
rect -8436 31018 -8254 31254
rect -8018 31018 29786 31254
rect 30022 31018 65786 31254
rect 66022 31018 101786 31254
rect 102022 31018 137786 31254
rect 138022 31018 173786 31254
rect 174022 31018 209786 31254
rect 210022 31018 245786 31254
rect 246022 31018 281786 31254
rect 282022 31018 317786 31254
rect 318022 31018 353786 31254
rect 354022 31018 389786 31254
rect 390022 31018 425786 31254
rect 426022 31018 461786 31254
rect 462022 31018 497786 31254
rect 498022 31018 533786 31254
rect 534022 31018 569786 31254
rect 570022 31018 591942 31254
rect 592178 31018 592360 31254
rect -8436 30934 592360 31018
rect -8436 30698 -8254 30934
rect -8018 30698 29786 30934
rect 30022 30698 65786 30934
rect 66022 30698 101786 30934
rect 102022 30698 137786 30934
rect 138022 30698 173786 30934
rect 174022 30698 209786 30934
rect 210022 30698 245786 30934
rect 246022 30698 281786 30934
rect 282022 30698 317786 30934
rect 318022 30698 353786 30934
rect 354022 30698 389786 30934
rect 390022 30698 425786 30934
rect 426022 30698 461786 30934
rect 462022 30698 497786 30934
rect 498022 30698 533786 30934
rect 534022 30698 569786 30934
rect 570022 30698 591942 30934
rect 592178 30698 592360 30934
rect -8436 30676 592360 30698
rect -8436 30674 -7836 30676
rect 29604 30674 30204 30676
rect 65604 30674 66204 30676
rect 101604 30674 102204 30676
rect 137604 30674 138204 30676
rect 173604 30674 174204 30676
rect 209604 30674 210204 30676
rect 245604 30674 246204 30676
rect 281604 30674 282204 30676
rect 317604 30674 318204 30676
rect 353604 30674 354204 30676
rect 389604 30674 390204 30676
rect 425604 30674 426204 30676
rect 461604 30674 462204 30676
rect 497604 30674 498204 30676
rect 533604 30674 534204 30676
rect 569604 30674 570204 30676
rect 591760 30674 592360 30676
rect -6596 27676 -5996 27678
rect 26004 27676 26604 27678
rect 62004 27676 62604 27678
rect 98004 27676 98604 27678
rect 134004 27676 134604 27678
rect 170004 27676 170604 27678
rect 206004 27676 206604 27678
rect 242004 27676 242604 27678
rect 278004 27676 278604 27678
rect 314004 27676 314604 27678
rect 350004 27676 350604 27678
rect 386004 27676 386604 27678
rect 422004 27676 422604 27678
rect 458004 27676 458604 27678
rect 494004 27676 494604 27678
rect 530004 27676 530604 27678
rect 566004 27676 566604 27678
rect 589920 27676 590520 27678
rect -6596 27654 590520 27676
rect -6596 27418 -6414 27654
rect -6178 27418 26186 27654
rect 26422 27418 62186 27654
rect 62422 27418 98186 27654
rect 98422 27418 134186 27654
rect 134422 27418 170186 27654
rect 170422 27418 206186 27654
rect 206422 27418 242186 27654
rect 242422 27418 278186 27654
rect 278422 27418 314186 27654
rect 314422 27418 350186 27654
rect 350422 27418 386186 27654
rect 386422 27418 422186 27654
rect 422422 27418 458186 27654
rect 458422 27418 494186 27654
rect 494422 27418 530186 27654
rect 530422 27418 566186 27654
rect 566422 27418 590102 27654
rect 590338 27418 590520 27654
rect -6596 27334 590520 27418
rect -6596 27098 -6414 27334
rect -6178 27098 26186 27334
rect 26422 27098 62186 27334
rect 62422 27098 98186 27334
rect 98422 27098 134186 27334
rect 134422 27098 170186 27334
rect 170422 27098 206186 27334
rect 206422 27098 242186 27334
rect 242422 27098 278186 27334
rect 278422 27098 314186 27334
rect 314422 27098 350186 27334
rect 350422 27098 386186 27334
rect 386422 27098 422186 27334
rect 422422 27098 458186 27334
rect 458422 27098 494186 27334
rect 494422 27098 530186 27334
rect 530422 27098 566186 27334
rect 566422 27098 590102 27334
rect 590338 27098 590520 27334
rect -6596 27076 590520 27098
rect -6596 27074 -5996 27076
rect 26004 27074 26604 27076
rect 62004 27074 62604 27076
rect 98004 27074 98604 27076
rect 134004 27074 134604 27076
rect 170004 27074 170604 27076
rect 206004 27074 206604 27076
rect 242004 27074 242604 27076
rect 278004 27074 278604 27076
rect 314004 27074 314604 27076
rect 350004 27074 350604 27076
rect 386004 27074 386604 27076
rect 422004 27074 422604 27076
rect 458004 27074 458604 27076
rect 494004 27074 494604 27076
rect 530004 27074 530604 27076
rect 566004 27074 566604 27076
rect 589920 27074 590520 27076
rect -4756 24076 -4156 24078
rect 22404 24076 23004 24078
rect 58404 24076 59004 24078
rect 94404 24076 95004 24078
rect 130404 24076 131004 24078
rect 166404 24076 167004 24078
rect 202404 24076 203004 24078
rect 238404 24076 239004 24078
rect 274404 24076 275004 24078
rect 310404 24076 311004 24078
rect 346404 24076 347004 24078
rect 382404 24076 383004 24078
rect 418404 24076 419004 24078
rect 454404 24076 455004 24078
rect 490404 24076 491004 24078
rect 526404 24076 527004 24078
rect 562404 24076 563004 24078
rect 588080 24076 588680 24078
rect -4756 24054 588680 24076
rect -4756 23818 -4574 24054
rect -4338 23818 22586 24054
rect 22822 23818 58586 24054
rect 58822 23818 94586 24054
rect 94822 23818 130586 24054
rect 130822 23818 166586 24054
rect 166822 23818 202586 24054
rect 202822 23818 238586 24054
rect 238822 23818 274586 24054
rect 274822 23818 310586 24054
rect 310822 23818 346586 24054
rect 346822 23818 382586 24054
rect 382822 23818 418586 24054
rect 418822 23818 454586 24054
rect 454822 23818 490586 24054
rect 490822 23818 526586 24054
rect 526822 23818 562586 24054
rect 562822 23818 588262 24054
rect 588498 23818 588680 24054
rect -4756 23734 588680 23818
rect -4756 23498 -4574 23734
rect -4338 23498 22586 23734
rect 22822 23498 58586 23734
rect 58822 23498 94586 23734
rect 94822 23498 130586 23734
rect 130822 23498 166586 23734
rect 166822 23498 202586 23734
rect 202822 23498 238586 23734
rect 238822 23498 274586 23734
rect 274822 23498 310586 23734
rect 310822 23498 346586 23734
rect 346822 23498 382586 23734
rect 382822 23498 418586 23734
rect 418822 23498 454586 23734
rect 454822 23498 490586 23734
rect 490822 23498 526586 23734
rect 526822 23498 562586 23734
rect 562822 23498 588262 23734
rect 588498 23498 588680 23734
rect -4756 23476 588680 23498
rect -4756 23474 -4156 23476
rect 22404 23474 23004 23476
rect 58404 23474 59004 23476
rect 94404 23474 95004 23476
rect 130404 23474 131004 23476
rect 166404 23474 167004 23476
rect 202404 23474 203004 23476
rect 238404 23474 239004 23476
rect 274404 23474 275004 23476
rect 310404 23474 311004 23476
rect 346404 23474 347004 23476
rect 382404 23474 383004 23476
rect 418404 23474 419004 23476
rect 454404 23474 455004 23476
rect 490404 23474 491004 23476
rect 526404 23474 527004 23476
rect 562404 23474 563004 23476
rect 588080 23474 588680 23476
rect -2916 20476 -2316 20478
rect 18804 20476 19404 20478
rect 54804 20476 55404 20478
rect 90804 20476 91404 20478
rect 126804 20476 127404 20478
rect 162804 20476 163404 20478
rect 198804 20476 199404 20478
rect 234804 20476 235404 20478
rect 270804 20476 271404 20478
rect 306804 20476 307404 20478
rect 342804 20476 343404 20478
rect 378804 20476 379404 20478
rect 414804 20476 415404 20478
rect 450804 20476 451404 20478
rect 486804 20476 487404 20478
rect 522804 20476 523404 20478
rect 558804 20476 559404 20478
rect 586240 20476 586840 20478
rect -2916 20454 586840 20476
rect -2916 20218 -2734 20454
rect -2498 20218 18986 20454
rect 19222 20218 54986 20454
rect 55222 20218 90986 20454
rect 91222 20218 126986 20454
rect 127222 20218 162986 20454
rect 163222 20218 198986 20454
rect 199222 20218 234986 20454
rect 235222 20218 270986 20454
rect 271222 20218 306986 20454
rect 307222 20218 342986 20454
rect 343222 20218 378986 20454
rect 379222 20218 414986 20454
rect 415222 20218 450986 20454
rect 451222 20218 486986 20454
rect 487222 20218 522986 20454
rect 523222 20218 558986 20454
rect 559222 20218 586422 20454
rect 586658 20218 586840 20454
rect -2916 20134 586840 20218
rect -2916 19898 -2734 20134
rect -2498 19898 18986 20134
rect 19222 19898 54986 20134
rect 55222 19898 90986 20134
rect 91222 19898 126986 20134
rect 127222 19898 162986 20134
rect 163222 19898 198986 20134
rect 199222 19898 234986 20134
rect 235222 19898 270986 20134
rect 271222 19898 306986 20134
rect 307222 19898 342986 20134
rect 343222 19898 378986 20134
rect 379222 19898 414986 20134
rect 415222 19898 450986 20134
rect 451222 19898 486986 20134
rect 487222 19898 522986 20134
rect 523222 19898 558986 20134
rect 559222 19898 586422 20134
rect 586658 19898 586840 20134
rect -2916 19876 586840 19898
rect -2916 19874 -2316 19876
rect 18804 19874 19404 19876
rect 54804 19874 55404 19876
rect 90804 19874 91404 19876
rect 126804 19874 127404 19876
rect 162804 19874 163404 19876
rect 198804 19874 199404 19876
rect 234804 19874 235404 19876
rect 270804 19874 271404 19876
rect 306804 19874 307404 19876
rect 342804 19874 343404 19876
rect 378804 19874 379404 19876
rect 414804 19874 415404 19876
rect 450804 19874 451404 19876
rect 486804 19874 487404 19876
rect 522804 19874 523404 19876
rect 558804 19874 559404 19876
rect 586240 19874 586840 19876
rect -7516 13276 -6916 13278
rect 11604 13276 12204 13278
rect 47604 13276 48204 13278
rect 83604 13276 84204 13278
rect 119604 13276 120204 13278
rect 155604 13276 156204 13278
rect 191604 13276 192204 13278
rect 227604 13276 228204 13278
rect 263604 13276 264204 13278
rect 299604 13276 300204 13278
rect 335604 13276 336204 13278
rect 371604 13276 372204 13278
rect 407604 13276 408204 13278
rect 443604 13276 444204 13278
rect 479604 13276 480204 13278
rect 515604 13276 516204 13278
rect 551604 13276 552204 13278
rect 590840 13276 591440 13278
rect -8436 13254 592360 13276
rect -8436 13018 -7334 13254
rect -7098 13018 11786 13254
rect 12022 13018 47786 13254
rect 48022 13018 83786 13254
rect 84022 13018 119786 13254
rect 120022 13018 155786 13254
rect 156022 13018 191786 13254
rect 192022 13018 227786 13254
rect 228022 13018 263786 13254
rect 264022 13018 299786 13254
rect 300022 13018 335786 13254
rect 336022 13018 371786 13254
rect 372022 13018 407786 13254
rect 408022 13018 443786 13254
rect 444022 13018 479786 13254
rect 480022 13018 515786 13254
rect 516022 13018 551786 13254
rect 552022 13018 591022 13254
rect 591258 13018 592360 13254
rect -8436 12934 592360 13018
rect -8436 12698 -7334 12934
rect -7098 12698 11786 12934
rect 12022 12698 47786 12934
rect 48022 12698 83786 12934
rect 84022 12698 119786 12934
rect 120022 12698 155786 12934
rect 156022 12698 191786 12934
rect 192022 12698 227786 12934
rect 228022 12698 263786 12934
rect 264022 12698 299786 12934
rect 300022 12698 335786 12934
rect 336022 12698 371786 12934
rect 372022 12698 407786 12934
rect 408022 12698 443786 12934
rect 444022 12698 479786 12934
rect 480022 12698 515786 12934
rect 516022 12698 551786 12934
rect 552022 12698 591022 12934
rect 591258 12698 592360 12934
rect -8436 12676 592360 12698
rect -7516 12674 -6916 12676
rect 11604 12674 12204 12676
rect 47604 12674 48204 12676
rect 83604 12674 84204 12676
rect 119604 12674 120204 12676
rect 155604 12674 156204 12676
rect 191604 12674 192204 12676
rect 227604 12674 228204 12676
rect 263604 12674 264204 12676
rect 299604 12674 300204 12676
rect 335604 12674 336204 12676
rect 371604 12674 372204 12676
rect 407604 12674 408204 12676
rect 443604 12674 444204 12676
rect 479604 12674 480204 12676
rect 515604 12674 516204 12676
rect 551604 12674 552204 12676
rect 590840 12674 591440 12676
rect -5676 9676 -5076 9678
rect 8004 9676 8604 9678
rect 44004 9676 44604 9678
rect 80004 9676 80604 9678
rect 116004 9676 116604 9678
rect 152004 9676 152604 9678
rect 188004 9676 188604 9678
rect 224004 9676 224604 9678
rect 260004 9676 260604 9678
rect 296004 9676 296604 9678
rect 332004 9676 332604 9678
rect 368004 9676 368604 9678
rect 404004 9676 404604 9678
rect 440004 9676 440604 9678
rect 476004 9676 476604 9678
rect 512004 9676 512604 9678
rect 548004 9676 548604 9678
rect 589000 9676 589600 9678
rect -6596 9654 590520 9676
rect -6596 9418 -5494 9654
rect -5258 9418 8186 9654
rect 8422 9418 44186 9654
rect 44422 9418 80186 9654
rect 80422 9418 116186 9654
rect 116422 9418 152186 9654
rect 152422 9418 188186 9654
rect 188422 9418 224186 9654
rect 224422 9418 260186 9654
rect 260422 9418 296186 9654
rect 296422 9418 332186 9654
rect 332422 9418 368186 9654
rect 368422 9418 404186 9654
rect 404422 9418 440186 9654
rect 440422 9418 476186 9654
rect 476422 9418 512186 9654
rect 512422 9418 548186 9654
rect 548422 9418 589182 9654
rect 589418 9418 590520 9654
rect -6596 9334 590520 9418
rect -6596 9098 -5494 9334
rect -5258 9098 8186 9334
rect 8422 9098 44186 9334
rect 44422 9098 80186 9334
rect 80422 9098 116186 9334
rect 116422 9098 152186 9334
rect 152422 9098 188186 9334
rect 188422 9098 224186 9334
rect 224422 9098 260186 9334
rect 260422 9098 296186 9334
rect 296422 9098 332186 9334
rect 332422 9098 368186 9334
rect 368422 9098 404186 9334
rect 404422 9098 440186 9334
rect 440422 9098 476186 9334
rect 476422 9098 512186 9334
rect 512422 9098 548186 9334
rect 548422 9098 589182 9334
rect 589418 9098 590520 9334
rect -6596 9076 590520 9098
rect -5676 9074 -5076 9076
rect 8004 9074 8604 9076
rect 44004 9074 44604 9076
rect 80004 9074 80604 9076
rect 116004 9074 116604 9076
rect 152004 9074 152604 9076
rect 188004 9074 188604 9076
rect 224004 9074 224604 9076
rect 260004 9074 260604 9076
rect 296004 9074 296604 9076
rect 332004 9074 332604 9076
rect 368004 9074 368604 9076
rect 404004 9074 404604 9076
rect 440004 9074 440604 9076
rect 476004 9074 476604 9076
rect 512004 9074 512604 9076
rect 548004 9074 548604 9076
rect 589000 9074 589600 9076
rect -3836 6076 -3236 6078
rect 4404 6076 5004 6078
rect 40404 6076 41004 6078
rect 76404 6076 77004 6078
rect 112404 6076 113004 6078
rect 148404 6076 149004 6078
rect 184404 6076 185004 6078
rect 220404 6076 221004 6078
rect 256404 6076 257004 6078
rect 292404 6076 293004 6078
rect 328404 6076 329004 6078
rect 364404 6076 365004 6078
rect 400404 6076 401004 6078
rect 436404 6076 437004 6078
rect 472404 6076 473004 6078
rect 508404 6076 509004 6078
rect 544404 6076 545004 6078
rect 580404 6076 581004 6078
rect 587160 6076 587760 6078
rect -4756 6054 588680 6076
rect -4756 5818 -3654 6054
rect -3418 5818 4586 6054
rect 4822 5818 40586 6054
rect 40822 5818 76586 6054
rect 76822 5818 112586 6054
rect 112822 5818 148586 6054
rect 148822 5818 184586 6054
rect 184822 5818 220586 6054
rect 220822 5818 256586 6054
rect 256822 5818 292586 6054
rect 292822 5818 328586 6054
rect 328822 5818 364586 6054
rect 364822 5818 400586 6054
rect 400822 5818 436586 6054
rect 436822 5818 472586 6054
rect 472822 5818 508586 6054
rect 508822 5818 544586 6054
rect 544822 5818 580586 6054
rect 580822 5818 587342 6054
rect 587578 5818 588680 6054
rect -4756 5734 588680 5818
rect -4756 5498 -3654 5734
rect -3418 5498 4586 5734
rect 4822 5498 40586 5734
rect 40822 5498 76586 5734
rect 76822 5498 112586 5734
rect 112822 5498 148586 5734
rect 148822 5498 184586 5734
rect 184822 5498 220586 5734
rect 220822 5498 256586 5734
rect 256822 5498 292586 5734
rect 292822 5498 328586 5734
rect 328822 5498 364586 5734
rect 364822 5498 400586 5734
rect 400822 5498 436586 5734
rect 436822 5498 472586 5734
rect 472822 5498 508586 5734
rect 508822 5498 544586 5734
rect 544822 5498 580586 5734
rect 580822 5498 587342 5734
rect 587578 5498 588680 5734
rect -4756 5476 588680 5498
rect -3836 5474 -3236 5476
rect 4404 5474 5004 5476
rect 40404 5474 41004 5476
rect 76404 5474 77004 5476
rect 112404 5474 113004 5476
rect 148404 5474 149004 5476
rect 184404 5474 185004 5476
rect 220404 5474 221004 5476
rect 256404 5474 257004 5476
rect 292404 5474 293004 5476
rect 328404 5474 329004 5476
rect 364404 5474 365004 5476
rect 400404 5474 401004 5476
rect 436404 5474 437004 5476
rect 472404 5474 473004 5476
rect 508404 5474 509004 5476
rect 544404 5474 545004 5476
rect 580404 5474 581004 5476
rect 587160 5474 587760 5476
rect -1996 2476 -1396 2478
rect 804 2476 1404 2478
rect 36804 2476 37404 2478
rect 72804 2476 73404 2478
rect 108804 2476 109404 2478
rect 144804 2476 145404 2478
rect 180804 2476 181404 2478
rect 216804 2476 217404 2478
rect 252804 2476 253404 2478
rect 288804 2476 289404 2478
rect 324804 2476 325404 2478
rect 360804 2476 361404 2478
rect 396804 2476 397404 2478
rect 432804 2476 433404 2478
rect 468804 2476 469404 2478
rect 504804 2476 505404 2478
rect 540804 2476 541404 2478
rect 576804 2476 577404 2478
rect 585320 2476 585920 2478
rect -2916 2454 586840 2476
rect -2916 2218 -1814 2454
rect -1578 2218 986 2454
rect 1222 2218 36986 2454
rect 37222 2218 72986 2454
rect 73222 2218 108986 2454
rect 109222 2218 144986 2454
rect 145222 2218 180986 2454
rect 181222 2218 216986 2454
rect 217222 2218 252986 2454
rect 253222 2218 288986 2454
rect 289222 2218 324986 2454
rect 325222 2218 360986 2454
rect 361222 2218 396986 2454
rect 397222 2218 432986 2454
rect 433222 2218 468986 2454
rect 469222 2218 504986 2454
rect 505222 2218 540986 2454
rect 541222 2218 576986 2454
rect 577222 2218 585502 2454
rect 585738 2218 586840 2454
rect -2916 2134 586840 2218
rect -2916 1898 -1814 2134
rect -1578 1898 986 2134
rect 1222 1898 36986 2134
rect 37222 1898 72986 2134
rect 73222 1898 108986 2134
rect 109222 1898 144986 2134
rect 145222 1898 180986 2134
rect 181222 1898 216986 2134
rect 217222 1898 252986 2134
rect 253222 1898 288986 2134
rect 289222 1898 324986 2134
rect 325222 1898 360986 2134
rect 361222 1898 396986 2134
rect 397222 1898 432986 2134
rect 433222 1898 468986 2134
rect 469222 1898 504986 2134
rect 505222 1898 540986 2134
rect 541222 1898 576986 2134
rect 577222 1898 585502 2134
rect 585738 1898 586840 2134
rect -2916 1876 586840 1898
rect -1996 1874 -1396 1876
rect 804 1874 1404 1876
rect 36804 1874 37404 1876
rect 72804 1874 73404 1876
rect 108804 1874 109404 1876
rect 144804 1874 145404 1876
rect 180804 1874 181404 1876
rect 216804 1874 217404 1876
rect 252804 1874 253404 1876
rect 288804 1874 289404 1876
rect 324804 1874 325404 1876
rect 360804 1874 361404 1876
rect 396804 1874 397404 1876
rect 432804 1874 433404 1876
rect 468804 1874 469404 1876
rect 504804 1874 505404 1876
rect 540804 1874 541404 1876
rect 576804 1874 577404 1876
rect 585320 1874 585920 1876
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 144804 -324 145404 -322
rect 180804 -324 181404 -322
rect 216804 -324 217404 -322
rect 252804 -324 253404 -322
rect 288804 -324 289404 -322
rect 324804 -324 325404 -322
rect 360804 -324 361404 -322
rect 396804 -324 397404 -322
rect 432804 -324 433404 -322
rect 468804 -324 469404 -322
rect 504804 -324 505404 -322
rect 540804 -324 541404 -322
rect 576804 -324 577404 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 986 -346
rect 1222 -582 36986 -346
rect 37222 -582 72986 -346
rect 73222 -582 108986 -346
rect 109222 -582 144986 -346
rect 145222 -582 180986 -346
rect 181222 -582 216986 -346
rect 217222 -582 252986 -346
rect 253222 -582 288986 -346
rect 289222 -582 324986 -346
rect 325222 -582 360986 -346
rect 361222 -582 396986 -346
rect 397222 -582 432986 -346
rect 433222 -582 468986 -346
rect 469222 -582 504986 -346
rect 505222 -582 540986 -346
rect 541222 -582 576986 -346
rect 577222 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 986 -666
rect 1222 -902 36986 -666
rect 37222 -902 72986 -666
rect 73222 -902 108986 -666
rect 109222 -902 144986 -666
rect 145222 -902 180986 -666
rect 181222 -902 216986 -666
rect 217222 -902 252986 -666
rect 253222 -902 288986 -666
rect 289222 -902 324986 -666
rect 325222 -902 360986 -666
rect 361222 -902 396986 -666
rect 397222 -902 432986 -666
rect 433222 -902 468986 -666
rect 469222 -902 504986 -666
rect 505222 -902 540986 -666
rect 541222 -902 576986 -666
rect 577222 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 144804 -926 145404 -924
rect 180804 -926 181404 -924
rect 216804 -926 217404 -924
rect 252804 -926 253404 -924
rect 288804 -926 289404 -924
rect 324804 -926 325404 -924
rect 360804 -926 361404 -924
rect 396804 -926 397404 -924
rect 432804 -926 433404 -924
rect 468804 -926 469404 -924
rect 504804 -926 505404 -924
rect 540804 -926 541404 -924
rect 576804 -926 577404 -924
rect 585320 -926 585920 -924
rect -2916 -1244 -2316 -1242
rect 18804 -1244 19404 -1242
rect 54804 -1244 55404 -1242
rect 90804 -1244 91404 -1242
rect 126804 -1244 127404 -1242
rect 162804 -1244 163404 -1242
rect 198804 -1244 199404 -1242
rect 234804 -1244 235404 -1242
rect 270804 -1244 271404 -1242
rect 306804 -1244 307404 -1242
rect 342804 -1244 343404 -1242
rect 378804 -1244 379404 -1242
rect 414804 -1244 415404 -1242
rect 450804 -1244 451404 -1242
rect 486804 -1244 487404 -1242
rect 522804 -1244 523404 -1242
rect 558804 -1244 559404 -1242
rect 586240 -1244 586840 -1242
rect -2916 -1266 586840 -1244
rect -2916 -1502 -2734 -1266
rect -2498 -1502 18986 -1266
rect 19222 -1502 54986 -1266
rect 55222 -1502 90986 -1266
rect 91222 -1502 126986 -1266
rect 127222 -1502 162986 -1266
rect 163222 -1502 198986 -1266
rect 199222 -1502 234986 -1266
rect 235222 -1502 270986 -1266
rect 271222 -1502 306986 -1266
rect 307222 -1502 342986 -1266
rect 343222 -1502 378986 -1266
rect 379222 -1502 414986 -1266
rect 415222 -1502 450986 -1266
rect 451222 -1502 486986 -1266
rect 487222 -1502 522986 -1266
rect 523222 -1502 558986 -1266
rect 559222 -1502 586422 -1266
rect 586658 -1502 586840 -1266
rect -2916 -1586 586840 -1502
rect -2916 -1822 -2734 -1586
rect -2498 -1822 18986 -1586
rect 19222 -1822 54986 -1586
rect 55222 -1822 90986 -1586
rect 91222 -1822 126986 -1586
rect 127222 -1822 162986 -1586
rect 163222 -1822 198986 -1586
rect 199222 -1822 234986 -1586
rect 235222 -1822 270986 -1586
rect 271222 -1822 306986 -1586
rect 307222 -1822 342986 -1586
rect 343222 -1822 378986 -1586
rect 379222 -1822 414986 -1586
rect 415222 -1822 450986 -1586
rect 451222 -1822 486986 -1586
rect 487222 -1822 522986 -1586
rect 523222 -1822 558986 -1586
rect 559222 -1822 586422 -1586
rect 586658 -1822 586840 -1586
rect -2916 -1844 586840 -1822
rect -2916 -1846 -2316 -1844
rect 18804 -1846 19404 -1844
rect 54804 -1846 55404 -1844
rect 90804 -1846 91404 -1844
rect 126804 -1846 127404 -1844
rect 162804 -1846 163404 -1844
rect 198804 -1846 199404 -1844
rect 234804 -1846 235404 -1844
rect 270804 -1846 271404 -1844
rect 306804 -1846 307404 -1844
rect 342804 -1846 343404 -1844
rect 378804 -1846 379404 -1844
rect 414804 -1846 415404 -1844
rect 450804 -1846 451404 -1844
rect 486804 -1846 487404 -1844
rect 522804 -1846 523404 -1844
rect 558804 -1846 559404 -1844
rect 586240 -1846 586840 -1844
rect -3836 -2164 -3236 -2162
rect 4404 -2164 5004 -2162
rect 40404 -2164 41004 -2162
rect 76404 -2164 77004 -2162
rect 112404 -2164 113004 -2162
rect 148404 -2164 149004 -2162
rect 184404 -2164 185004 -2162
rect 220404 -2164 221004 -2162
rect 256404 -2164 257004 -2162
rect 292404 -2164 293004 -2162
rect 328404 -2164 329004 -2162
rect 364404 -2164 365004 -2162
rect 400404 -2164 401004 -2162
rect 436404 -2164 437004 -2162
rect 472404 -2164 473004 -2162
rect 508404 -2164 509004 -2162
rect 544404 -2164 545004 -2162
rect 580404 -2164 581004 -2162
rect 587160 -2164 587760 -2162
rect -3836 -2186 587760 -2164
rect -3836 -2422 -3654 -2186
rect -3418 -2422 4586 -2186
rect 4822 -2422 40586 -2186
rect 40822 -2422 76586 -2186
rect 76822 -2422 112586 -2186
rect 112822 -2422 148586 -2186
rect 148822 -2422 184586 -2186
rect 184822 -2422 220586 -2186
rect 220822 -2422 256586 -2186
rect 256822 -2422 292586 -2186
rect 292822 -2422 328586 -2186
rect 328822 -2422 364586 -2186
rect 364822 -2422 400586 -2186
rect 400822 -2422 436586 -2186
rect 436822 -2422 472586 -2186
rect 472822 -2422 508586 -2186
rect 508822 -2422 544586 -2186
rect 544822 -2422 580586 -2186
rect 580822 -2422 587342 -2186
rect 587578 -2422 587760 -2186
rect -3836 -2506 587760 -2422
rect -3836 -2742 -3654 -2506
rect -3418 -2742 4586 -2506
rect 4822 -2742 40586 -2506
rect 40822 -2742 76586 -2506
rect 76822 -2742 112586 -2506
rect 112822 -2742 148586 -2506
rect 148822 -2742 184586 -2506
rect 184822 -2742 220586 -2506
rect 220822 -2742 256586 -2506
rect 256822 -2742 292586 -2506
rect 292822 -2742 328586 -2506
rect 328822 -2742 364586 -2506
rect 364822 -2742 400586 -2506
rect 400822 -2742 436586 -2506
rect 436822 -2742 472586 -2506
rect 472822 -2742 508586 -2506
rect 508822 -2742 544586 -2506
rect 544822 -2742 580586 -2506
rect 580822 -2742 587342 -2506
rect 587578 -2742 587760 -2506
rect -3836 -2764 587760 -2742
rect -3836 -2766 -3236 -2764
rect 4404 -2766 5004 -2764
rect 40404 -2766 41004 -2764
rect 76404 -2766 77004 -2764
rect 112404 -2766 113004 -2764
rect 148404 -2766 149004 -2764
rect 184404 -2766 185004 -2764
rect 220404 -2766 221004 -2764
rect 256404 -2766 257004 -2764
rect 292404 -2766 293004 -2764
rect 328404 -2766 329004 -2764
rect 364404 -2766 365004 -2764
rect 400404 -2766 401004 -2764
rect 436404 -2766 437004 -2764
rect 472404 -2766 473004 -2764
rect 508404 -2766 509004 -2764
rect 544404 -2766 545004 -2764
rect 580404 -2766 581004 -2764
rect 587160 -2766 587760 -2764
rect -4756 -3084 -4156 -3082
rect 22404 -3084 23004 -3082
rect 58404 -3084 59004 -3082
rect 94404 -3084 95004 -3082
rect 130404 -3084 131004 -3082
rect 166404 -3084 167004 -3082
rect 202404 -3084 203004 -3082
rect 238404 -3084 239004 -3082
rect 274404 -3084 275004 -3082
rect 310404 -3084 311004 -3082
rect 346404 -3084 347004 -3082
rect 382404 -3084 383004 -3082
rect 418404 -3084 419004 -3082
rect 454404 -3084 455004 -3082
rect 490404 -3084 491004 -3082
rect 526404 -3084 527004 -3082
rect 562404 -3084 563004 -3082
rect 588080 -3084 588680 -3082
rect -4756 -3106 588680 -3084
rect -4756 -3342 -4574 -3106
rect -4338 -3342 22586 -3106
rect 22822 -3342 58586 -3106
rect 58822 -3342 94586 -3106
rect 94822 -3342 130586 -3106
rect 130822 -3342 166586 -3106
rect 166822 -3342 202586 -3106
rect 202822 -3342 238586 -3106
rect 238822 -3342 274586 -3106
rect 274822 -3342 310586 -3106
rect 310822 -3342 346586 -3106
rect 346822 -3342 382586 -3106
rect 382822 -3342 418586 -3106
rect 418822 -3342 454586 -3106
rect 454822 -3342 490586 -3106
rect 490822 -3342 526586 -3106
rect 526822 -3342 562586 -3106
rect 562822 -3342 588262 -3106
rect 588498 -3342 588680 -3106
rect -4756 -3426 588680 -3342
rect -4756 -3662 -4574 -3426
rect -4338 -3662 22586 -3426
rect 22822 -3662 58586 -3426
rect 58822 -3662 94586 -3426
rect 94822 -3662 130586 -3426
rect 130822 -3662 166586 -3426
rect 166822 -3662 202586 -3426
rect 202822 -3662 238586 -3426
rect 238822 -3662 274586 -3426
rect 274822 -3662 310586 -3426
rect 310822 -3662 346586 -3426
rect 346822 -3662 382586 -3426
rect 382822 -3662 418586 -3426
rect 418822 -3662 454586 -3426
rect 454822 -3662 490586 -3426
rect 490822 -3662 526586 -3426
rect 526822 -3662 562586 -3426
rect 562822 -3662 588262 -3426
rect 588498 -3662 588680 -3426
rect -4756 -3684 588680 -3662
rect -4756 -3686 -4156 -3684
rect 22404 -3686 23004 -3684
rect 58404 -3686 59004 -3684
rect 94404 -3686 95004 -3684
rect 130404 -3686 131004 -3684
rect 166404 -3686 167004 -3684
rect 202404 -3686 203004 -3684
rect 238404 -3686 239004 -3684
rect 274404 -3686 275004 -3684
rect 310404 -3686 311004 -3684
rect 346404 -3686 347004 -3684
rect 382404 -3686 383004 -3684
rect 418404 -3686 419004 -3684
rect 454404 -3686 455004 -3684
rect 490404 -3686 491004 -3684
rect 526404 -3686 527004 -3684
rect 562404 -3686 563004 -3684
rect 588080 -3686 588680 -3684
rect -5676 -4004 -5076 -4002
rect 8004 -4004 8604 -4002
rect 44004 -4004 44604 -4002
rect 80004 -4004 80604 -4002
rect 116004 -4004 116604 -4002
rect 152004 -4004 152604 -4002
rect 188004 -4004 188604 -4002
rect 224004 -4004 224604 -4002
rect 260004 -4004 260604 -4002
rect 296004 -4004 296604 -4002
rect 332004 -4004 332604 -4002
rect 368004 -4004 368604 -4002
rect 404004 -4004 404604 -4002
rect 440004 -4004 440604 -4002
rect 476004 -4004 476604 -4002
rect 512004 -4004 512604 -4002
rect 548004 -4004 548604 -4002
rect 589000 -4004 589600 -4002
rect -5676 -4026 589600 -4004
rect -5676 -4262 -5494 -4026
rect -5258 -4262 8186 -4026
rect 8422 -4262 44186 -4026
rect 44422 -4262 80186 -4026
rect 80422 -4262 116186 -4026
rect 116422 -4262 152186 -4026
rect 152422 -4262 188186 -4026
rect 188422 -4262 224186 -4026
rect 224422 -4262 260186 -4026
rect 260422 -4262 296186 -4026
rect 296422 -4262 332186 -4026
rect 332422 -4262 368186 -4026
rect 368422 -4262 404186 -4026
rect 404422 -4262 440186 -4026
rect 440422 -4262 476186 -4026
rect 476422 -4262 512186 -4026
rect 512422 -4262 548186 -4026
rect 548422 -4262 589182 -4026
rect 589418 -4262 589600 -4026
rect -5676 -4346 589600 -4262
rect -5676 -4582 -5494 -4346
rect -5258 -4582 8186 -4346
rect 8422 -4582 44186 -4346
rect 44422 -4582 80186 -4346
rect 80422 -4582 116186 -4346
rect 116422 -4582 152186 -4346
rect 152422 -4582 188186 -4346
rect 188422 -4582 224186 -4346
rect 224422 -4582 260186 -4346
rect 260422 -4582 296186 -4346
rect 296422 -4582 332186 -4346
rect 332422 -4582 368186 -4346
rect 368422 -4582 404186 -4346
rect 404422 -4582 440186 -4346
rect 440422 -4582 476186 -4346
rect 476422 -4582 512186 -4346
rect 512422 -4582 548186 -4346
rect 548422 -4582 589182 -4346
rect 589418 -4582 589600 -4346
rect -5676 -4604 589600 -4582
rect -5676 -4606 -5076 -4604
rect 8004 -4606 8604 -4604
rect 44004 -4606 44604 -4604
rect 80004 -4606 80604 -4604
rect 116004 -4606 116604 -4604
rect 152004 -4606 152604 -4604
rect 188004 -4606 188604 -4604
rect 224004 -4606 224604 -4604
rect 260004 -4606 260604 -4604
rect 296004 -4606 296604 -4604
rect 332004 -4606 332604 -4604
rect 368004 -4606 368604 -4604
rect 404004 -4606 404604 -4604
rect 440004 -4606 440604 -4604
rect 476004 -4606 476604 -4604
rect 512004 -4606 512604 -4604
rect 548004 -4606 548604 -4604
rect 589000 -4606 589600 -4604
rect -6596 -4924 -5996 -4922
rect 26004 -4924 26604 -4922
rect 62004 -4924 62604 -4922
rect 98004 -4924 98604 -4922
rect 134004 -4924 134604 -4922
rect 170004 -4924 170604 -4922
rect 206004 -4924 206604 -4922
rect 242004 -4924 242604 -4922
rect 278004 -4924 278604 -4922
rect 314004 -4924 314604 -4922
rect 350004 -4924 350604 -4922
rect 386004 -4924 386604 -4922
rect 422004 -4924 422604 -4922
rect 458004 -4924 458604 -4922
rect 494004 -4924 494604 -4922
rect 530004 -4924 530604 -4922
rect 566004 -4924 566604 -4922
rect 589920 -4924 590520 -4922
rect -6596 -4946 590520 -4924
rect -6596 -5182 -6414 -4946
rect -6178 -5182 26186 -4946
rect 26422 -5182 62186 -4946
rect 62422 -5182 98186 -4946
rect 98422 -5182 134186 -4946
rect 134422 -5182 170186 -4946
rect 170422 -5182 206186 -4946
rect 206422 -5182 242186 -4946
rect 242422 -5182 278186 -4946
rect 278422 -5182 314186 -4946
rect 314422 -5182 350186 -4946
rect 350422 -5182 386186 -4946
rect 386422 -5182 422186 -4946
rect 422422 -5182 458186 -4946
rect 458422 -5182 494186 -4946
rect 494422 -5182 530186 -4946
rect 530422 -5182 566186 -4946
rect 566422 -5182 590102 -4946
rect 590338 -5182 590520 -4946
rect -6596 -5266 590520 -5182
rect -6596 -5502 -6414 -5266
rect -6178 -5502 26186 -5266
rect 26422 -5502 62186 -5266
rect 62422 -5502 98186 -5266
rect 98422 -5502 134186 -5266
rect 134422 -5502 170186 -5266
rect 170422 -5502 206186 -5266
rect 206422 -5502 242186 -5266
rect 242422 -5502 278186 -5266
rect 278422 -5502 314186 -5266
rect 314422 -5502 350186 -5266
rect 350422 -5502 386186 -5266
rect 386422 -5502 422186 -5266
rect 422422 -5502 458186 -5266
rect 458422 -5502 494186 -5266
rect 494422 -5502 530186 -5266
rect 530422 -5502 566186 -5266
rect 566422 -5502 590102 -5266
rect 590338 -5502 590520 -5266
rect -6596 -5524 590520 -5502
rect -6596 -5526 -5996 -5524
rect 26004 -5526 26604 -5524
rect 62004 -5526 62604 -5524
rect 98004 -5526 98604 -5524
rect 134004 -5526 134604 -5524
rect 170004 -5526 170604 -5524
rect 206004 -5526 206604 -5524
rect 242004 -5526 242604 -5524
rect 278004 -5526 278604 -5524
rect 314004 -5526 314604 -5524
rect 350004 -5526 350604 -5524
rect 386004 -5526 386604 -5524
rect 422004 -5526 422604 -5524
rect 458004 -5526 458604 -5524
rect 494004 -5526 494604 -5524
rect 530004 -5526 530604 -5524
rect 566004 -5526 566604 -5524
rect 589920 -5526 590520 -5524
rect -7516 -5844 -6916 -5842
rect 11604 -5844 12204 -5842
rect 47604 -5844 48204 -5842
rect 83604 -5844 84204 -5842
rect 119604 -5844 120204 -5842
rect 155604 -5844 156204 -5842
rect 191604 -5844 192204 -5842
rect 227604 -5844 228204 -5842
rect 263604 -5844 264204 -5842
rect 299604 -5844 300204 -5842
rect 335604 -5844 336204 -5842
rect 371604 -5844 372204 -5842
rect 407604 -5844 408204 -5842
rect 443604 -5844 444204 -5842
rect 479604 -5844 480204 -5842
rect 515604 -5844 516204 -5842
rect 551604 -5844 552204 -5842
rect 590840 -5844 591440 -5842
rect -7516 -5866 591440 -5844
rect -7516 -6102 -7334 -5866
rect -7098 -6102 11786 -5866
rect 12022 -6102 47786 -5866
rect 48022 -6102 83786 -5866
rect 84022 -6102 119786 -5866
rect 120022 -6102 155786 -5866
rect 156022 -6102 191786 -5866
rect 192022 -6102 227786 -5866
rect 228022 -6102 263786 -5866
rect 264022 -6102 299786 -5866
rect 300022 -6102 335786 -5866
rect 336022 -6102 371786 -5866
rect 372022 -6102 407786 -5866
rect 408022 -6102 443786 -5866
rect 444022 -6102 479786 -5866
rect 480022 -6102 515786 -5866
rect 516022 -6102 551786 -5866
rect 552022 -6102 591022 -5866
rect 591258 -6102 591440 -5866
rect -7516 -6186 591440 -6102
rect -7516 -6422 -7334 -6186
rect -7098 -6422 11786 -6186
rect 12022 -6422 47786 -6186
rect 48022 -6422 83786 -6186
rect 84022 -6422 119786 -6186
rect 120022 -6422 155786 -6186
rect 156022 -6422 191786 -6186
rect 192022 -6422 227786 -6186
rect 228022 -6422 263786 -6186
rect 264022 -6422 299786 -6186
rect 300022 -6422 335786 -6186
rect 336022 -6422 371786 -6186
rect 372022 -6422 407786 -6186
rect 408022 -6422 443786 -6186
rect 444022 -6422 479786 -6186
rect 480022 -6422 515786 -6186
rect 516022 -6422 551786 -6186
rect 552022 -6422 591022 -6186
rect 591258 -6422 591440 -6186
rect -7516 -6444 591440 -6422
rect -7516 -6446 -6916 -6444
rect 11604 -6446 12204 -6444
rect 47604 -6446 48204 -6444
rect 83604 -6446 84204 -6444
rect 119604 -6446 120204 -6444
rect 155604 -6446 156204 -6444
rect 191604 -6446 192204 -6444
rect 227604 -6446 228204 -6444
rect 263604 -6446 264204 -6444
rect 299604 -6446 300204 -6444
rect 335604 -6446 336204 -6444
rect 371604 -6446 372204 -6444
rect 407604 -6446 408204 -6444
rect 443604 -6446 444204 -6444
rect 479604 -6446 480204 -6444
rect 515604 -6446 516204 -6444
rect 551604 -6446 552204 -6444
rect 590840 -6446 591440 -6444
rect -8436 -6764 -7836 -6762
rect 29604 -6764 30204 -6762
rect 65604 -6764 66204 -6762
rect 101604 -6764 102204 -6762
rect 137604 -6764 138204 -6762
rect 173604 -6764 174204 -6762
rect 209604 -6764 210204 -6762
rect 245604 -6764 246204 -6762
rect 281604 -6764 282204 -6762
rect 317604 -6764 318204 -6762
rect 353604 -6764 354204 -6762
rect 389604 -6764 390204 -6762
rect 425604 -6764 426204 -6762
rect 461604 -6764 462204 -6762
rect 497604 -6764 498204 -6762
rect 533604 -6764 534204 -6762
rect 569604 -6764 570204 -6762
rect 591760 -6764 592360 -6762
rect -8436 -6786 592360 -6764
rect -8436 -7022 -8254 -6786
rect -8018 -7022 29786 -6786
rect 30022 -7022 65786 -6786
rect 66022 -7022 101786 -6786
rect 102022 -7022 137786 -6786
rect 138022 -7022 173786 -6786
rect 174022 -7022 209786 -6786
rect 210022 -7022 245786 -6786
rect 246022 -7022 281786 -6786
rect 282022 -7022 317786 -6786
rect 318022 -7022 353786 -6786
rect 354022 -7022 389786 -6786
rect 390022 -7022 425786 -6786
rect 426022 -7022 461786 -6786
rect 462022 -7022 497786 -6786
rect 498022 -7022 533786 -6786
rect 534022 -7022 569786 -6786
rect 570022 -7022 591942 -6786
rect 592178 -7022 592360 -6786
rect -8436 -7106 592360 -7022
rect -8436 -7342 -8254 -7106
rect -8018 -7342 29786 -7106
rect 30022 -7342 65786 -7106
rect 66022 -7342 101786 -7106
rect 102022 -7342 137786 -7106
rect 138022 -7342 173786 -7106
rect 174022 -7342 209786 -7106
rect 210022 -7342 245786 -7106
rect 246022 -7342 281786 -7106
rect 282022 -7342 317786 -7106
rect 318022 -7342 353786 -7106
rect 354022 -7342 389786 -7106
rect 390022 -7342 425786 -7106
rect 426022 -7342 461786 -7106
rect 462022 -7342 497786 -7106
rect 498022 -7342 533786 -7106
rect 534022 -7342 569786 -7106
rect 570022 -7342 591942 -7106
rect 592178 -7342 592360 -7106
rect -8436 -7364 592360 -7342
rect -8436 -7366 -7836 -7364
rect 29604 -7366 30204 -7364
rect 65604 -7366 66204 -7364
rect 101604 -7366 102204 -7364
rect 137604 -7366 138204 -7364
rect 173604 -7366 174204 -7364
rect 209604 -7366 210204 -7364
rect 245604 -7366 246204 -7364
rect 281604 -7366 282204 -7364
rect 317604 -7366 318204 -7364
rect 353604 -7366 354204 -7364
rect 389604 -7366 390204 -7364
rect 425604 -7366 426204 -7364
rect 461604 -7366 462204 -7364
rect 497604 -7366 498204 -7364
rect 533604 -7366 534204 -7364
rect 569604 -7366 570204 -7364
rect 591760 -7366 592360 -7364
use user_proj_example  mprj
timestamp 1607892876
transform 1 0 229999 0 1 340000
box 1 0 219578 220000
<< labels >>
rlabel metal3 s 583520 5796 584960 6036 6 analog_io[0]
port 0 nsew default bidirectional
rlabel metal3 s 583520 474996 584960 475236 6 analog_io[10]
port 1 nsew default bidirectional
rlabel metal3 s 583520 521916 584960 522156 6 analog_io[11]
port 2 nsew default bidirectional
rlabel metal3 s 583520 568836 584960 569076 6 analog_io[12]
port 3 nsew default bidirectional
rlabel metal3 s 583520 615756 584960 615996 6 analog_io[13]
port 4 nsew default bidirectional
rlabel metal3 s 583520 662676 584960 662916 6 analog_io[14]
port 5 nsew default bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[15]
port 6 nsew default bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[16]
port 7 nsew default bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[17]
port 8 nsew default bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[18]
port 9 nsew default bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[19]
port 10 nsew default bidirectional
rlabel metal3 s 583520 52716 584960 52956 6 analog_io[1]
port 11 nsew default bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[20]
port 12 nsew default bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[21]
port 13 nsew default bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[22]
port 14 nsew default bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[23]
port 15 nsew default bidirectional
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 16 nsew default bidirectional
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 17 nsew default bidirectional
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 18 nsew default bidirectional
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 19 nsew default bidirectional
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 20 nsew default bidirectional
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 21 nsew default bidirectional
rlabel metal3 s 583520 99636 584960 99876 6 analog_io[2]
port 22 nsew default bidirectional
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 23 nsew default bidirectional
rlabel metal3 s 583520 146556 584960 146796 6 analog_io[3]
port 24 nsew default bidirectional
rlabel metal3 s 583520 193476 584960 193716 6 analog_io[4]
port 25 nsew default bidirectional
rlabel metal3 s 583520 240396 584960 240636 6 analog_io[5]
port 26 nsew default bidirectional
rlabel metal3 s 583520 287316 584960 287556 6 analog_io[6]
port 27 nsew default bidirectional
rlabel metal3 s 583520 334236 584960 334476 6 analog_io[7]
port 28 nsew default bidirectional
rlabel metal3 s 583520 381156 584960 381396 6 analog_io[8]
port 29 nsew default bidirectional
rlabel metal3 s 583520 428076 584960 428316 6 analog_io[9]
port 30 nsew default bidirectional
rlabel metal3 s 583520 17492 584960 17732 6 io_in[0]
port 31 nsew default input
rlabel metal3 s 583520 486692 584960 486932 6 io_in[10]
port 32 nsew default input
rlabel metal3 s 583520 533748 584960 533988 6 io_in[11]
port 33 nsew default input
rlabel metal3 s 583520 580668 584960 580908 6 io_in[12]
port 34 nsew default input
rlabel metal3 s 583520 627588 584960 627828 6 io_in[13]
port 35 nsew default input
rlabel metal3 s 583520 674508 584960 674748 6 io_in[14]
port 36 nsew default input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 37 nsew default input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 38 nsew default input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 39 nsew default input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 40 nsew default input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 41 nsew default input
rlabel metal3 s 583520 64412 584960 64652 6 io_in[1]
port 42 nsew default input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 43 nsew default input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 44 nsew default input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 45 nsew default input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 46 nsew default input
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 47 nsew default input
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 48 nsew default input
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 49 nsew default input
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 50 nsew default input
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 51 nsew default input
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 52 nsew default input
rlabel metal3 s 583520 111332 584960 111572 6 io_in[2]
port 53 nsew default input
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 54 nsew default input
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 55 nsew default input
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 56 nsew default input
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 57 nsew default input
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 58 nsew default input
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 59 nsew default input
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 60 nsew default input
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 61 nsew default input
rlabel metal3 s 583520 158252 584960 158492 6 io_in[3]
port 62 nsew default input
rlabel metal3 s 583520 205172 584960 205412 6 io_in[4]
port 63 nsew default input
rlabel metal3 s 583520 252092 584960 252332 6 io_in[5]
port 64 nsew default input
rlabel metal3 s 583520 299012 584960 299252 6 io_in[6]
port 65 nsew default input
rlabel metal3 s 583520 345932 584960 346172 6 io_in[7]
port 66 nsew default input
rlabel metal3 s 583520 392852 584960 393092 6 io_in[8]
port 67 nsew default input
rlabel metal3 s 583520 439772 584960 440012 6 io_in[9]
port 68 nsew default input
rlabel metal3 s 583520 40884 584960 41124 6 io_oeb[0]
port 69 nsew default tristate
rlabel metal3 s 583520 510220 584960 510460 6 io_oeb[10]
port 70 nsew default tristate
rlabel metal3 s 583520 557140 584960 557380 6 io_oeb[11]
port 71 nsew default tristate
rlabel metal3 s 583520 604060 584960 604300 6 io_oeb[12]
port 72 nsew default tristate
rlabel metal3 s 583520 650980 584960 651220 6 io_oeb[13]
port 73 nsew default tristate
rlabel metal3 s 583520 697900 584960 698140 6 io_oeb[14]
port 74 nsew default tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 75 nsew default tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 76 nsew default tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 77 nsew default tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 78 nsew default tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 79 nsew default tristate
rlabel metal3 s 583520 87804 584960 88044 6 io_oeb[1]
port 80 nsew default tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 81 nsew default tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 82 nsew default tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 83 nsew default tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 84 nsew default tristate
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 85 nsew default tristate
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 86 nsew default tristate
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 87 nsew default tristate
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 88 nsew default tristate
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 89 nsew default tristate
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 90 nsew default tristate
rlabel metal3 s 583520 134724 584960 134964 6 io_oeb[2]
port 91 nsew default tristate
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 92 nsew default tristate
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 93 nsew default tristate
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 94 nsew default tristate
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 95 nsew default tristate
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 96 nsew default tristate
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 97 nsew default tristate
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 98 nsew default tristate
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 99 nsew default tristate
rlabel metal3 s 583520 181780 584960 182020 6 io_oeb[3]
port 100 nsew default tristate
rlabel metal3 s 583520 228700 584960 228940 6 io_oeb[4]
port 101 nsew default tristate
rlabel metal3 s 583520 275620 584960 275860 6 io_oeb[5]
port 102 nsew default tristate
rlabel metal3 s 583520 322540 584960 322780 6 io_oeb[6]
port 103 nsew default tristate
rlabel metal3 s 583520 369460 584960 369700 6 io_oeb[7]
port 104 nsew default tristate
rlabel metal3 s 583520 416380 584960 416620 6 io_oeb[8]
port 105 nsew default tristate
rlabel metal3 s 583520 463300 584960 463540 6 io_oeb[9]
port 106 nsew default tristate
rlabel metal3 s 583520 29188 584960 29428 6 io_out[0]
port 107 nsew default tristate
rlabel metal3 s 583520 498524 584960 498764 6 io_out[10]
port 108 nsew default tristate
rlabel metal3 s 583520 545444 584960 545684 6 io_out[11]
port 109 nsew default tristate
rlabel metal3 s 583520 592364 584960 592604 6 io_out[12]
port 110 nsew default tristate
rlabel metal3 s 583520 639284 584960 639524 6 io_out[13]
port 111 nsew default tristate
rlabel metal3 s 583520 686204 584960 686444 6 io_out[14]
port 112 nsew default tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 113 nsew default tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 114 nsew default tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 115 nsew default tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 116 nsew default tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 117 nsew default tristate
rlabel metal3 s 583520 76108 584960 76348 6 io_out[1]
port 118 nsew default tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 119 nsew default tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 120 nsew default tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 121 nsew default tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 122 nsew default tristate
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 123 nsew default tristate
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 124 nsew default tristate
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 125 nsew default tristate
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 126 nsew default tristate
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 127 nsew default tristate
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 128 nsew default tristate
rlabel metal3 s 583520 123028 584960 123268 6 io_out[2]
port 129 nsew default tristate
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 130 nsew default tristate
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 131 nsew default tristate
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 132 nsew default tristate
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 133 nsew default tristate
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 134 nsew default tristate
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 135 nsew default tristate
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 136 nsew default tristate
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 137 nsew default tristate
rlabel metal3 s 583520 169948 584960 170188 6 io_out[3]
port 138 nsew default tristate
rlabel metal3 s 583520 216868 584960 217108 6 io_out[4]
port 139 nsew default tristate
rlabel metal3 s 583520 263788 584960 264028 6 io_out[5]
port 140 nsew default tristate
rlabel metal3 s 583520 310708 584960 310948 6 io_out[6]
port 141 nsew default tristate
rlabel metal3 s 583520 357764 584960 358004 6 io_out[7]
port 142 nsew default tristate
rlabel metal3 s 583520 404684 584960 404924 6 io_out[8]
port 143 nsew default tristate
rlabel metal3 s 583520 451604 584960 451844 6 io_out[9]
port 144 nsew default tristate
rlabel metal2 s 126582 -960 126694 480 8 la_data_in[0]
port 145 nsew default input
rlabel metal2 s 483450 -960 483562 480 8 la_data_in[100]
port 146 nsew default input
rlabel metal2 s 486946 -960 487058 480 8 la_data_in[101]
port 147 nsew default input
rlabel metal2 s 490534 -960 490646 480 8 la_data_in[102]
port 148 nsew default input
rlabel metal2 s 494122 -960 494234 480 8 la_data_in[103]
port 149 nsew default input
rlabel metal2 s 497710 -960 497822 480 8 la_data_in[104]
port 150 nsew default input
rlabel metal2 s 501206 -960 501318 480 8 la_data_in[105]
port 151 nsew default input
rlabel metal2 s 504794 -960 504906 480 8 la_data_in[106]
port 152 nsew default input
rlabel metal2 s 508382 -960 508494 480 8 la_data_in[107]
port 153 nsew default input
rlabel metal2 s 511970 -960 512082 480 8 la_data_in[108]
port 154 nsew default input
rlabel metal2 s 515558 -960 515670 480 8 la_data_in[109]
port 155 nsew default input
rlabel metal2 s 162278 -960 162390 480 8 la_data_in[10]
port 156 nsew default input
rlabel metal2 s 519054 -960 519166 480 8 la_data_in[110]
port 157 nsew default input
rlabel metal2 s 522642 -960 522754 480 8 la_data_in[111]
port 158 nsew default input
rlabel metal2 s 526230 -960 526342 480 8 la_data_in[112]
port 159 nsew default input
rlabel metal2 s 529818 -960 529930 480 8 la_data_in[113]
port 160 nsew default input
rlabel metal2 s 533406 -960 533518 480 8 la_data_in[114]
port 161 nsew default input
rlabel metal2 s 536902 -960 537014 480 8 la_data_in[115]
port 162 nsew default input
rlabel metal2 s 540490 -960 540602 480 8 la_data_in[116]
port 163 nsew default input
rlabel metal2 s 544078 -960 544190 480 8 la_data_in[117]
port 164 nsew default input
rlabel metal2 s 547666 -960 547778 480 8 la_data_in[118]
port 165 nsew default input
rlabel metal2 s 551162 -960 551274 480 8 la_data_in[119]
port 166 nsew default input
rlabel metal2 s 165866 -960 165978 480 8 la_data_in[11]
port 167 nsew default input
rlabel metal2 s 554750 -960 554862 480 8 la_data_in[120]
port 168 nsew default input
rlabel metal2 s 558338 -960 558450 480 8 la_data_in[121]
port 169 nsew default input
rlabel metal2 s 561926 -960 562038 480 8 la_data_in[122]
port 170 nsew default input
rlabel metal2 s 565514 -960 565626 480 8 la_data_in[123]
port 171 nsew default input
rlabel metal2 s 569010 -960 569122 480 8 la_data_in[124]
port 172 nsew default input
rlabel metal2 s 572598 -960 572710 480 8 la_data_in[125]
port 173 nsew default input
rlabel metal2 s 576186 -960 576298 480 8 la_data_in[126]
port 174 nsew default input
rlabel metal2 s 579774 -960 579886 480 8 la_data_in[127]
port 175 nsew default input
rlabel metal2 s 169362 -960 169474 480 8 la_data_in[12]
port 176 nsew default input
rlabel metal2 s 172950 -960 173062 480 8 la_data_in[13]
port 177 nsew default input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[14]
port 178 nsew default input
rlabel metal2 s 180126 -960 180238 480 8 la_data_in[15]
port 179 nsew default input
rlabel metal2 s 183714 -960 183826 480 8 la_data_in[16]
port 180 nsew default input
rlabel metal2 s 187210 -960 187322 480 8 la_data_in[17]
port 181 nsew default input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[18]
port 182 nsew default input
rlabel metal2 s 194386 -960 194498 480 8 la_data_in[19]
port 183 nsew default input
rlabel metal2 s 130170 -960 130282 480 8 la_data_in[1]
port 184 nsew default input
rlabel metal2 s 197974 -960 198086 480 8 la_data_in[20]
port 185 nsew default input
rlabel metal2 s 201470 -960 201582 480 8 la_data_in[21]
port 186 nsew default input
rlabel metal2 s 205058 -960 205170 480 8 la_data_in[22]
port 187 nsew default input
rlabel metal2 s 208646 -960 208758 480 8 la_data_in[23]
port 188 nsew default input
rlabel metal2 s 212234 -960 212346 480 8 la_data_in[24]
port 189 nsew default input
rlabel metal2 s 215822 -960 215934 480 8 la_data_in[25]
port 190 nsew default input
rlabel metal2 s 219318 -960 219430 480 8 la_data_in[26]
port 191 nsew default input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[27]
port 192 nsew default input
rlabel metal2 s 226494 -960 226606 480 8 la_data_in[28]
port 193 nsew default input
rlabel metal2 s 230082 -960 230194 480 8 la_data_in[29]
port 194 nsew default input
rlabel metal2 s 133758 -960 133870 480 8 la_data_in[2]
port 195 nsew default input
rlabel metal2 s 233670 -960 233782 480 8 la_data_in[30]
port 196 nsew default input
rlabel metal2 s 237166 -960 237278 480 8 la_data_in[31]
port 197 nsew default input
rlabel metal2 s 240754 -960 240866 480 8 la_data_in[32]
port 198 nsew default input
rlabel metal2 s 244342 -960 244454 480 8 la_data_in[33]
port 199 nsew default input
rlabel metal2 s 247930 -960 248042 480 8 la_data_in[34]
port 200 nsew default input
rlabel metal2 s 251426 -960 251538 480 8 la_data_in[35]
port 201 nsew default input
rlabel metal2 s 255014 -960 255126 480 8 la_data_in[36]
port 202 nsew default input
rlabel metal2 s 258602 -960 258714 480 8 la_data_in[37]
port 203 nsew default input
rlabel metal2 s 262190 -960 262302 480 8 la_data_in[38]
port 204 nsew default input
rlabel metal2 s 265778 -960 265890 480 8 la_data_in[39]
port 205 nsew default input
rlabel metal2 s 137254 -960 137366 480 8 la_data_in[3]
port 206 nsew default input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 207 nsew default input
rlabel metal2 s 272862 -960 272974 480 8 la_data_in[41]
port 208 nsew default input
rlabel metal2 s 276450 -960 276562 480 8 la_data_in[42]
port 209 nsew default input
rlabel metal2 s 280038 -960 280150 480 8 la_data_in[43]
port 210 nsew default input
rlabel metal2 s 283626 -960 283738 480 8 la_data_in[44]
port 211 nsew default input
rlabel metal2 s 287122 -960 287234 480 8 la_data_in[45]
port 212 nsew default input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[46]
port 213 nsew default input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[47]
port 214 nsew default input
rlabel metal2 s 297886 -960 297998 480 8 la_data_in[48]
port 215 nsew default input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[49]
port 216 nsew default input
rlabel metal2 s 140842 -960 140954 480 8 la_data_in[4]
port 217 nsew default input
rlabel metal2 s 304970 -960 305082 480 8 la_data_in[50]
port 218 nsew default input
rlabel metal2 s 308558 -960 308670 480 8 la_data_in[51]
port 219 nsew default input
rlabel metal2 s 312146 -960 312258 480 8 la_data_in[52]
port 220 nsew default input
rlabel metal2 s 315734 -960 315846 480 8 la_data_in[53]
port 221 nsew default input
rlabel metal2 s 319230 -960 319342 480 8 la_data_in[54]
port 222 nsew default input
rlabel metal2 s 322818 -960 322930 480 8 la_data_in[55]
port 223 nsew default input
rlabel metal2 s 326406 -960 326518 480 8 la_data_in[56]
port 224 nsew default input
rlabel metal2 s 329994 -960 330106 480 8 la_data_in[57]
port 225 nsew default input
rlabel metal2 s 333582 -960 333694 480 8 la_data_in[58]
port 226 nsew default input
rlabel metal2 s 337078 -960 337190 480 8 la_data_in[59]
port 227 nsew default input
rlabel metal2 s 144430 -960 144542 480 8 la_data_in[5]
port 228 nsew default input
rlabel metal2 s 340666 -960 340778 480 8 la_data_in[60]
port 229 nsew default input
rlabel metal2 s 344254 -960 344366 480 8 la_data_in[61]
port 230 nsew default input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[62]
port 231 nsew default input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[63]
port 232 nsew default input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[64]
port 233 nsew default input
rlabel metal2 s 358514 -960 358626 480 8 la_data_in[65]
port 234 nsew default input
rlabel metal2 s 362102 -960 362214 480 8 la_data_in[66]
port 235 nsew default input
rlabel metal2 s 365690 -960 365802 480 8 la_data_in[67]
port 236 nsew default input
rlabel metal2 s 369186 -960 369298 480 8 la_data_in[68]
port 237 nsew default input
rlabel metal2 s 372774 -960 372886 480 8 la_data_in[69]
port 238 nsew default input
rlabel metal2 s 148018 -960 148130 480 8 la_data_in[6]
port 239 nsew default input
rlabel metal2 s 376362 -960 376474 480 8 la_data_in[70]
port 240 nsew default input
rlabel metal2 s 379950 -960 380062 480 8 la_data_in[71]
port 241 nsew default input
rlabel metal2 s 383538 -960 383650 480 8 la_data_in[72]
port 242 nsew default input
rlabel metal2 s 387034 -960 387146 480 8 la_data_in[73]
port 243 nsew default input
rlabel metal2 s 390622 -960 390734 480 8 la_data_in[74]
port 244 nsew default input
rlabel metal2 s 394210 -960 394322 480 8 la_data_in[75]
port 245 nsew default input
rlabel metal2 s 397798 -960 397910 480 8 la_data_in[76]
port 246 nsew default input
rlabel metal2 s 401294 -960 401406 480 8 la_data_in[77]
port 247 nsew default input
rlabel metal2 s 404882 -960 404994 480 8 la_data_in[78]
port 248 nsew default input
rlabel metal2 s 408470 -960 408582 480 8 la_data_in[79]
port 249 nsew default input
rlabel metal2 s 151514 -960 151626 480 8 la_data_in[7]
port 250 nsew default input
rlabel metal2 s 412058 -960 412170 480 8 la_data_in[80]
port 251 nsew default input
rlabel metal2 s 415646 -960 415758 480 8 la_data_in[81]
port 252 nsew default input
rlabel metal2 s 419142 -960 419254 480 8 la_data_in[82]
port 253 nsew default input
rlabel metal2 s 422730 -960 422842 480 8 la_data_in[83]
port 254 nsew default input
rlabel metal2 s 426318 -960 426430 480 8 la_data_in[84]
port 255 nsew default input
rlabel metal2 s 429906 -960 430018 480 8 la_data_in[85]
port 256 nsew default input
rlabel metal2 s 433494 -960 433606 480 8 la_data_in[86]
port 257 nsew default input
rlabel metal2 s 436990 -960 437102 480 8 la_data_in[87]
port 258 nsew default input
rlabel metal2 s 440578 -960 440690 480 8 la_data_in[88]
port 259 nsew default input
rlabel metal2 s 444166 -960 444278 480 8 la_data_in[89]
port 260 nsew default input
rlabel metal2 s 155102 -960 155214 480 8 la_data_in[8]
port 261 nsew default input
rlabel metal2 s 447754 -960 447866 480 8 la_data_in[90]
port 262 nsew default input
rlabel metal2 s 451250 -960 451362 480 8 la_data_in[91]
port 263 nsew default input
rlabel metal2 s 454838 -960 454950 480 8 la_data_in[92]
port 264 nsew default input
rlabel metal2 s 458426 -960 458538 480 8 la_data_in[93]
port 265 nsew default input
rlabel metal2 s 462014 -960 462126 480 8 la_data_in[94]
port 266 nsew default input
rlabel metal2 s 465602 -960 465714 480 8 la_data_in[95]
port 267 nsew default input
rlabel metal2 s 469098 -960 469210 480 8 la_data_in[96]
port 268 nsew default input
rlabel metal2 s 472686 -960 472798 480 8 la_data_in[97]
port 269 nsew default input
rlabel metal2 s 476274 -960 476386 480 8 la_data_in[98]
port 270 nsew default input
rlabel metal2 s 479862 -960 479974 480 8 la_data_in[99]
port 271 nsew default input
rlabel metal2 s 158690 -960 158802 480 8 la_data_in[9]
port 272 nsew default input
rlabel metal2 s 127778 -960 127890 480 8 la_data_out[0]
port 273 nsew default tristate
rlabel metal2 s 484554 -960 484666 480 8 la_data_out[100]
port 274 nsew default tristate
rlabel metal2 s 488142 -960 488254 480 8 la_data_out[101]
port 275 nsew default tristate
rlabel metal2 s 491730 -960 491842 480 8 la_data_out[102]
port 276 nsew default tristate
rlabel metal2 s 495318 -960 495430 480 8 la_data_out[103]
port 277 nsew default tristate
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[104]
port 278 nsew default tristate
rlabel metal2 s 502402 -960 502514 480 8 la_data_out[105]
port 279 nsew default tristate
rlabel metal2 s 505990 -960 506102 480 8 la_data_out[106]
port 280 nsew default tristate
rlabel metal2 s 509578 -960 509690 480 8 la_data_out[107]
port 281 nsew default tristate
rlabel metal2 s 513166 -960 513278 480 8 la_data_out[108]
port 282 nsew default tristate
rlabel metal2 s 516754 -960 516866 480 8 la_data_out[109]
port 283 nsew default tristate
rlabel metal2 s 163474 -960 163586 480 8 la_data_out[10]
port 284 nsew default tristate
rlabel metal2 s 520250 -960 520362 480 8 la_data_out[110]
port 285 nsew default tristate
rlabel metal2 s 523838 -960 523950 480 8 la_data_out[111]
port 286 nsew default tristate
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[112]
port 287 nsew default tristate
rlabel metal2 s 531014 -960 531126 480 8 la_data_out[113]
port 288 nsew default tristate
rlabel metal2 s 534510 -960 534622 480 8 la_data_out[114]
port 289 nsew default tristate
rlabel metal2 s 538098 -960 538210 480 8 la_data_out[115]
port 290 nsew default tristate
rlabel metal2 s 541686 -960 541798 480 8 la_data_out[116]
port 291 nsew default tristate
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[117]
port 292 nsew default tristate
rlabel metal2 s 548862 -960 548974 480 8 la_data_out[118]
port 293 nsew default tristate
rlabel metal2 s 552358 -960 552470 480 8 la_data_out[119]
port 294 nsew default tristate
rlabel metal2 s 167062 -960 167174 480 8 la_data_out[11]
port 295 nsew default tristate
rlabel metal2 s 555946 -960 556058 480 8 la_data_out[120]
port 296 nsew default tristate
rlabel metal2 s 559534 -960 559646 480 8 la_data_out[121]
port 297 nsew default tristate
rlabel metal2 s 563122 -960 563234 480 8 la_data_out[122]
port 298 nsew default tristate
rlabel metal2 s 566710 -960 566822 480 8 la_data_out[123]
port 299 nsew default tristate
rlabel metal2 s 570206 -960 570318 480 8 la_data_out[124]
port 300 nsew default tristate
rlabel metal2 s 573794 -960 573906 480 8 la_data_out[125]
port 301 nsew default tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[126]
port 302 nsew default tristate
rlabel metal2 s 580970 -960 581082 480 8 la_data_out[127]
port 303 nsew default tristate
rlabel metal2 s 170558 -960 170670 480 8 la_data_out[12]
port 304 nsew default tristate
rlabel metal2 s 174146 -960 174258 480 8 la_data_out[13]
port 305 nsew default tristate
rlabel metal2 s 177734 -960 177846 480 8 la_data_out[14]
port 306 nsew default tristate
rlabel metal2 s 181322 -960 181434 480 8 la_data_out[15]
port 307 nsew default tristate
rlabel metal2 s 184818 -960 184930 480 8 la_data_out[16]
port 308 nsew default tristate
rlabel metal2 s 188406 -960 188518 480 8 la_data_out[17]
port 309 nsew default tristate
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[18]
port 310 nsew default tristate
rlabel metal2 s 195582 -960 195694 480 8 la_data_out[19]
port 311 nsew default tristate
rlabel metal2 s 131366 -960 131478 480 8 la_data_out[1]
port 312 nsew default tristate
rlabel metal2 s 199170 -960 199282 480 8 la_data_out[20]
port 313 nsew default tristate
rlabel metal2 s 202666 -960 202778 480 8 la_data_out[21]
port 314 nsew default tristate
rlabel metal2 s 206254 -960 206366 480 8 la_data_out[22]
port 315 nsew default tristate
rlabel metal2 s 209842 -960 209954 480 8 la_data_out[23]
port 316 nsew default tristate
rlabel metal2 s 213430 -960 213542 480 8 la_data_out[24]
port 317 nsew default tristate
rlabel metal2 s 217018 -960 217130 480 8 la_data_out[25]
port 318 nsew default tristate
rlabel metal2 s 220514 -960 220626 480 8 la_data_out[26]
port 319 nsew default tristate
rlabel metal2 s 224102 -960 224214 480 8 la_data_out[27]
port 320 nsew default tristate
rlabel metal2 s 227690 -960 227802 480 8 la_data_out[28]
port 321 nsew default tristate
rlabel metal2 s 231278 -960 231390 480 8 la_data_out[29]
port 322 nsew default tristate
rlabel metal2 s 134862 -960 134974 480 8 la_data_out[2]
port 323 nsew default tristate
rlabel metal2 s 234774 -960 234886 480 8 la_data_out[30]
port 324 nsew default tristate
rlabel metal2 s 238362 -960 238474 480 8 la_data_out[31]
port 325 nsew default tristate
rlabel metal2 s 241950 -960 242062 480 8 la_data_out[32]
port 326 nsew default tristate
rlabel metal2 s 245538 -960 245650 480 8 la_data_out[33]
port 327 nsew default tristate
rlabel metal2 s 249126 -960 249238 480 8 la_data_out[34]
port 328 nsew default tristate
rlabel metal2 s 252622 -960 252734 480 8 la_data_out[35]
port 329 nsew default tristate
rlabel metal2 s 256210 -960 256322 480 8 la_data_out[36]
port 330 nsew default tristate
rlabel metal2 s 259798 -960 259910 480 8 la_data_out[37]
port 331 nsew default tristate
rlabel metal2 s 263386 -960 263498 480 8 la_data_out[38]
port 332 nsew default tristate
rlabel metal2 s 266974 -960 267086 480 8 la_data_out[39]
port 333 nsew default tristate
rlabel metal2 s 138450 -960 138562 480 8 la_data_out[3]
port 334 nsew default tristate
rlabel metal2 s 270470 -960 270582 480 8 la_data_out[40]
port 335 nsew default tristate
rlabel metal2 s 274058 -960 274170 480 8 la_data_out[41]
port 336 nsew default tristate
rlabel metal2 s 277646 -960 277758 480 8 la_data_out[42]
port 337 nsew default tristate
rlabel metal2 s 281234 -960 281346 480 8 la_data_out[43]
port 338 nsew default tristate
rlabel metal2 s 284730 -960 284842 480 8 la_data_out[44]
port 339 nsew default tristate
rlabel metal2 s 288318 -960 288430 480 8 la_data_out[45]
port 340 nsew default tristate
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[46]
port 341 nsew default tristate
rlabel metal2 s 295494 -960 295606 480 8 la_data_out[47]
port 342 nsew default tristate
rlabel metal2 s 299082 -960 299194 480 8 la_data_out[48]
port 343 nsew default tristate
rlabel metal2 s 302578 -960 302690 480 8 la_data_out[49]
port 344 nsew default tristate
rlabel metal2 s 142038 -960 142150 480 8 la_data_out[4]
port 345 nsew default tristate
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[50]
port 346 nsew default tristate
rlabel metal2 s 309754 -960 309866 480 8 la_data_out[51]
port 347 nsew default tristate
rlabel metal2 s 313342 -960 313454 480 8 la_data_out[52]
port 348 nsew default tristate
rlabel metal2 s 316930 -960 317042 480 8 la_data_out[53]
port 349 nsew default tristate
rlabel metal2 s 320426 -960 320538 480 8 la_data_out[54]
port 350 nsew default tristate
rlabel metal2 s 324014 -960 324126 480 8 la_data_out[55]
port 351 nsew default tristate
rlabel metal2 s 327602 -960 327714 480 8 la_data_out[56]
port 352 nsew default tristate
rlabel metal2 s 331190 -960 331302 480 8 la_data_out[57]
port 353 nsew default tristate
rlabel metal2 s 334686 -960 334798 480 8 la_data_out[58]
port 354 nsew default tristate
rlabel metal2 s 338274 -960 338386 480 8 la_data_out[59]
port 355 nsew default tristate
rlabel metal2 s 145626 -960 145738 480 8 la_data_out[5]
port 356 nsew default tristate
rlabel metal2 s 341862 -960 341974 480 8 la_data_out[60]
port 357 nsew default tristate
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[61]
port 358 nsew default tristate
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[62]
port 359 nsew default tristate
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[63]
port 360 nsew default tristate
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[64]
port 361 nsew default tristate
rlabel metal2 s 359710 -960 359822 480 8 la_data_out[65]
port 362 nsew default tristate
rlabel metal2 s 363298 -960 363410 480 8 la_data_out[66]
port 363 nsew default tristate
rlabel metal2 s 366886 -960 366998 480 8 la_data_out[67]
port 364 nsew default tristate
rlabel metal2 s 370382 -960 370494 480 8 la_data_out[68]
port 365 nsew default tristate
rlabel metal2 s 373970 -960 374082 480 8 la_data_out[69]
port 366 nsew default tristate
rlabel metal2 s 149214 -960 149326 480 8 la_data_out[6]
port 367 nsew default tristate
rlabel metal2 s 377558 -960 377670 480 8 la_data_out[70]
port 368 nsew default tristate
rlabel metal2 s 381146 -960 381258 480 8 la_data_out[71]
port 369 nsew default tristate
rlabel metal2 s 384642 -960 384754 480 8 la_data_out[72]
port 370 nsew default tristate
rlabel metal2 s 388230 -960 388342 480 8 la_data_out[73]
port 371 nsew default tristate
rlabel metal2 s 391818 -960 391930 480 8 la_data_out[74]
port 372 nsew default tristate
rlabel metal2 s 395406 -960 395518 480 8 la_data_out[75]
port 373 nsew default tristate
rlabel metal2 s 398994 -960 399106 480 8 la_data_out[76]
port 374 nsew default tristate
rlabel metal2 s 402490 -960 402602 480 8 la_data_out[77]
port 375 nsew default tristate
rlabel metal2 s 406078 -960 406190 480 8 la_data_out[78]
port 376 nsew default tristate
rlabel metal2 s 409666 -960 409778 480 8 la_data_out[79]
port 377 nsew default tristate
rlabel metal2 s 152710 -960 152822 480 8 la_data_out[7]
port 378 nsew default tristate
rlabel metal2 s 413254 -960 413366 480 8 la_data_out[80]
port 379 nsew default tristate
rlabel metal2 s 416842 -960 416954 480 8 la_data_out[81]
port 380 nsew default tristate
rlabel metal2 s 420338 -960 420450 480 8 la_data_out[82]
port 381 nsew default tristate
rlabel metal2 s 423926 -960 424038 480 8 la_data_out[83]
port 382 nsew default tristate
rlabel metal2 s 427514 -960 427626 480 8 la_data_out[84]
port 383 nsew default tristate
rlabel metal2 s 431102 -960 431214 480 8 la_data_out[85]
port 384 nsew default tristate
rlabel metal2 s 434598 -960 434710 480 8 la_data_out[86]
port 385 nsew default tristate
rlabel metal2 s 438186 -960 438298 480 8 la_data_out[87]
port 386 nsew default tristate
rlabel metal2 s 441774 -960 441886 480 8 la_data_out[88]
port 387 nsew default tristate
rlabel metal2 s 445362 -960 445474 480 8 la_data_out[89]
port 388 nsew default tristate
rlabel metal2 s 156298 -960 156410 480 8 la_data_out[8]
port 389 nsew default tristate
rlabel metal2 s 448950 -960 449062 480 8 la_data_out[90]
port 390 nsew default tristate
rlabel metal2 s 452446 -960 452558 480 8 la_data_out[91]
port 391 nsew default tristate
rlabel metal2 s 456034 -960 456146 480 8 la_data_out[92]
port 392 nsew default tristate
rlabel metal2 s 459622 -960 459734 480 8 la_data_out[93]
port 393 nsew default tristate
rlabel metal2 s 463210 -960 463322 480 8 la_data_out[94]
port 394 nsew default tristate
rlabel metal2 s 466798 -960 466910 480 8 la_data_out[95]
port 395 nsew default tristate
rlabel metal2 s 470294 -960 470406 480 8 la_data_out[96]
port 396 nsew default tristate
rlabel metal2 s 473882 -960 473994 480 8 la_data_out[97]
port 397 nsew default tristate
rlabel metal2 s 477470 -960 477582 480 8 la_data_out[98]
port 398 nsew default tristate
rlabel metal2 s 481058 -960 481170 480 8 la_data_out[99]
port 399 nsew default tristate
rlabel metal2 s 159886 -960 159998 480 8 la_data_out[9]
port 400 nsew default tristate
rlabel metal2 s 128974 -960 129086 480 8 la_oen[0]
port 401 nsew default input
rlabel metal2 s 485750 -960 485862 480 8 la_oen[100]
port 402 nsew default input
rlabel metal2 s 489338 -960 489450 480 8 la_oen[101]
port 403 nsew default input
rlabel metal2 s 492926 -960 493038 480 8 la_oen[102]
port 404 nsew default input
rlabel metal2 s 496514 -960 496626 480 8 la_oen[103]
port 405 nsew default input
rlabel metal2 s 500102 -960 500214 480 8 la_oen[104]
port 406 nsew default input
rlabel metal2 s 503598 -960 503710 480 8 la_oen[105]
port 407 nsew default input
rlabel metal2 s 507186 -960 507298 480 8 la_oen[106]
port 408 nsew default input
rlabel metal2 s 510774 -960 510886 480 8 la_oen[107]
port 409 nsew default input
rlabel metal2 s 514362 -960 514474 480 8 la_oen[108]
port 410 nsew default input
rlabel metal2 s 517858 -960 517970 480 8 la_oen[109]
port 411 nsew default input
rlabel metal2 s 164670 -960 164782 480 8 la_oen[10]
port 412 nsew default input
rlabel metal2 s 521446 -960 521558 480 8 la_oen[110]
port 413 nsew default input
rlabel metal2 s 525034 -960 525146 480 8 la_oen[111]
port 414 nsew default input
rlabel metal2 s 528622 -960 528734 480 8 la_oen[112]
port 415 nsew default input
rlabel metal2 s 532210 -960 532322 480 8 la_oen[113]
port 416 nsew default input
rlabel metal2 s 535706 -960 535818 480 8 la_oen[114]
port 417 nsew default input
rlabel metal2 s 539294 -960 539406 480 8 la_oen[115]
port 418 nsew default input
rlabel metal2 s 542882 -960 542994 480 8 la_oen[116]
port 419 nsew default input
rlabel metal2 s 546470 -960 546582 480 8 la_oen[117]
port 420 nsew default input
rlabel metal2 s 550058 -960 550170 480 8 la_oen[118]
port 421 nsew default input
rlabel metal2 s 553554 -960 553666 480 8 la_oen[119]
port 422 nsew default input
rlabel metal2 s 168166 -960 168278 480 8 la_oen[11]
port 423 nsew default input
rlabel metal2 s 557142 -960 557254 480 8 la_oen[120]
port 424 nsew default input
rlabel metal2 s 560730 -960 560842 480 8 la_oen[121]
port 425 nsew default input
rlabel metal2 s 564318 -960 564430 480 8 la_oen[122]
port 426 nsew default input
rlabel metal2 s 567814 -960 567926 480 8 la_oen[123]
port 427 nsew default input
rlabel metal2 s 571402 -960 571514 480 8 la_oen[124]
port 428 nsew default input
rlabel metal2 s 574990 -960 575102 480 8 la_oen[125]
port 429 nsew default input
rlabel metal2 s 578578 -960 578690 480 8 la_oen[126]
port 430 nsew default input
rlabel metal2 s 582166 -960 582278 480 8 la_oen[127]
port 431 nsew default input
rlabel metal2 s 171754 -960 171866 480 8 la_oen[12]
port 432 nsew default input
rlabel metal2 s 175342 -960 175454 480 8 la_oen[13]
port 433 nsew default input
rlabel metal2 s 178930 -960 179042 480 8 la_oen[14]
port 434 nsew default input
rlabel metal2 s 182518 -960 182630 480 8 la_oen[15]
port 435 nsew default input
rlabel metal2 s 186014 -960 186126 480 8 la_oen[16]
port 436 nsew default input
rlabel metal2 s 189602 -960 189714 480 8 la_oen[17]
port 437 nsew default input
rlabel metal2 s 193190 -960 193302 480 8 la_oen[18]
port 438 nsew default input
rlabel metal2 s 196778 -960 196890 480 8 la_oen[19]
port 439 nsew default input
rlabel metal2 s 132562 -960 132674 480 8 la_oen[1]
port 440 nsew default input
rlabel metal2 s 200366 -960 200478 480 8 la_oen[20]
port 441 nsew default input
rlabel metal2 s 203862 -960 203974 480 8 la_oen[21]
port 442 nsew default input
rlabel metal2 s 207450 -960 207562 480 8 la_oen[22]
port 443 nsew default input
rlabel metal2 s 211038 -960 211150 480 8 la_oen[23]
port 444 nsew default input
rlabel metal2 s 214626 -960 214738 480 8 la_oen[24]
port 445 nsew default input
rlabel metal2 s 218122 -960 218234 480 8 la_oen[25]
port 446 nsew default input
rlabel metal2 s 221710 -960 221822 480 8 la_oen[26]
port 447 nsew default input
rlabel metal2 s 225298 -960 225410 480 8 la_oen[27]
port 448 nsew default input
rlabel metal2 s 228886 -960 228998 480 8 la_oen[28]
port 449 nsew default input
rlabel metal2 s 232474 -960 232586 480 8 la_oen[29]
port 450 nsew default input
rlabel metal2 s 136058 -960 136170 480 8 la_oen[2]
port 451 nsew default input
rlabel metal2 s 235970 -960 236082 480 8 la_oen[30]
port 452 nsew default input
rlabel metal2 s 239558 -960 239670 480 8 la_oen[31]
port 453 nsew default input
rlabel metal2 s 243146 -960 243258 480 8 la_oen[32]
port 454 nsew default input
rlabel metal2 s 246734 -960 246846 480 8 la_oen[33]
port 455 nsew default input
rlabel metal2 s 250322 -960 250434 480 8 la_oen[34]
port 456 nsew default input
rlabel metal2 s 253818 -960 253930 480 8 la_oen[35]
port 457 nsew default input
rlabel metal2 s 257406 -960 257518 480 8 la_oen[36]
port 458 nsew default input
rlabel metal2 s 260994 -960 261106 480 8 la_oen[37]
port 459 nsew default input
rlabel metal2 s 264582 -960 264694 480 8 la_oen[38]
port 460 nsew default input
rlabel metal2 s 268078 -960 268190 480 8 la_oen[39]
port 461 nsew default input
rlabel metal2 s 139646 -960 139758 480 8 la_oen[3]
port 462 nsew default input
rlabel metal2 s 271666 -960 271778 480 8 la_oen[40]
port 463 nsew default input
rlabel metal2 s 275254 -960 275366 480 8 la_oen[41]
port 464 nsew default input
rlabel metal2 s 278842 -960 278954 480 8 la_oen[42]
port 465 nsew default input
rlabel metal2 s 282430 -960 282542 480 8 la_oen[43]
port 466 nsew default input
rlabel metal2 s 285926 -960 286038 480 8 la_oen[44]
port 467 nsew default input
rlabel metal2 s 289514 -960 289626 480 8 la_oen[45]
port 468 nsew default input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[46]
port 469 nsew default input
rlabel metal2 s 296690 -960 296802 480 8 la_oen[47]
port 470 nsew default input
rlabel metal2 s 300278 -960 300390 480 8 la_oen[48]
port 471 nsew default input
rlabel metal2 s 303774 -960 303886 480 8 la_oen[49]
port 472 nsew default input
rlabel metal2 s 143234 -960 143346 480 8 la_oen[4]
port 473 nsew default input
rlabel metal2 s 307362 -960 307474 480 8 la_oen[50]
port 474 nsew default input
rlabel metal2 s 310950 -960 311062 480 8 la_oen[51]
port 475 nsew default input
rlabel metal2 s 314538 -960 314650 480 8 la_oen[52]
port 476 nsew default input
rlabel metal2 s 318034 -960 318146 480 8 la_oen[53]
port 477 nsew default input
rlabel metal2 s 321622 -960 321734 480 8 la_oen[54]
port 478 nsew default input
rlabel metal2 s 325210 -960 325322 480 8 la_oen[55]
port 479 nsew default input
rlabel metal2 s 328798 -960 328910 480 8 la_oen[56]
port 480 nsew default input
rlabel metal2 s 332386 -960 332498 480 8 la_oen[57]
port 481 nsew default input
rlabel metal2 s 335882 -960 335994 480 8 la_oen[58]
port 482 nsew default input
rlabel metal2 s 339470 -960 339582 480 8 la_oen[59]
port 483 nsew default input
rlabel metal2 s 146822 -960 146934 480 8 la_oen[5]
port 484 nsew default input
rlabel metal2 s 343058 -960 343170 480 8 la_oen[60]
port 485 nsew default input
rlabel metal2 s 346646 -960 346758 480 8 la_oen[61]
port 486 nsew default input
rlabel metal2 s 350234 -960 350346 480 8 la_oen[62]
port 487 nsew default input
rlabel metal2 s 353730 -960 353842 480 8 la_oen[63]
port 488 nsew default input
rlabel metal2 s 357318 -960 357430 480 8 la_oen[64]
port 489 nsew default input
rlabel metal2 s 360906 -960 361018 480 8 la_oen[65]
port 490 nsew default input
rlabel metal2 s 364494 -960 364606 480 8 la_oen[66]
port 491 nsew default input
rlabel metal2 s 367990 -960 368102 480 8 la_oen[67]
port 492 nsew default input
rlabel metal2 s 371578 -960 371690 480 8 la_oen[68]
port 493 nsew default input
rlabel metal2 s 375166 -960 375278 480 8 la_oen[69]
port 494 nsew default input
rlabel metal2 s 150410 -960 150522 480 8 la_oen[6]
port 495 nsew default input
rlabel metal2 s 378754 -960 378866 480 8 la_oen[70]
port 496 nsew default input
rlabel metal2 s 382342 -960 382454 480 8 la_oen[71]
port 497 nsew default input
rlabel metal2 s 385838 -960 385950 480 8 la_oen[72]
port 498 nsew default input
rlabel metal2 s 389426 -960 389538 480 8 la_oen[73]
port 499 nsew default input
rlabel metal2 s 393014 -960 393126 480 8 la_oen[74]
port 500 nsew default input
rlabel metal2 s 396602 -960 396714 480 8 la_oen[75]
port 501 nsew default input
rlabel metal2 s 400190 -960 400302 480 8 la_oen[76]
port 502 nsew default input
rlabel metal2 s 403686 -960 403798 480 8 la_oen[77]
port 503 nsew default input
rlabel metal2 s 407274 -960 407386 480 8 la_oen[78]
port 504 nsew default input
rlabel metal2 s 410862 -960 410974 480 8 la_oen[79]
port 505 nsew default input
rlabel metal2 s 153906 -960 154018 480 8 la_oen[7]
port 506 nsew default input
rlabel metal2 s 414450 -960 414562 480 8 la_oen[80]
port 507 nsew default input
rlabel metal2 s 417946 -960 418058 480 8 la_oen[81]
port 508 nsew default input
rlabel metal2 s 421534 -960 421646 480 8 la_oen[82]
port 509 nsew default input
rlabel metal2 s 425122 -960 425234 480 8 la_oen[83]
port 510 nsew default input
rlabel metal2 s 428710 -960 428822 480 8 la_oen[84]
port 511 nsew default input
rlabel metal2 s 432298 -960 432410 480 8 la_oen[85]
port 512 nsew default input
rlabel metal2 s 435794 -960 435906 480 8 la_oen[86]
port 513 nsew default input
rlabel metal2 s 439382 -960 439494 480 8 la_oen[87]
port 514 nsew default input
rlabel metal2 s 442970 -960 443082 480 8 la_oen[88]
port 515 nsew default input
rlabel metal2 s 446558 -960 446670 480 8 la_oen[89]
port 516 nsew default input
rlabel metal2 s 157494 -960 157606 480 8 la_oen[8]
port 517 nsew default input
rlabel metal2 s 450146 -960 450258 480 8 la_oen[90]
port 518 nsew default input
rlabel metal2 s 453642 -960 453754 480 8 la_oen[91]
port 519 nsew default input
rlabel metal2 s 457230 -960 457342 480 8 la_oen[92]
port 520 nsew default input
rlabel metal2 s 460818 -960 460930 480 8 la_oen[93]
port 521 nsew default input
rlabel metal2 s 464406 -960 464518 480 8 la_oen[94]
port 522 nsew default input
rlabel metal2 s 467902 -960 468014 480 8 la_oen[95]
port 523 nsew default input
rlabel metal2 s 471490 -960 471602 480 8 la_oen[96]
port 524 nsew default input
rlabel metal2 s 475078 -960 475190 480 8 la_oen[97]
port 525 nsew default input
rlabel metal2 s 478666 -960 478778 480 8 la_oen[98]
port 526 nsew default input
rlabel metal2 s 482254 -960 482366 480 8 la_oen[99]
port 527 nsew default input
rlabel metal2 s 161082 -960 161194 480 8 la_oen[9]
port 528 nsew default input
rlabel metal2 s 583362 -960 583474 480 8 user_clock2
port 529 nsew default input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 530 nsew default input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 531 nsew default input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 532 nsew default tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 533 nsew default input
rlabel metal2 s 48106 -960 48218 480 8 wbs_adr_i[10]
port 534 nsew default input
rlabel metal2 s 51602 -960 51714 480 8 wbs_adr_i[11]
port 535 nsew default input
rlabel metal2 s 55190 -960 55302 480 8 wbs_adr_i[12]
port 536 nsew default input
rlabel metal2 s 58778 -960 58890 480 8 wbs_adr_i[13]
port 537 nsew default input
rlabel metal2 s 62366 -960 62478 480 8 wbs_adr_i[14]
port 538 nsew default input
rlabel metal2 s 65954 -960 66066 480 8 wbs_adr_i[15]
port 539 nsew default input
rlabel metal2 s 69450 -960 69562 480 8 wbs_adr_i[16]
port 540 nsew default input
rlabel metal2 s 73038 -960 73150 480 8 wbs_adr_i[17]
port 541 nsew default input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[18]
port 542 nsew default input
rlabel metal2 s 80214 -960 80326 480 8 wbs_adr_i[19]
port 543 nsew default input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 544 nsew default input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[20]
port 545 nsew default input
rlabel metal2 s 87298 -960 87410 480 8 wbs_adr_i[21]
port 546 nsew default input
rlabel metal2 s 90886 -960 90998 480 8 wbs_adr_i[22]
port 547 nsew default input
rlabel metal2 s 94474 -960 94586 480 8 wbs_adr_i[23]
port 548 nsew default input
rlabel metal2 s 98062 -960 98174 480 8 wbs_adr_i[24]
port 549 nsew default input
rlabel metal2 s 101558 -960 101670 480 8 wbs_adr_i[25]
port 550 nsew default input
rlabel metal2 s 105146 -960 105258 480 8 wbs_adr_i[26]
port 551 nsew default input
rlabel metal2 s 108734 -960 108846 480 8 wbs_adr_i[27]
port 552 nsew default input
rlabel metal2 s 112322 -960 112434 480 8 wbs_adr_i[28]
port 553 nsew default input
rlabel metal2 s 115910 -960 116022 480 8 wbs_adr_i[29]
port 554 nsew default input
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[2]
port 555 nsew default input
rlabel metal2 s 119406 -960 119518 480 8 wbs_adr_i[30]
port 556 nsew default input
rlabel metal2 s 122994 -960 123106 480 8 wbs_adr_i[31]
port 557 nsew default input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 558 nsew default input
rlabel metal2 s 26670 -960 26782 480 8 wbs_adr_i[4]
port 559 nsew default input
rlabel metal2 s 30258 -960 30370 480 8 wbs_adr_i[5]
port 560 nsew default input
rlabel metal2 s 33846 -960 33958 480 8 wbs_adr_i[6]
port 561 nsew default input
rlabel metal2 s 37342 -960 37454 480 8 wbs_adr_i[7]
port 562 nsew default input
rlabel metal2 s 40930 -960 41042 480 8 wbs_adr_i[8]
port 563 nsew default input
rlabel metal2 s 44518 -960 44630 480 8 wbs_adr_i[9]
port 564 nsew default input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 565 nsew default input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 566 nsew default input
rlabel metal2 s 49302 -960 49414 480 8 wbs_dat_i[10]
port 567 nsew default input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_i[11]
port 568 nsew default input
rlabel metal2 s 56386 -960 56498 480 8 wbs_dat_i[12]
port 569 nsew default input
rlabel metal2 s 59974 -960 60086 480 8 wbs_dat_i[13]
port 570 nsew default input
rlabel metal2 s 63562 -960 63674 480 8 wbs_dat_i[14]
port 571 nsew default input
rlabel metal2 s 67150 -960 67262 480 8 wbs_dat_i[15]
port 572 nsew default input
rlabel metal2 s 70646 -960 70758 480 8 wbs_dat_i[16]
port 573 nsew default input
rlabel metal2 s 74234 -960 74346 480 8 wbs_dat_i[17]
port 574 nsew default input
rlabel metal2 s 77822 -960 77934 480 8 wbs_dat_i[18]
port 575 nsew default input
rlabel metal2 s 81410 -960 81522 480 8 wbs_dat_i[19]
port 576 nsew default input
rlabel metal2 s 13606 -960 13718 480 8 wbs_dat_i[1]
port 577 nsew default input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[20]
port 578 nsew default input
rlabel metal2 s 88494 -960 88606 480 8 wbs_dat_i[21]
port 579 nsew default input
rlabel metal2 s 92082 -960 92194 480 8 wbs_dat_i[22]
port 580 nsew default input
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_i[23]
port 581 nsew default input
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_i[24]
port 582 nsew default input
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_i[25]
port 583 nsew default input
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_i[26]
port 584 nsew default input
rlabel metal2 s 109930 -960 110042 480 8 wbs_dat_i[27]
port 585 nsew default input
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_i[28]
port 586 nsew default input
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_i[29]
port 587 nsew default input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 588 nsew default input
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_i[30]
port 589 nsew default input
rlabel metal2 s 124190 -960 124302 480 8 wbs_dat_i[31]
port 590 nsew default input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 591 nsew default input
rlabel metal2 s 27866 -960 27978 480 8 wbs_dat_i[4]
port 592 nsew default input
rlabel metal2 s 31454 -960 31566 480 8 wbs_dat_i[5]
port 593 nsew default input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 594 nsew default input
rlabel metal2 s 38538 -960 38650 480 8 wbs_dat_i[7]
port 595 nsew default input
rlabel metal2 s 42126 -960 42238 480 8 wbs_dat_i[8]
port 596 nsew default input
rlabel metal2 s 45714 -960 45826 480 8 wbs_dat_i[9]
port 597 nsew default input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 598 nsew default tristate
rlabel metal2 s 50498 -960 50610 480 8 wbs_dat_o[10]
port 599 nsew default tristate
rlabel metal2 s 53994 -960 54106 480 8 wbs_dat_o[11]
port 600 nsew default tristate
rlabel metal2 s 57582 -960 57694 480 8 wbs_dat_o[12]
port 601 nsew default tristate
rlabel metal2 s 61170 -960 61282 480 8 wbs_dat_o[13]
port 602 nsew default tristate
rlabel metal2 s 64758 -960 64870 480 8 wbs_dat_o[14]
port 603 nsew default tristate
rlabel metal2 s 68254 -960 68366 480 8 wbs_dat_o[15]
port 604 nsew default tristate
rlabel metal2 s 71842 -960 71954 480 8 wbs_dat_o[16]
port 605 nsew default tristate
rlabel metal2 s 75430 -960 75542 480 8 wbs_dat_o[17]
port 606 nsew default tristate
rlabel metal2 s 79018 -960 79130 480 8 wbs_dat_o[18]
port 607 nsew default tristate
rlabel metal2 s 82606 -960 82718 480 8 wbs_dat_o[19]
port 608 nsew default tristate
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[1]
port 609 nsew default tristate
rlabel metal2 s 86102 -960 86214 480 8 wbs_dat_o[20]
port 610 nsew default tristate
rlabel metal2 s 89690 -960 89802 480 8 wbs_dat_o[21]
port 611 nsew default tristate
rlabel metal2 s 93278 -960 93390 480 8 wbs_dat_o[22]
port 612 nsew default tristate
rlabel metal2 s 96866 -960 96978 480 8 wbs_dat_o[23]
port 613 nsew default tristate
rlabel metal2 s 100454 -960 100566 480 8 wbs_dat_o[24]
port 614 nsew default tristate
rlabel metal2 s 103950 -960 104062 480 8 wbs_dat_o[25]
port 615 nsew default tristate
rlabel metal2 s 107538 -960 107650 480 8 wbs_dat_o[26]
port 616 nsew default tristate
rlabel metal2 s 111126 -960 111238 480 8 wbs_dat_o[27]
port 617 nsew default tristate
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_o[28]
port 618 nsew default tristate
rlabel metal2 s 118210 -960 118322 480 8 wbs_dat_o[29]
port 619 nsew default tristate
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 620 nsew default tristate
rlabel metal2 s 121798 -960 121910 480 8 wbs_dat_o[30]
port 621 nsew default tristate
rlabel metal2 s 125386 -960 125498 480 8 wbs_dat_o[31]
port 622 nsew default tristate
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 623 nsew default tristate
rlabel metal2 s 29062 -960 29174 480 8 wbs_dat_o[4]
port 624 nsew default tristate
rlabel metal2 s 32650 -960 32762 480 8 wbs_dat_o[5]
port 625 nsew default tristate
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 626 nsew default tristate
rlabel metal2 s 39734 -960 39846 480 8 wbs_dat_o[7]
port 627 nsew default tristate
rlabel metal2 s 43322 -960 43434 480 8 wbs_dat_o[8]
port 628 nsew default tristate
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_o[9]
port 629 nsew default tristate
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 630 nsew default input
rlabel metal2 s 15998 -960 16110 480 8 wbs_sel_i[1]
port 631 nsew default input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 632 nsew default input
rlabel metal2 s 25474 -960 25586 480 8 wbs_sel_i[3]
port 633 nsew default input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 634 nsew default input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 635 nsew default input
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 636 nsew default input
rlabel metal5 s -2916 -1844 586840 -1244 8 vssd1
port 637 nsew default input
rlabel metal5 s -3836 -2764 587760 -2164 8 vccd2
port 638 nsew default input
rlabel metal5 s -4756 -3684 588680 -3084 8 vssd2
port 639 nsew default input
rlabel metal5 s -5676 -4604 589600 -4004 8 vdda1
port 640 nsew default input
rlabel metal5 s -6596 -5524 590520 -4924 8 vssa1
port 641 nsew default input
rlabel metal5 s -7516 -6444 591440 -5844 8 vdda2
port 642 nsew default input
rlabel metal5 s -8436 -7364 592360 -6764 8 vssa2
port 643 nsew default input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
